module AHB_Lite_2s (
	HCLK, 
	HRESETn, 
	HADDR, 
	HBURST, 
	HMASTLOCK, 
	HPROT, 
	HSIZE, 
	HTRANS, 
	HWDATA, 
	HWRITE, 
	hsel_s1, 
	hready_resp_s1, 
	hresp_s1, 
	hrdata_s1, 
	hsel_s2, 
	hready_resp_s2, 
	hresp_s2, 
	hrdata_s2, 
	haddr_s, 
	hburst_s, 
	hprot_s, 
	hsize_s, 
	htrans_s, 
	hwdata_s, 
	hwrite_s, 
	HREADY, 
	hresp_ahb, 
	HRDATA, 
	hmaster, 
	hmaster_data, 
	hmastlock_s, 
	FE_OFN114_HADDR_29_, 
	FE_OFN119_HADDR_31_);
   input HCLK;
   input HRESETn;
   input [31:0] HADDR;
   input [2:0] HBURST;
   input HMASTLOCK;
   input [3:0] HPROT;
   input [2:0] HSIZE;
   input [1:0] HTRANS;
   input [31:0] HWDATA;
   input HWRITE;
   output hsel_s1;
   input hready_resp_s1;
   input [1:0] hresp_s1;
   input [31:0] hrdata_s1;
   output hsel_s2;
   input hready_resp_s2;
   input [1:0] hresp_s2;
   input [31:0] hrdata_s2;
   output [31:0] haddr_s;
   output [2:0] hburst_s;
   output [3:0] hprot_s;
   output [2:0] hsize_s;
   output [1:0] htrans_s;
   output [31:0] hwdata_s;
   output hwrite_s;
   inout HREADY;
   output [1:0] hresp_ahb;
   output [31:0] HRDATA;
   output [3:0] hmaster;
   output [3:0] hmaster_data;
   output hmastlock_s;
   input FE_OFN114_HADDR_29_;
   input FE_OFN119_HADDR_31_;

   // Internal wires
   wire FE_PHN692_hrdata_s1_20_;
   wire FE_PHN688_hrdata_s1_17_;
   wire FE_PHN681_hrdata_s1_24_;
   wire FE_OFN122_hsel_s2;
   wire FE_OFN121_hsel_s2;
   wire FE_OFN120_HADDR_31_;
   wire FE_OFN116_HADDR_29_;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;

   assign HREADY = hready_resp_s1 ;
   assign htrans_s[0] = 1'b0 ;
   assign hsize_s[2] = 1'b0 ;

   BUF_X32 FE_PHC692_hrdata_s1_20_ (.Z(FE_PHN692_hrdata_s1_20_), 
	.A(hrdata_s1[20]));
   BUF_X32 FE_PHC688_hrdata_s1_17_ (.Z(FE_PHN688_hrdata_s1_17_), 
	.A(hrdata_s1[17]));
   BUF_X32 FE_PHC681_hrdata_s1_24_ (.Z(FE_PHN681_hrdata_s1_24_), 
	.A(hrdata_s1[24]));
   INV_X4 FE_OFC122_hsel_s2 (.ZN(hsel_s2), 
	.A(FE_OFN122_hsel_s2));
   INV_X4 FE_OFC121_hsel_s2 (.ZN(FE_OFN122_hsel_s2), 
	.A(FE_OFN121_hsel_s2));
   INV_X8 FE_OFC119_HADDR_31_ (.ZN(FE_OFN120_HADDR_31_), 
	.A(FE_OFN119_HADDR_31_));
   INV_X4 FE_OFC116_HADDR_29_ (.ZN(FE_OFN116_HADDR_29_), 
	.A(FE_OFN114_HADDR_29_));
   NOR3_X4 U92 (.ZN(hsel_s1), 
	.A3(FE_OFN116_HADDR_29_), 
	.A2(FE_OFN120_HADDR_31_), 
	.A1(HADDR[30]));
   INV_X4 U93 (.ZN(HRDATA[31]), 
	.A(n377));
   INV_X4 U94 (.ZN(HRDATA[30]), 
	.A(n378));
   INV_X4 U95 (.ZN(HRDATA[29]), 
	.A(n380));
   INV_X4 U96 (.ZN(HRDATA[28]), 
	.A(n381));
   INV_X4 U97 (.ZN(HRDATA[27]), 
	.A(n382));
   INV_X4 U98 (.ZN(HRDATA[26]), 
	.A(n383));
   INV_X4 U99 (.ZN(HRDATA[25]), 
	.A(n384));
   INV_X4 U100 (.ZN(HRDATA[24]), 
	.A(n385));
   INV_X4 U101 (.ZN(HRDATA[23]), 
	.A(n386));
   INV_X4 U102 (.ZN(HRDATA[22]), 
	.A(n387));
   INV_X4 U103 (.ZN(HRDATA[21]), 
	.A(n388));
   INV_X4 U104 (.ZN(HRDATA[20]), 
	.A(n389));
   INV_X4 U105 (.ZN(HRDATA[19]), 
	.A(n391));
   INV_X4 U106 (.ZN(HRDATA[18]), 
	.A(n392));
   INV_X4 U107 (.ZN(HRDATA[17]), 
	.A(n393));
   INV_X4 U108 (.ZN(HRDATA[16]), 
	.A(n394));
   INV_X4 U109 (.ZN(HRDATA[15]), 
	.A(n395));
   INV_X4 U110 (.ZN(HRDATA[14]), 
	.A(n396));
   INV_X4 U111 (.ZN(HRDATA[13]), 
	.A(n397));
   INV_X4 U112 (.ZN(HRDATA[12]), 
	.A(n398));
   INV_X4 U113 (.ZN(HRDATA[11]), 
	.A(n399));
   INV_X4 U114 (.ZN(HRDATA[10]), 
	.A(n400));
   INV_X4 U115 (.ZN(HRDATA[9]), 
	.A(n371));
   INV_X4 U116 (.ZN(HRDATA[8]), 
	.A(n372));
   INV_X4 U117 (.ZN(HRDATA[7]), 
	.A(n373));
   INV_X4 U118 (.ZN(HRDATA[6]), 
	.A(n374));
   INV_X4 U119 (.ZN(HRDATA[5]), 
	.A(n375));
   INV_X4 U120 (.ZN(HRDATA[4]), 
	.A(n376));
   INV_X4 U121 (.ZN(HRDATA[3]), 
	.A(n379));
   INV_X4 U122 (.ZN(HRDATA[2]), 
	.A(n390));
   INV_X4 U123 (.ZN(HRDATA[1]), 
	.A(n401));
   INV_X4 U124 (.ZN(HRDATA[0]), 
	.A(n402));
   NOR3_X4 U125 (.ZN(FE_OFN121_hsel_s2), 
	.A3(n403), 
	.A2(FE_OFN120_HADDR_31_), 
	.A1(FE_OFN116_HADDR_29_));
   BUF_X2 U126 (.Z(haddr_s[31]), 
	.A(HADDR[31]));
   BUF_X2 U127 (.Z(haddr_s[30]), 
	.A(HADDR[30]));
   BUF_X2 U128 (.Z(haddr_s[29]), 
	.A(HADDR[29]));
   BUF_X2 U129 (.Z(haddr_s[28]), 
	.A(HADDR[28]));
   BUF_X2 U130 (.Z(haddr_s[27]), 
	.A(HADDR[27]));
   BUF_X2 U131 (.Z(haddr_s[26]), 
	.A(HADDR[26]));
   BUF_X2 U132 (.Z(haddr_s[25]), 
	.A(HADDR[25]));
   BUF_X2 U133 (.Z(haddr_s[24]), 
	.A(HADDR[24]));
   BUF_X2 U134 (.Z(haddr_s[23]), 
	.A(HADDR[23]));
   BUF_X2 U135 (.Z(haddr_s[22]), 
	.A(HADDR[22]));
   BUF_X2 U136 (.Z(haddr_s[21]), 
	.A(HADDR[21]));
   BUF_X2 U137 (.Z(haddr_s[20]), 
	.A(HADDR[20]));
   BUF_X2 U138 (.Z(haddr_s[19]), 
	.A(HADDR[19]));
   BUF_X2 U139 (.Z(haddr_s[18]), 
	.A(HADDR[18]));
   BUF_X2 U140 (.Z(haddr_s[17]), 
	.A(HADDR[17]));
   BUF_X2 U141 (.Z(haddr_s[16]), 
	.A(HADDR[16]));
   BUF_X2 U142 (.Z(haddr_s[15]), 
	.A(HADDR[15]));
   BUF_X2 U143 (.Z(haddr_s[14]), 
	.A(HADDR[14]));
   BUF_X2 U144 (.Z(haddr_s[13]), 
	.A(HADDR[13]));
   BUF_X2 U145 (.Z(haddr_s[12]), 
	.A(HADDR[12]));
   BUF_X2 U146 (.Z(haddr_s[11]), 
	.A(HADDR[11]));
   BUF_X2 U147 (.Z(haddr_s[10]), 
	.A(HADDR[10]));
   BUF_X2 U148 (.Z(haddr_s[9]), 
	.A(HADDR[9]));
   BUF_X2 U149 (.Z(haddr_s[8]), 
	.A(HADDR[8]));
   BUF_X2 U150 (.Z(haddr_s[7]), 
	.A(HADDR[7]));
   BUF_X2 U151 (.Z(haddr_s[6]), 
	.A(HADDR[6]));
   BUF_X2 U152 (.Z(haddr_s[5]), 
	.A(HADDR[5]));
   BUF_X2 U153 (.Z(haddr_s[4]), 
	.A(HADDR[4]));
   BUF_X2 U154 (.Z(haddr_s[3]), 
	.A(HADDR[3]));
   BUF_X2 U155 (.Z(haddr_s[2]), 
	.A(HADDR[2]));
   BUF_X2 U156 (.Z(haddr_s[1]), 
	.A(HADDR[1]));
   BUF_X2 U157 (.Z(haddr_s[0]), 
	.A(HADDR[0]));
   BUF_X2 U166 (.Z(hsize_s[1]), 
	.A(HSIZE[1]));
   BUF_X2 U167 (.Z(hsize_s[0]), 
	.A(HSIZE[0]));
   BUF_X2 U168 (.Z(htrans_s[1]), 
	.A(HTRANS[1]));
   BUF_X2 U170 (.Z(hwdata_s[31]), 
	.A(HWDATA[31]));
   BUF_X2 U171 (.Z(hwdata_s[30]), 
	.A(HWDATA[30]));
   BUF_X2 U172 (.Z(hwdata_s[29]), 
	.A(HWDATA[29]));
   BUF_X2 U173 (.Z(hwdata_s[28]), 
	.A(HWDATA[28]));
   BUF_X2 U174 (.Z(hwdata_s[27]), 
	.A(HWDATA[27]));
   BUF_X2 U175 (.Z(hwdata_s[26]), 
	.A(HWDATA[26]));
   BUF_X2 U176 (.Z(hwdata_s[25]), 
	.A(HWDATA[25]));
   BUF_X2 U177 (.Z(hwdata_s[24]), 
	.A(HWDATA[24]));
   BUF_X2 U178 (.Z(hwdata_s[23]), 
	.A(HWDATA[23]));
   BUF_X2 U179 (.Z(hwdata_s[22]), 
	.A(HWDATA[22]));
   BUF_X2 U180 (.Z(hwdata_s[21]), 
	.A(HWDATA[21]));
   BUF_X2 U181 (.Z(hwdata_s[20]), 
	.A(HWDATA[20]));
   BUF_X2 U182 (.Z(hwdata_s[19]), 
	.A(HWDATA[19]));
   BUF_X2 U183 (.Z(hwdata_s[18]), 
	.A(HWDATA[18]));
   BUF_X2 U184 (.Z(hwdata_s[17]), 
	.A(HWDATA[17]));
   BUF_X2 U185 (.Z(hwdata_s[16]), 
	.A(HWDATA[16]));
   BUF_X2 U186 (.Z(hwdata_s[15]), 
	.A(HWDATA[15]));
   BUF_X2 U187 (.Z(hwdata_s[14]), 
	.A(HWDATA[14]));
   BUF_X2 U188 (.Z(hwdata_s[13]), 
	.A(HWDATA[13]));
   BUF_X2 U189 (.Z(hwdata_s[12]), 
	.A(HWDATA[12]));
   BUF_X2 U190 (.Z(hwdata_s[11]), 
	.A(HWDATA[11]));
   BUF_X2 U191 (.Z(hwdata_s[10]), 
	.A(HWDATA[10]));
   BUF_X2 U192 (.Z(hwdata_s[9]), 
	.A(HWDATA[9]));
   BUF_X2 U193 (.Z(hwdata_s[8]), 
	.A(HWDATA[8]));
   BUF_X2 U194 (.Z(hwdata_s[7]), 
	.A(HWDATA[7]));
   BUF_X2 U195 (.Z(hwdata_s[6]), 
	.A(HWDATA[6]));
   BUF_X2 U196 (.Z(hwdata_s[5]), 
	.A(HWDATA[5]));
   BUF_X2 U197 (.Z(hwdata_s[4]), 
	.A(HWDATA[4]));
   BUF_X2 U198 (.Z(hwdata_s[3]), 
	.A(HWDATA[3]));
   BUF_X2 U199 (.Z(hwdata_s[2]), 
	.A(HWDATA[2]));
   BUF_X2 U200 (.Z(hwdata_s[1]), 
	.A(HWDATA[1]));
   BUF_X2 U201 (.Z(hwdata_s[0]), 
	.A(HWDATA[0]));
   BUF_X2 U202 (.Z(hwrite_s), 
	.A(HWRITE));
   AOI22_X1 U203 (.ZN(n371), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[9]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[9]));
   AOI22_X1 U204 (.ZN(n372), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[8]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[8]));
   AOI22_X1 U205 (.ZN(n373), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[7]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[7]));
   AOI22_X1 U206 (.ZN(n374), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[6]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[6]));
   AOI22_X1 U207 (.ZN(n375), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[5]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[5]));
   AOI22_X1 U208 (.ZN(n376), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[4]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[4]));
   AOI22_X1 U209 (.ZN(n377), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[31]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[31]));
   AOI22_X1 U210 (.ZN(n378), 
	.B2(hsel_s2), 
	.B1(hrdata_s2[30]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[30]));
   AOI22_X1 U211 (.ZN(n379), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[3]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[3]));
   AOI22_X1 U212 (.ZN(n380), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[29]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[29]));
   AOI22_X1 U213 (.ZN(n381), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[28]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[28]));
   AOI22_X1 U214 (.ZN(n382), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[27]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[27]));
   AOI22_X1 U215 (.ZN(n383), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[26]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[26]));
   AOI22_X1 U216 (.ZN(n384), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[25]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[25]));
   AOI22_X1 U217 (.ZN(n385), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[24]), 
	.A2(hsel_s1), 
	.A1(FE_PHN681_hrdata_s1_24_));
   AOI22_X1 U218 (.ZN(n386), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[23]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[23]));
   AOI22_X1 U219 (.ZN(n387), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[22]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[22]));
   AOI22_X1 U220 (.ZN(n388), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[21]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[21]));
   AOI22_X1 U221 (.ZN(n389), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[20]), 
	.A2(hsel_s1), 
	.A1(FE_PHN692_hrdata_s1_20_));
   AOI22_X1 U222 (.ZN(n390), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[2]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[2]));
   AOI22_X1 U223 (.ZN(n391), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[19]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[19]));
   AOI22_X1 U224 (.ZN(n392), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[18]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[18]));
   AOI22_X1 U225 (.ZN(n393), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[17]), 
	.A2(hsel_s1), 
	.A1(FE_PHN688_hrdata_s1_17_));
   AOI22_X1 U226 (.ZN(n394), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[16]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[16]));
   AOI22_X1 U227 (.ZN(n395), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[15]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[15]));
   AOI22_X1 U228 (.ZN(n396), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[14]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[14]));
   AOI22_X1 U229 (.ZN(n397), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[13]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[13]));
   AOI22_X1 U230 (.ZN(n398), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[12]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[12]));
   AOI22_X1 U231 (.ZN(n399), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[11]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[11]));
   AOI22_X1 U232 (.ZN(n400), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[10]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[10]));
   AOI22_X1 U233 (.ZN(n401), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[1]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[1]));
   AOI22_X1 U234 (.ZN(n402), 
	.B2(FE_OFN121_hsel_s2), 
	.B1(hrdata_s2[0]), 
	.A2(hsel_s1), 
	.A1(hrdata_s1[0]));
   INV_X1 U235 (.ZN(n403), 
	.A(HADDR[30]));
endmodule

module DW_memctl_hiu (
	hclk, 
	hresetn, 
	hsel_mem, 
	hsel_reg, 
	htrans, 
	hwrite, 
	hsize, 
	hburst, 
	hready, 
	hready_resp, 
	hresp, 
	haddr, 
	hwdata, 
	hrdata, 
	hiu_req, 
	hiu_burst_size, 
	hiu_wrap_burst, 
	hiu_rw, 
	hiu_terminate, 
	hiu_addr, 
	hiu_data, 
	hiu_haddr, 
	hiu_hsize, 
	miu_burst_done, 
	miu_push_n, 
	miu_pop_n, 
	miu_data, 
	miu_data_width, 
	miu_col_width, 
	big_endian, 
	FE_OFN28_HRESETn, 
	FE_OFN29_HRESETn, 
	FE_OFN30_HRESETn, 
	FE_OFN34_HRESETn, 
	FE_OFN42_HRESETn, 
	FE_OFN43_HRESETn, 
	FE_OFN55_HRESETn, 
	FE_OFN31_HRESETn, 
	FE_OFN35_HRESETn, 
	FE_OFN46_HRESETn, 
	FE_OFN51_HRESETn, 
	FE_OFN53_HRESETn, 
	FE_OFN57_HRESETn, 
	HCLK__L5_N14, 
	HCLK__L5_N15, 
	HCLK__L5_N16, 
	HCLK__L5_N17, 
	HCLK__L5_N18, 
	HCLK__L5_N27, 
	HCLK__L5_N32, 
	HCLK__L5_N33, 
	HCLK__L5_N34, 
	HCLK__L5_N35, 
	HCLK__L5_N36, 
	HCLK__L5_N37, 
	HCLK__L5_N38, 
	HCLK__L5_N39, 
	HCLK__L5_N4, 
	HCLK__L5_N5, 
	HCLK__L5_N6, 
	FE_OFN151_HRESETn, 
	FE_OFN160_HRESETn, 
	FE_OFN191_HRESETn, 
	FE_OFN214_hiu_burst_size_4_, 
	FE_OFN217_hiu_burst_size_2_, 
	FE_OFN220_hiu_burst_size_0_);
   input hclk;
   input hresetn;
   input hsel_mem;
   input hsel_reg;
   input [1:0] htrans;
   input hwrite;
   input [2:0] hsize;
   input [2:0] hburst;
   input hready;
   output hready_resp;
   output [1:0] hresp;
   input [31:0] haddr;
   input [31:0] hwdata;
   output [31:0] hrdata;
   output [1:0] hiu_req;
   output [5:0] hiu_burst_size;
   output hiu_wrap_burst;
   output hiu_rw;
   output hiu_terminate;
   output [31:0] hiu_addr;
   output [31:0] hiu_data;
   output [3:0] hiu_haddr;
   output [2:0] hiu_hsize;
   input miu_burst_done;
   input miu_push_n;
   input miu_pop_n;
   input [31:0] miu_data;
   input [1:0] miu_data_width;
   input [3:0] miu_col_width;
   input big_endian;
   input FE_OFN28_HRESETn;
   input FE_OFN29_HRESETn;
   input FE_OFN30_HRESETn;
   input FE_OFN34_HRESETn;
   input FE_OFN42_HRESETn;
   input FE_OFN43_HRESETn;
   input FE_OFN55_HRESETn;
   input FE_OFN31_HRESETn;
   input FE_OFN35_HRESETn;
   input FE_OFN46_HRESETn;
   input FE_OFN51_HRESETn;
   input FE_OFN53_HRESETn;
   input FE_OFN57_HRESETn;
   input HCLK__L5_N14;
   input HCLK__L5_N15;
   input HCLK__L5_N16;
   input HCLK__L5_N17;
   input HCLK__L5_N18;
   input HCLK__L5_N27;
   input HCLK__L5_N32;
   input HCLK__L5_N33;
   input HCLK__L5_N34;
   input HCLK__L5_N35;
   input HCLK__L5_N36;
   input HCLK__L5_N37;
   input HCLK__L5_N38;
   input HCLK__L5_N39;
   input HCLK__L5_N4;
   input HCLK__L5_N5;
   input HCLK__L5_N6;
   input FE_OFN151_HRESETn;
   input FE_OFN160_HRESETn;
   input FE_OFN191_HRESETn;
   input FE_OFN214_hiu_burst_size_4_;
   input FE_OFN217_hiu_burst_size_2_;
   input FE_OFN220_hiu_burst_size_0_;

   // Internal wires
   wire FE_PHN5241_U_rbuf_n175;
   wire FE_PHN5240_U_rbuf_n69;
   wire FE_PHN5239_U_ctl_n299;
   wire FE_PHN5218_U_ctl_N89;
   wire FE_PHN5203_U_ctl_n299;
   wire FE_PHN5191_miu_data_27_;
   wire FE_PHN5190_U_rbuf_n69;
   wire FE_PHN5189_U_rbuf_n175;
   wire FE_PHN5181_hsel_reg;
   wire FE_PHN5180_U_rbuf_n63;
   wire FE_PHN5179_U_rbuf_n72;
   wire FE_PHN5175_U_rbuf_n188;
   wire FE_PHN5165_U_afifo_U_acore_U_sub_fifo_n282;
   wire FE_PHN5164_U_afifo_U_acore_U_sub_fifo_n260;
   wire FE_PHN5162_U_afifo_U_acore_U_sub_fifo_n316;
   wire FE_PHN5159_U_dfifo_U_dcore_U_sub_fifo_n275;
   wire FE_PHN5157_U_dfifo_U_dcore_U_sub_fifo_n299;
   wire FE_PHN5154_U_afifo_U_acore_U_sub_fifo_n249;
   wire FE_PHN5153_U_afifo_U_acore_U_sub_fifo_n209;
   wire FE_PHN5152_U_afifo_U_acore_U_sub_fifo_n294;
   wire FE_PHN5148_U_dfifo_U_dcore_U_sub_fifo_n257;
   wire FE_PHN5147_U_dfifo_U_dcore_U_sub_fifo_n259;
   wire FE_PHN5143_U_afifo_U_acore_U_sub_fifo_n188;
   wire FE_PHN5140_U_afifo_U_acore_U_sub_fifo_n245;
   wire FE_PHN5138_U_dfifo_U_dcore_U_sub_fifo_n307;
   wire FE_PHN5133_U_afifo_U_acore_U_sub_fifo_n236;
   wire FE_PHN5132_U_afifo_n158;
   wire FE_PHN5128_U_dfifo_U_dcore_U_sub_fifo_n251;
   wire FE_PHN5118_U_afifo_U_acore_U_sub_fifo_n250;
   wire FE_PHN5117_U_afifo_U_acore_U_sub_fifo_n275;
   wire FE_PHN5116_U_dfifo_U_dcore_U_sub_fifo_n247;
   wire FE_PHN5115_U_dfifo_U_dcore_U_sub_fifo_n292;
   wire FE_PHN5111_U_afifo_U_acore_U_sub_fifo_n220;
   wire FE_PHN5109_U_dfifo_U_dcore_U_sub_fifo_n310;
   wire FE_PHN5103_U_afifo_U_acore_U_sub_fifo_n308;
   wire FE_PHN5101_U_afifo_U_acore_U_sub_fifo_n177;
   wire FE_PHN5100_U_afifo_n159;
   wire FE_PHN5098_U_afifo_U_acore_U_sub_fifo_n251;
   wire FE_PHN5095_U_afifo_U_acore_U_sub_fifo_n194;
   wire FE_PHN5092_U_dfifo_U_dcore_U_sub_fifo_n287;
   wire FE_PHN5087_U_afifo_U_acore_U_sub_fifo_n265;
   wire FE_PHN5083_U_dfifo_U_dcore_U_sub_fifo_n274;
   wire FE_PHN5082_U_dfifo_U_dcore_U_sub_fifo_n280;
   wire FE_PHN5081_U_afifo_U_acore_U_sub_fifo_n309;
   wire FE_PHN5079_U_afifo_U_acore_U_sub_fifo_n231;
   wire FE_PHN5078_U_afifo_U_acore_U_sub_fifo_n246;
   wire FE_PHN5075_U_afifo_U_acore_U_sub_fifo_n213;
   wire FE_PHN5073_U_afifo_U_acore_U_sub_fifo_n180;
   wire FE_PHN5072_U_dfifo_U_dcore_U_sub_fifo_n263;
   wire FE_PHN5071_U_afifo_U_acore_U_sub_fifo_n264;
   wire FE_PHN5070_U_dfifo_U_dcore_U_sub_fifo_n308;
   wire FE_PHN5069_U_afifo_U_acore_U_sub_fifo_n185;
   wire FE_PHN5068_U_afifo_U_acore_U_sub_fifo_n243;
   wire FE_PHN5067_U_afifo_U_acore_U_sub_fifo_n307;
   wire FE_PHN5063_U_afifo_U_acore_U_sub_fifo_n227;
   wire FE_PHN5062_U_dfifo_U_dcore_U_sub_fifo_n297;
   wire FE_PHN5058_U_afifo_U_acore_U_sub_fifo_n205;
   wire FE_PHN5057_U_dfifo_U_dcore_U_sub_fifo_n285;
   wire FE_PHN5054_U_dfifo_U_dcore_n153;
   wire FE_PHN5051_U_dfifo_U_dcore_U_sub_fifo_n254;
   wire FE_PHN5048_U_afifo_U_acore_U_sub_fifo_n255;
   wire FE_PHN5041_U_dfifo_U_dcore_U_sub_fifo_n178;
   wire FE_PHN5040_U_afifo_U_acore_U_sub_fifo_n237;
   wire FE_PHN5038_U_afifo_U_acore_U_sub_fifo_n274;
   wire FE_PHN5037_U_afifo_U_acore_U_sub_fifo_n315;
   wire FE_PHN5036_U_dfifo_U_dcore_U_sub_fifo_n255;
   wire FE_PHN5033_U_dfifo_U_dcore_U_sub_fifo_n281;
   wire FE_PHN5032_U_afifo_U_acore_U_sub_fifo_n192;
   wire FE_PHN5030_U_dfifo_U_dcore_U_sub_fifo_n304;
   wire FE_PHN5024_U_afifo_n17;
   wire FE_PHN5022_U_afifo_U_acore_U_sub_fifo_n191;
   wire FE_PHN5021_U_afifo_n166;
   wire FE_PHN5020_U_afifo_U_acore_U_sub_fifo_n184;
   wire FE_PHN5016_U_dfifo_U_dcore_n156;
   wire FE_PHN5009_U_afifo_U_acore_U_sub_fifo_n273;
   wire FE_PHN5007_U_afifo_U_acore_U_sub_fifo_n285;
   wire FE_PHN5005_U_afifo_U_acore_U_sub_fifo_n187;
   wire FE_PHN5004_U_afifo_n165;
   wire FE_PHN5003_U_afifo_U_acore_U_sub_fifo_n283;
   wire FE_PHN4998_U_dfifo_U_dcore_U_sub_fifo_n302;
   wire FE_PHN4996_U_afifo_U_acore_U_sub_fifo_n202;
   wire FE_PHN4993_U_dfifo_U_dcore_U_sub_fifo_n279;
   wire FE_PHN4992_U_afifo_U_acore_U_sub_fifo_n235;
   wire FE_PHN4987_U_afifo_U_acore_U_sub_fifo_n210;
   wire FE_PHN4981_U_afifo_U_acore_U_sub_fifo_n277;
   wire FE_PHN4979_U_afifo_U_acore_U_sub_fifo_n173;
   wire FE_PHN4978_U_afifo_U_acore_U_sub_fifo_n247;
   wire FE_PHN4975_U_dfifo_U_dcore_U_sub_fifo_n213;
   wire FE_PHN4973_U_afifo_U_acore_U_sub_fifo_n218;
   wire FE_PHN4968_U_dfifo_U_dcore_U_sub_fifo_n266;
   wire FE_PHN4965_U_afifo_U_acore_U_sub_fifo_n203;
   wire FE_PHN4964_U_afifo_U_acore_U_sub_fifo_n240;
   wire FE_PHN4961_U_dfifo_U_dcore_U_sub_fifo_n291;
   wire FE_PHN4957_U_afifo_n192;
   wire FE_PHN4951_U_afifo_U_acore_U_sub_fifo_n229;
   wire FE_PHN4948_U_dfifo_U_dcore_U_sub_fifo_n261;
   wire FE_PHN4945_U_dfifo_U_dcore_n151;
   wire FE_PHN4942_U_afifo_U_acore_U_sub_fifo_n258;
   wire FE_PHN4939_U_dfifo_U_dcore_U_sub_fifo_n253;
   wire FE_PHN4936_U_afifo_U_acore_U_sub_fifo_n222;
   wire FE_PHN4929_U_dfifo_U_dcore_U_sub_fifo_n210;
   wire FE_PHN4928_U_dfifo_U_dcore_n157;
   wire FE_PHN4926_U_dfifo_U_dcore_n154;
   wire FE_PHN4925_U_dfifo_U_dcore_U_sub_fifo_n267;
   wire FE_PHN4918_U_dfifo_U_dcore_U_sub_fifo_n296;
   wire FE_PHN4917_U_afifo_n191;
   wire FE_PHN4908_U_dfifo_U_dcore_U_sub_fifo_n216;
   wire FE_PHN4903_U_dfifo_U_dcore_U_sub_fifo_n164;
   wire FE_PHN4901_U_dfifo_U_dcore_n155;
   wire FE_PHN4899_U_afifo_U_acore_U_sub_fifo_n256;
   wire FE_PHN4892_U_dfifo_U_dcore_U_sub_fifo_n202;
   wire FE_PHN4889_U_dfifo_U_dcore_U_sub_fifo_n314;
   wire FE_PHN4881_U_dfifo_U_dcore_U_sub_fifo_n256;
   wire FE_PHN4880_U_dfifo_U_dcore_U_sub_fifo_n174;
   wire FE_PHN4879_U_dfifo_U_dcore_U_sub_fifo_n176;
   wire FE_PHN4877_U_afifo_U_acore_U_sub_fifo_n320;
   wire FE_PHN4875_U_dfifo_U_dcore_U_sub_fifo_n172;
   wire FE_PHN4872_U_dfifo_U_dcore_U_sub_fifo_n163;
   wire FE_PHN4858_U_afifo_U_acore_U_sub_fifo_n214;
   wire FE_PHN4856_U_dfifo_U_dcore_U_sub_fifo_n413;
   wire FE_PHN4852_U_dfifo_U_dcore_U_sub_fifo_n207;
   wire FE_PHN4848_U_dfifo_U_dcore_U_sub_fifo_n179;
   wire FE_PHN4846_U_dfifo_U_dcore_U_sub_fifo_n166;
   wire FE_PHN4843_U_dfifo_U_dcore_U_sub_fifo_n298;
   wire FE_PHN4837_U_dfifo_U_dcore_U_sub_fifo_n214;
   wire FE_PHN4836_U_dfifo_U_dcore_U_sub_fifo_n212;
   wire FE_PHN4832_U_dfifo_U_dcore_U_sub_fifo_n338;
   wire FE_PHN4826_U_dfifo_U_dcore_U_sub_fifo_n169;
   wire FE_PHN4825_U_dfifo_U_dcore_U_sub_fifo_n168;
   wire FE_PHN4824_U_dfifo_U_dcore_U_sub_fifo_n445;
   wire FE_PHN4819_U_afifo_U_acore_U_sub_fifo_n267;
   wire FE_PHN4817_U_dfifo_U_dcore_U_sub_fifo_n218;
   wire FE_PHN4816_U_dfifo_U_dcore_U_sub_fifo_n209;
   wire FE_PHN4812_U_dfifo_U_dcore_U_sub_fifo_n450;
   wire FE_PHN4811_U_dfifo_U_dcore_U_sub_fifo_n165;
   wire FE_PHN4806_U_dfifo_U_dcore_U_sub_fifo_n401;
   wire FE_PHN4803_U_dfifo_U_dcore_U_sub_fifo_n170;
   wire FE_PHN4800_U_dfifo_U_dcore_U_sub_fifo_n173;
   wire FE_PHN4799_U_dfifo_U_dcore_U_sub_fifo_n175;
   wire FE_PHN4793_U_afifo_U_acore_U_sub_fifo_n266;
   wire FE_PHN4791_U_dfifo_U_dcore_U_sub_fifo_n205;
   wire FE_PHN4789_U_afifo_U_acore_U_sub_fifo_n296;
   wire FE_PHN4786_U_dfifo_U_dcore_U_sub_fifo_n211;
   wire FE_PHN4780_U_dfifo_U_dcore_n145;
   wire FE_PHN4773_U_dfifo_U_dcore_U_sub_fifo_n215;
   wire FE_PHN4771_U_dfifo_U_dcore_U_sub_fifo_n219;
   wire FE_PHN4770_U_dfifo_U_dcore_U_sub_fifo_n344;
   wire FE_PHN4769_U_dfifo_U_dcore_U_sub_fifo_n333;
   wire FE_PHN4768_U_dfifo_U_dcore_U_sub_fifo_n403;
   wire FE_PHN4766_U_dfifo_U_dcore_U_sub_fifo_n397;
   wire FE_PHN4765_U_dfifo_U_dcore_U_sub_fifo_n398;
   wire FE_PHN4764_U_dfifo_U_dcore_U_sub_fifo_n208;
   wire FE_PHN4762_U_dfifo_U_dcore_U_sub_fifo_n220;
   wire FE_PHN4758_U_afifo_U_acore_U_sub_fifo_n269;
   wire FE_PHN4757_U_dfifo_U_dcore_U_sub_fifo_n206;
   wire FE_PHN4755_U_dfifo_U_dcore_U_sub_fifo_n442;
   wire FE_PHN4754_U_dfifo_U_dcore_U_sub_fifo_n356;
   wire FE_PHN4753_U_dfifo_U_dcore_U_sub_fifo_n167;
   wire FE_PHN4752_U_dfifo_U_dcore_U_sub_fifo_n440;
   wire FE_PHN4751_U_dfifo_U_dcore_U_sub_fifo_n327;
   wire FE_PHN4747_U_dfifo_U_dcore_U_sub_fifo_n412;
   wire FE_PHN4746_U_dfifo_U_dcore_U_sub_fifo_n320;
   wire FE_PHN4745_U_dfifo_U_dcore_U_sub_fifo_n452;
   wire FE_PHN4744_U_dfifo_U_dcore_U_sub_fifo_n402;
   wire FE_PHN4742_U_dfifo_U_dcore_U_sub_fifo_n316;
   wire FE_PHN4741_U_dfifo_U_dcore_U_sub_fifo_n204;
   wire FE_PHN4740_U_dfifo_U_dcore_U_sub_fifo_n340;
   wire FE_PHN4738_U_dfifo_U_dcore_U_sub_fifo_n446;
   wire FE_PHN4719_U_afifo_U_acore_n97;
   wire FE_PHN4705_U_ctl_N89;
   wire FE_PHN4677_U_afifo_U_acore_U_sub_fifo_n297;
   wire FE_PHN4665_U_rbuf_n69;
   wire FE_PHN4664_miu_data_27_;
   wire FE_PHN4663_U_rbuf_n175;
   wire FE_PHN4650_U_rbuf_n63;
   wire FE_PHN4649_U_rbuf_n59;
   wire FE_PHN4647_U_rbuf_n174;
   wire FE_PHN4646_U_rbuf_n179;
   wire FE_PHN4644_U_rbuf_n182;
   wire FE_PHN4643_U_rbuf_n56;
   wire FE_PHN4642_U_rbuf_n75;
   wire FE_PHN4640_U_ctl_n_bh_state_0_;
   wire FE_PHN4636_hsel_reg;
   wire FE_PHN4635_U_rbuf_n188;
   wire FE_PHN4633_U_ctl_n212;
   wire FE_PHN4632_U_ctl_n_sel_buf;
   wire FE_PHN4628_U_ctl_n382;
   wire FE_PHN4626_m_af_push1_n;
   wire FE_PHN4619_U_ctl_f_burst_done;
   wire FE_PHN4384_U_dfifo_U_dcore_n_empty;
   wire FE_PHN4370_U_dfifo_U_dcore_U_sub_fifo_n272;
   wire FE_PHN4347_U_dfifo_U_dcore_U_sub_fifo_n303;
   wire FE_PHN4341_U_dfifo_U_dcore_U_sub_fifo_n262;
   wire FE_PHN4321_U_dfifo_U_dcore_U_sub_fifo_n55;
   wire FE_PHN4310_U_dfifo_U_dcore_U_sub_fifo_n258;
   wire FE_PHN4309_U_dfifo_U_dcore_U_sub_fifo_n278;
   wire FE_PHN4300_U_dfifo_U_dcore_U_sub_fifo_n306;
   wire FE_PHN4299_U_dfifo_U_dcore_U_sub_fifo_n451;
   wire FE_PHN4296_U_dfifo_U_dcore_U_sub_fifo_n276;
   wire FE_PHN4294_U_dfifo_U_dcore_U_sub_fifo_n448;
   wire FE_PHN4292_U_dfifo_U_dcore_U_sub_fifo_n271;
   wire FE_PHN4290_U_dfifo_U_dcore_U_sub_fifo_n270;
   wire FE_PHN4285_U_dfifo_U_dcore_U_sub_fifo_n294;
   wire FE_PHN4284_U_dfifo_U_dcore_U_sub_fifo_n260;
   wire FE_PHN4281_U_dfifo_U_dcore_U_sub_fifo_n264;
   wire FE_PHN4278_U_dfifo_U_dcore_U_sub_fifo_n265;
   wire FE_PHN4276_U_dfifo_U_dcore_U_sub_fifo_n283;
   wire FE_PHN4275_U_dfifo_U_dcore_U_sub_fifo_n295;
   wire FE_PHN4268_U_dfifo_U_dcore_U_sub_fifo_n277;
   wire FE_PHN4256_U_dfifo_U_dcore_U_sub_fifo_n243;
   wire FE_PHN4255_U_dfifo_U_dcore_U_sub_fifo_n259;
   wire FE_PHN4254_U_dfifo_U_dcore_U_sub_fifo_n282;
   wire FE_PHN4253_U_dfifo_U_dcore_U_sub_fifo_n268;
   wire FE_PHN4252_U_dfifo_U_dcore_U_sub_fifo_n309;
   wire FE_PHN4251_U_dfifo_U_dcore_U_sub_fifo_n250;
   wire FE_PHN4250_U_dfifo_U_dcore_U_sub_fifo_n248;
   wire FE_PHN4245_U_dfifo_U_dcore_U_sub_fifo_n269;
   wire FE_PHN4244_U_dfifo_U_dcore_U_sub_fifo_n299;
   wire FE_PHN4243_U_dfifo_U_dcore_U_sub_fifo_n305;
   wire FE_PHN4242_U_dfifo_U_dcore_U_sub_fifo_n300;
   wire FE_PHN4241_U_dfifo_U_dcore_U_sub_fifo_n286;
   wire FE_PHN4239_U_dfifo_U_dcore_U_sub_fifo_n273;
   wire FE_PHN4238_U_dfifo_U_dcore_U_sub_fifo_n284;
   wire FE_PHN4236_U_dfifo_U_dcore_U_sub_fifo_n257;
   wire FE_PHN4228_U_dfifo_U_dcore_U_sub_fifo_n254;
   wire FE_PHN4226_U_afifo_U_acore_U_sub_fifo_n279;
   wire FE_PHN4225_U_dfifo_U_dcore_U_sub_fifo_n310;
   wire FE_PHN4224_U_dfifo_U_dcore_U_sub_fifo_n293;
   wire FE_PHN4223_U_afifo_U_acore_U_sub_fifo_n309;
   wire FE_PHN4222_U_dfifo_U_dcore_U_sub_fifo_n274;
   wire FE_PHN4211_U_dfifo_U_dcore_U_sub_fifo_n292;
   wire FE_PHN4210_U_dfifo_U_dcore_U_sub_fifo_n255;
   wire FE_PHN4209_U_dfifo_U_dcore_U_sub_fifo_n288;
   wire FE_PHN4208_U_dfifo_U_dcore_U_sub_fifo_n245;
   wire FE_PHN4207_U_dfifo_U_dcore_n156;
   wire FE_PHN4206_U_dfifo_U_dcore_U_sub_fifo_n290;
   wire FE_PHN4203_U_afifo_U_acore_U_sub_fifo_n196;
   wire FE_PHN4197_U_afifo_U_acore_U_sub_fifo_n208;
   wire FE_PHN4195_U_dfifo_U_dcore_U_sub_fifo_n308;
   wire FE_PHN4194_U_dfifo_U_dcore_U_sub_fifo_n307;
   wire FE_PHN4190_U_dfifo_U_dcore_U_sub_fifo_n285;
   wire FE_PHN4189_U_dfifo_U_dcore_U_sub_fifo_n249;
   wire FE_PHN4188_U_dfifo_U_dcore_U_sub_fifo_n280;
   wire FE_PHN4186_U_afifo_n159;
   wire FE_PHN4184_U_dfifo_U_dcore_U_sub_fifo_n247;
   wire FE_PHN4183_U_dfifo_U_dcore_U_sub_fifo_n246;
   wire FE_PHN4179_U_afifo_U_acore_U_sub_fifo_n192;
   wire FE_PHN4173_U_dfifo_U_dcore_U_sub_fifo_n251;
   wire FE_PHN4164_U_afifo_U_acore_U_sub_fifo_n275;
   wire FE_PHN4163_U_afifo_U_acore_U_sub_fifo_n205;
   wire FE_PHN4162_U_dfifo_U_dcore_n154;
   wire FE_PHN4159_U_afifo_U_acore_U_sub_fifo_n187;
   wire FE_PHN4158_U_afifo_U_acore_U_sub_fifo_n191;
   wire FE_PHN4157_U_dfifo_U_dcore_U_sub_fifo_n275;
   wire FE_PHN4156_U_dfifo_U_dcore_U_sub_fifo_n291;
   wire FE_PHN4155_U_dfifo_U_dcore_n153;
   wire FE_PHN4153_U_afifo_U_acore_U_sub_fifo_n184;
   wire FE_PHN4151_U_dfifo_U_dcore_U_sub_fifo_n304;
   wire FE_PHN4144_U_dfifo_U_dcore_U_sub_fifo_n267;
   wire FE_PHN4143_U_dfifo_U_dcore_U_sub_fifo_n279;
   wire FE_PHN4137_U_dfifo_U_dcore_U_sub_fifo_n253;
   wire FE_PHN4134_U_afifo_U_acore_U_sub_fifo_n210;
   wire FE_PHN4131_U_dfifo_U_dcore_U_sub_fifo_n296;
   wire FE_PHN4130_U_dfifo_U_dcore_U_sub_fifo_n281;
   wire FE_PHN4128_U_afifo_U_acore_U_sub_fifo_n188;
   wire FE_PHN4127_U_afifo_U_acore_U_sub_fifo_n291;
   wire FE_PHN4125_U_dfifo_U_dcore_U_sub_fifo_n263;
   wire FE_PHN4121_U_afifo_U_acore_U_sub_fifo_n265;
   wire FE_PHN4116_U_dfifo_U_dcore_U_sub_fifo_n261;
   wire FE_PHN4114_U_afifo_U_acore_U_sub_fifo_n218;
   wire FE_PHN4113_U_afifo_U_acore_U_sub_fifo_n314;
   wire FE_PHN4112_U_afifo_U_acore_U_sub_fifo_n317;
   wire FE_PHN4111_U_afifo_U_acore_U_sub_fifo_n180;
   wire FE_PHN4107_U_afifo_U_acore_U_sub_fifo_n190;
   wire FE_PHN4106_U_afifo_U_acore_U_sub_fifo_n285;
   wire FE_PHN4105_U_afifo_n17;
   wire FE_PHN4103_U_dfifo_U_dcore_U_sub_fifo_n266;
   wire FE_PHN4100_U_afifo_U_acore_U_sub_fifo_n263;
   wire FE_PHN4099_U_afifo_U_acore_U_sub_fifo_n264;
   wire FE_PHN4098_U_afifo_U_acore_U_sub_fifo_n283;
   wire FE_PHN4097_U_afifo_U_acore_U_sub_fifo_n284;
   wire FE_PHN4095_U_dfifo_U_dcore_U_sub_fifo_n287;
   wire FE_PHN4092_U_afifo_U_acore_U_sub_fifo_n288;
   wire FE_PHN4091_U_dfifo_U_dcore_U_sub_fifo_n289;
   wire FE_PHN4087_U_afifo_U_acore_U_sub_fifo_n214;
   wire FE_PHN4086_U_afifo_n191;
   wire FE_PHN4081_U_afifo_U_acore_U_sub_fifo_n213;
   wire FE_PHN4080_U_afifo_U_acore_U_sub_fifo_n230;
   wire FE_PHN4079_U_afifo_n166;
   wire FE_PHN4074_U_afifo_U_acore_U_sub_fifo_n232;
   wire FE_PHN4073_U_dfifo_U_dcore_U_sub_fifo_n297;
   wire FE_PHN4071_U_afifo_U_acore_U_sub_fifo_n224;
   wire FE_PHN4070_U_afifo_U_acore_U_sub_fifo_n181;
   wire FE_PHN4069_U_afifo_U_acore_U_sub_fifo_n315;
   wire FE_PHN4068_U_dfifo_U_dcore_U_sub_fifo_n301;
   wire FE_PHN4066_U_afifo_U_acore_U_sub_fifo_n178;
   wire FE_PHN4065_U_afifo_U_acore_U_sub_fifo_n175;
   wire FE_PHN4064_U_dfifo_U_dcore_U_sub_fifo_n179;
   wire FE_PHN4063_U_dfifo_U_dcore_U_sub_fifo_n244;
   wire FE_PHN4062_U_dfifo_U_dcore_U_sub_fifo_n256;
   wire FE_PHN4056_U_afifo_U_acore_U_sub_fifo_n215;
   wire FE_PHN4055_U_afifo_U_acore_U_sub_fifo_n290;
   wire FE_PHN4049_U_afifo_U_acore_U_sub_fifo_n247;
   wire FE_PHN4046_U_dfifo_U_dcore_n150;
   wire FE_PHN4038_U_afifo_U_acore_U_sub_fifo_n259;
   wire FE_PHN4037_U_afifo_U_acore_U_sub_fifo_n320;
   wire FE_PHN4036_U_afifo_U_acore_U_sub_fifo_n197;
   wire FE_PHN4033_U_dfifo_U_dcore_U_sub_fifo_n302;
   wire FE_PHN4030_U_afifo_U_acore_U_sub_fifo_n257;
   wire FE_PHN4028_U_afifo_n192;
   wire FE_PHN4025_U_afifo_n165;
   wire FE_PHN4019_U_afifo_U_acore_U_sub_fifo_n304;
   wire FE_PHN4016_U_afifo_U_acore_U_sub_fifo_n211;
   wire FE_PHN4015_U_afifo_U_acore_U_sub_fifo_n183;
   wire FE_PHN4014_U_afifo_U_acore_U_sub_fifo_n207;
   wire FE_PHN4011_U_afifo_U_acore_U_sub_fifo_n195;
   wire FE_PHN4010_U_afifo_U_acore_U_sub_fifo_n182;
   wire FE_PHN4009_U_afifo_U_acore_U_sub_fifo_n242;
   wire FE_PHN4008_U_dfifo_U_dcore_U_sub_fifo_n298;
   wire FE_PHN4007_U_dfifo_U_dcore_U_sub_fifo_n252;
   wire FE_PHN3999_U_afifo_U_acore_U_sub_fifo_n261;
   wire FE_PHN3998_U_afifo_U_acore_U_sub_fifo_n174;
   wire FE_PHN3997_U_afifo_U_acore_U_sub_fifo_n179;
   wire FE_PHN3996_U_afifo_U_acore_U_sub_fifo_n204;
   wire FE_PHN3995_U_afifo_U_acore_U_sub_fifo_n238;
   wire FE_PHN3994_U_afifo_U_acore_U_sub_fifo_n229;
   wire FE_PHN3993_U_afifo_U_acore_U_sub_fifo_n254;
   wire FE_PHN3992_U_afifo_U_acore_U_sub_fifo_n240;
   wire FE_PHN3991_U_afifo_U_acore_U_sub_fifo_n189;
   wire FE_PHN3990_U_afifo_U_acore_U_sub_fifo_n222;
   wire FE_PHN3984_U_afifo_U_acore_U_sub_fifo_n216;
   wire FE_PHN3980_U_afifo_U_acore_U_sub_fifo_n289;
   wire FE_PHN3979_U_afifo_U_acore_U_sub_fifo_n258;
   wire FE_PHN3978_U_afifo_U_acore_U_sub_fifo_n244;
   wire FE_PHN3967_U_afifo_U_acore_U_sub_fifo_n245;
   wire FE_PHN3966_U_afifo_U_acore_U_sub_fifo_n228;
   wire FE_PHN3965_U_dfifo_U_dcore_n152;
   wire FE_PHN3964_U_dfifo_U_dcore_U_sub_fifo_n205;
   wire FE_PHN3957_U_afifo_U_acore_U_sub_fifo_n186;
   wire FE_PHN3956_U_afifo_U_acore_U_sub_fifo_n233;
   wire FE_PHN3955_U_afifo_U_acore_U_sub_fifo_n281;
   wire FE_PHN3953_U_afifo_U_acore_U_sub_fifo_n234;
   wire FE_PHN3952_U_afifo_U_acore_U_sub_fifo_n286;
   wire FE_PHN3947_U_afifo_U_acore_U_sub_fifo_n194;
   wire FE_PHN3946_U_afifo_U_acore_U_sub_fifo_n282;
   wire FE_PHN3945_U_afifo_U_acore_U_sub_fifo_n225;
   wire FE_PHN3944_U_dfifo_U_dcore_U_sub_fifo_n171;
   wire FE_PHN3940_U_afifo_U_acore_U_sub_fifo_n239;
   wire FE_PHN3939_U_afifo_U_acore_U_sub_fifo_n209;
   wire FE_PHN3936_U_afifo_U_acore_U_sub_fifo_n231;
   wire FE_PHN3935_U_afifo_U_acore_U_sub_fifo_n220;
   wire FE_PHN3933_U_dfifo_U_dcore_U_sub_fifo_n210;
   wire FE_PHN3932_U_dfifo_U_dcore_U_sub_fifo_n170;
   wire FE_PHN3929_U_afifo_U_acore_U_sub_fifo_n241;
   wire FE_PHN3920_U_afifo_U_acore_U_sub_fifo_n260;
   wire FE_PHN3914_U_afifo_U_acore_U_sub_fifo_n217;
   wire FE_PHN3913_U_dfifo_U_dcore_U_sub_fifo_n164;
   wire FE_PHN3905_U_afifo_U_acore_U_sub_fifo_n237;
   wire FE_PHN3901_U_afifo_U_acore_U_sub_fifo_n236;
   wire FE_PHN3899_U_dfifo_U_dcore_U_sub_fifo_n213;
   wire FE_PHN3897_U_afifo_n158;
   wire FE_PHN3895_U_afifo_U_acore_U_sub_fifo_n235;
   wire FE_PHN3894_U_dfifo_U_dcore_U_sub_fifo_n216;
   wire FE_PHN3891_U_afifo_U_acore_U_sub_fifo_n185;
   wire FE_PHN3890_U_afifo_U_acore_U_sub_fifo_n255;
   wire FE_PHN3881_U_afifo_U_acore_U_sub_fifo_n246;
   wire FE_PHN3873_U_dfifo_U_dcore_n151;
   wire FE_PHN3861_U_dfifo_U_dcore_U_sub_fifo_n214;
   wire FE_PHN3860_U_dfifo_U_dcore_U_sub_fifo_n218;
   wire FE_PHN3859_U_dfifo_U_dcore_U_sub_fifo_n163;
   wire FE_PHN3858_U_dfifo_U_dcore_U_sub_fifo_n209;
   wire FE_PHN3855_U_dfifo_U_dcore_U_sub_fifo_n215;
   wire FE_PHN3854_U_dfifo_U_dcore_U_sub_fifo_n219;
   wire FE_PHN3852_U_dfifo_U_dcore_U_sub_fifo_n202;
   wire FE_PHN3850_U_dfifo_U_dcore_U_sub_fifo_n178;
   wire FE_PHN3849_U_dfifo_U_dcore_U_sub_fifo_n175;
   wire FE_PHN3848_U_dfifo_U_dcore_U_sub_fifo_n166;
   wire FE_PHN3846_U_dfifo_U_dcore_U_sub_fifo_n211;
   wire FE_PHN3841_U_dfifo_U_dcore_U_sub_fifo_n207;
   wire FE_PHN3840_U_dfifo_U_dcore_U_sub_fifo_n314;
   wire FE_PHN3838_U_dfifo_U_dcore_U_sub_fifo_n177;
   wire FE_PHN3837_U_afifo_U_acore_U_sub_fifo_n268;
   wire FE_PHN3835_U_dfifo_U_dcore_U_sub_fifo_n169;
   wire FE_PHN3834_U_dfifo_U_dcore_U_sub_fifo_n206;
   wire FE_PHN3832_U_dfifo_U_dcore_U_sub_fifo_n174;
   wire FE_PHN3829_U_dfifo_U_dcore_U_sub_fifo_n337;
   wire FE_PHN3827_U_dfifo_U_dcore_U_sub_fifo_n162;
   wire FE_PHN3825_U_dfifo_U_dcore_U_sub_fifo_n445;
   wire FE_PHN3824_U_dfifo_U_dcore_U_sub_fifo_n168;
   wire FE_PHN3822_U_dfifo_U_dcore_U_sub_fifo_n413;
   wire FE_PHN3820_U_dfifo_U_dcore_U_sub_fifo_n220;
   wire FE_PHN3819_U_dfifo_U_dcore_U_sub_fifo_n165;
   wire FE_PHN3818_U_dfifo_U_dcore_U_sub_fifo_n173;
   wire FE_PHN3817_U_afifo_U_acore_U_sub_fifo_n267;
   wire FE_PHN3815_U_dfifo_U_dcore_U_sub_fifo_n212;
   wire FE_PHN3813_U_afifo_U_acore_U_sub_fifo_n272;
   wire FE_PHN3812_U_dfifo_U_dcore_U_sub_fifo_n176;
   wire FE_PHN3809_U_dfifo_U_dcore_U_sub_fifo_n329;
   wire FE_PHN3807_U_dfifo_U_dcore_U_sub_fifo_n172;
   wire FE_PHN3805_U_dfifo_U_dcore_U_sub_fifo_n204;
   wire FE_PHN3804_U_dfifo_U_dcore_U_sub_fifo_n330;
   wire FE_PHN3801_U_dfifo_U_dcore_U_sub_fifo_n415;
   wire FE_PHN3795_U_afifo_U_acore_U_sub_fifo_n266;
   wire FE_PHN3794_U_dfifo_U_dcore_U_sub_fifo_n321;
   wire FE_PHN3792_U_dfifo_U_dcore_U_sub_fifo_n217;
   wire FE_PHN3791_U_dfifo_U_dcore_U_sub_fifo_n401;
   wire FE_PHN3790_U_dfifo_U_dcore_U_sub_fifo_n338;
   wire FE_PHN3789_U_dfifo_U_dcore_n144;
   wire FE_PHN3788_U_dfifo_U_dcore_U_sub_fifo_n317;
   wire FE_PHN3783_U_dfifo_U_dcore_U_sub_fifo_n333;
   wire FE_PHN3772_U_afifo_U_acore_U_sub_fifo_n270;
   wire FE_PHN3770_U_afifo_n20;
   wire FE_PHN3767_U_dfifo_U_dcore_U_sub_fifo_n344;
   wire FE_PHN3761_U_dfifo_U_dcore_U_sub_fifo_n203;
   wire FE_PHN3756_U_dfifo_U_dcore_n143;
   wire FE_PHN3754_U_dfifo_U_dcore_U_sub_fifo_n315;
   wire FE_PHN3752_U_dfifo_U_dcore_U_sub_fifo_n416;
   wire FE_PHN3750_U_dfifo_U_dcore_U_sub_fifo_n407;
   wire FE_PHN3749_U_dfifo_U_dcore_U_sub_fifo_n167;
   wire FE_PHN3748_U_dfifo_U_dcore_U_sub_fifo_n313;
   wire FE_PHN3747_U_dfifo_U_dcore_U_sub_fifo_n403;
   wire FE_PHN3746_U_dfifo_U_dcore_U_sub_fifo_n397;
   wire FE_PHN3743_U_dfifo_U_dcore_U_sub_fifo_n417;
   wire FE_PHN3742_U_dfifo_U_dcore_U_sub_fifo_n324;
   wire FE_PHN3741_U_dfifo_U_dcore_U_sub_fifo_n325;
   wire FE_PHN3740_U_dfifo_U_dcore_U_sub_fifo_n398;
   wire FE_PHN3734_U_dfifo_U_dcore_U_sub_fifo_n208;
   wire FE_PHN3732_U_dfifo_U_dcore_U_sub_fifo_n326;
   wire FE_PHN3731_U_dfifo_U_dcore_U_sub_fifo_n442;
   wire FE_PHN3729_U_dfifo_U_dcore_U_sub_fifo_n356;
   wire FE_PHN3728_U_dfifo_U_dcore_U_sub_fifo_n318;
   wire FE_PHN3727_U_dfifo_U_dcore_U_sub_fifo_n443;
   wire FE_PHN3723_U_dfifo_U_dcore_U_sub_fifo_n340;
   wire FE_PHN3721_U_dfifo_U_dcore_U_sub_fifo_n411;
   wire FE_PHN3720_U_dfifo_U_dcore_U_sub_fifo_n402;
   wire FE_PHN3719_U_dfifo_U_dcore_U_sub_fifo_n440;
   wire FE_PHN3716_U_dfifo_U_dcore_n147;
   wire FE_PHN3715_U_dfifo_U_dcore_U_sub_fifo_n127;
   wire FE_PHN3711_U_dfifo_U_dcore_U_sub_fifo_n405;
   wire FE_PHN3710_U_dfifo_U_dcore_U_sub_fifo_n406;
   wire FE_PHN3709_U_dfifo_U_dcore_U_sub_fifo_n412;
   wire FE_PHN3708_U_dfifo_U_dcore_U_sub_fifo_n327;
   wire FE_PHN3706_U_dfifo_U_dcore_U_sub_fifo_n399;
   wire FE_PHN3705_U_dfifo_U_dcore_U_sub_fifo_n339;
   wire FE_PHN3703_U_dfifo_U_dcore_U_sub_fifo_n414;
   wire FE_PHN3701_U_dfifo_U_dcore_U_sub_fifo_n400;
   wire FE_PHN3700_U_dfifo_U_dcore_U_sub_fifo_n320;
   wire FE_PHN3696_U_dfifo_U_dcore_U_sub_fifo_n323;
   wire FE_PHN3695_U_dfifo_U_dcore_U_sub_fifo_n311;
   wire FE_PHN3694_U_dfifo_U_dcore_U_sub_fifo_n404;
   wire FE_PHN3693_U_dfifo_U_dcore_U_sub_fifo_n331;
   wire FE_PHN3691_U_dfifo_U_dcore_U_sub_fifo_n334;
   wire FE_PHN3689_U_dfifo_U_dcore_U_sub_fifo_n441;
   wire FE_PHN3688_U_dfifo_U_dcore_U_sub_fifo_n439;
   wire FE_PHN3685_U_dfifo_U_dcore_U_sub_fifo_n418;
   wire FE_PHN3679_U_dfifo_U_dcore_U_sub_fifo_n343;
   wire FE_PHN3678_U_dfifo_U_dcore_U_sub_fifo_n319;
   wire FE_PHN3677_U_dfifo_U_dcore_U_sub_fifo_n332;
   wire FE_PHN3676_U_dfifo_U_dcore_U_sub_fifo_n444;
   wire FE_PHN3675_U_dfifo_U_dcore_U_sub_fifo_n438;
   wire FE_PHN3674_U_dfifo_U_dcore_U_sub_fifo_n322;
   wire FE_PHN3673_U_dfifo_U_dcore_U_sub_fifo_n446;
   wire FE_PHN3671_U_afifo_n18;
   wire FE_PHN3670_U_dfifo_U_dcore_U_sub_fifo_n328;
   wire FE_PHN3668_U_dfifo_U_dcore_U_sub_fifo_n341;
   wire FE_PHN3667_U_dfifo_U_dcore_U_sub_fifo_n408;
   wire FE_PHN3664_U_dfifo_U_dcore_U_sub_fifo_n410;
   wire FE_PHN3658_U_dfifo_U_dcore_U_sub_fifo_n409;
   wire FE_PHN3656_U_dfifo_U_dcore_U_sub_fifo_n335;
   wire FE_PHN3655_U_dfifo_U_dcore_n146;
   wire FE_PHN3652_U_dfifo_U_dcore_U_sub_fifo_n312;
   wire FE_PHN3650_U_dfifo_U_dcore_U_sub_fifo_n342;
   wire FE_PHN3649_U_dfifo_U_dcore_U_sub_fifo_n336;
   wire FE_PHN3646_U_afifo_n19;
   wire FE_PHN3644_U_dfifo_U_dcore_U_sub_fifo_n316;
   wire FE_PHN3632_U_dfifo_U_dcore_n13;
   wire FE_PHN3618_U_dfifo_U_dcore_n14;
   wire FE_PHN3543_U_afifo_n164;
   wire FE_PHN3504_U_afifo_U_acore_U_sub_fifo_n223;
   wire FE_PHN3499_U_afifo_U_acore_U_sub_fifo_n248;
   wire FE_PHN3498_U_afifo_U_acore_U_sub_fifo_n250;
   wire FE_PHN3495_U_afifo_U_acore_U_sub_fifo_n173;
   wire FE_PHN3494_U_afifo_U_acore_U_sub_fifo_n219;
   wire FE_PHN3493_U_afifo_U_acore_U_sub_fifo_n253;
   wire FE_PHN3492_U_afifo_U_acore_U_sub_fifo_n226;
   wire FE_PHN3491_U_afifo_U_acore_U_sub_fifo_n177;
   wire FE_PHN3490_U_afifo_U_acore_U_sub_fifo_n227;
   wire FE_PHN3489_U_afifo_U_acore_U_sub_fifo_n256;
   wire FE_PHN3488_U_afifo_U_acore_U_sub_fifo_n252;
   wire FE_PHN3487_U_afifo_U_acore_U_sub_fifo_n199;
   wire FE_PHN3486_U_afifo_U_acore_U_sub_fifo_n193;
   wire FE_PHN3484_U_afifo_U_acore_U_sub_fifo_n251;
   wire FE_PHN3483_U_afifo_U_acore_U_sub_fifo_n243;
   wire FE_PHN3481_U_afifo_n157;
   wire FE_PHN3471_U_afifo_m_data_in_49_;
   wire FE_PHN3469_U_ctl_n136;
   wire FE_PHN3468_U_ctl_n103;
   wire FE_PHN3465_U_afifo_U_acore_f_obuf_34_;
   wire FE_PHN3462_U_ctl_n101;
   wire FE_PHN3460_U_afifo_U_acore_n157;
   wire FE_PHN3459_U_afifo_U_acore_n91;
   wire FE_PHN3458_U_afifo_n186;
   wire FE_PHN3457_U_afifo_U_acore_n69;
   wire FE_PHN3455_U_afifo_U_acore_n164;
   wire FE_PHN3453_U_afifo_U_acore_n75;
   wire FE_PHN3451_U_ctl_n102;
   wire FE_PHN3448_U_afifo_U_acore_n89;
   wire FE_PHN3447_U_afifo_U_acore_n101;
   wire FE_PHN3444_U_afifo_U_acore_n87;
   wire FE_PHN3441_U_afifo_n202;
   wire FE_PHN3439_U_afifo_n212;
   wire FE_PHN3438_U_dfifo_U_dcore_n200;
   wire FE_PHN3436_U_afifo_n208;
   wire FE_PHN3435_U_afifo_n198;
   wire FE_PHN3434_U_afifo_n210;
   wire FE_PHN3433_U_afifo_U_acore_n155;
   wire FE_PHN3430_U_afifo_U_acore_n143;
   wire FE_PHN3429_U_afifo_n220;
   wire FE_PHN3428_U_dfifo_U_dcore_n140;
   wire FE_PHN3426_U_afifo_U_acore_n_obuf_empty;
   wire FE_PHN3425_U_afifo_n188;
   wire FE_PHN3424_U_afifo_n232;
   wire FE_PHN3423_U_afifo_U_acore_n29;
   wire FE_PHN3422_U_afifo_n226;
   wire FE_PHN3420_U_afifo_n206;
   wire FE_PHN3419_U_afifo_n248;
   wire FE_PHN3418_U_afifo_n236;
   wire FE_PHN3417_U_dfifo_U_dcore_n194;
   wire FE_PHN3416_U_afifo_U_acore_n67;
   wire FE_PHN3413_U_afifo_n204;
   wire FE_PHN3412_U_afifo_U_acore_n158;
   wire FE_PHN3410_U_afifo_n230;
   wire FE_PHN3409_U_afifo_U_acore_n153;
   wire FE_PHN3408_U_afifo_n234;
   wire FE_PHN3406_U_afifo_U_acore_n99;
   wire FE_PHN3404_U_afifo_n218;
   wire FE_PHN3403_U_afifo_n224;
   wire FE_PHN3402_U_afifo_n238;
   wire FE_PHN3401_U_afifo_U_acore_n77;
   wire FE_PHN3400_U_afifo_n250;
   wire FE_PHN3398_U_dfifo_U_dcore_n195;
   wire FE_PHN3397_U_afifo_n200;
   wire FE_PHN3396_U_afifo_n240;
   wire FE_PHN3395_U_afifo_n244;
   wire FE_PHN3394_U_afifo_n246;
   wire FE_PHN3393_U_afifo_n216;
   wire FE_PHN3392_U_afifo_n222;
   wire FE_PHN3390_U_afifo_n173;
   wire FE_PHN3388_U_afifo_n214;
   wire FE_PHN3386_U_afifo_U_acore_n71;
   wire FE_PHN3385_U_afifo_n228;
   wire FE_PHN3384_U_afifo_U_acore_n156;
   wire FE_PHN3383_U_afifo_n242;
   wire FE_PHN3382_U_ctl_n105;
   wire FE_PHN3381_U_afifo_n171;
   wire FE_PHN3380_U_afifo_U_acore_n73;
   wire FE_PHN3376_U_afifo_U_acore_n200;
   wire FE_PHN3374_U_afifo_f_clr_pers;
   wire FE_PHN3372_U_dfifo_U_dcore_n178;
   wire FE_PHN3369_U_afifo_U_acore_n183;
   wire FE_PHN3368_U_dfifo_U_dcore_n192;
   wire FE_PHN3367_U_afifo_U_acore_n189;
   wire FE_PHN3366_U_afifo_U_acore_n180;
   wire FE_PHN3365_U_afifo_U_acore_n171;
   wire FE_PHN3364_U_dfifo_U_dcore_n180;
   wire FE_PHN3363_U_dfifo_U_dcore_n184;
   wire FE_PHN3362_U_afifo_U_acore_n193;
   wire FE_PHN3361_U_afifo_U_acore_n209;
   wire FE_PHN3360_U_afifo_U_acore_n182;
   wire FE_PHN3359_U_afifo_U_acore_n174;
   wire FE_PHN3358_U_dfifo_U_dcore_n176;
   wire FE_PHN3357_U_afifo_U_acore_f_afull;
   wire FE_PHN3356_U_afifo_U_acore_n187;
   wire FE_PHN3354_U_dfifo_U_dcore_n181;
   wire FE_PHN3351_U_dfifo_U_dcore_n193;
   wire FE_PHN3350_U_afifo_U_acore_n206;
   wire FE_PHN3348_U_afifo_U_acore_n202;
   wire FE_PHN3347_U_afifo_U_acore_n172;
   wire FE_PHN3344_U_afifo_U_acore_n191;
   wire FE_PHN3342_U_afifo_U_acore_n196;
   wire FE_PHN3341_U_dfifo_U_dcore_n189;
   wire FE_PHN3340_U_afifo_U_acore_n185;
   wire FE_PHN3339_U_dfifo_U_dcore_n182;
   wire FE_PHN3338_U_dfifo_U_dcore_n186;
   wire FE_PHN3336_U_afifo_U_acore_n208;
   wire FE_PHN3335_U_afifo_U_acore_n178;
   wire FE_PHN3334_U_dfifo_U_dcore_n188;
   wire FE_PHN3333_U_afifo_U_acore_n176;
   wire FE_PHN3332_U_dfifo_U_dcore_n197;
   wire FE_PHN3331_U_afifo_U_acore_n204;
   wire FE_PHN3330_U_dfifo_U_dcore_n179;
   wire FE_PHN3329_U_dfifo_U_dcore_n191;
   wire FE_PHN3323_U_afifo_U_acore_n95;
   wire FE_PHN3310_U_afifo_U_acore_n97;
   wire FE_PHN3308_U_afifo_U_acore_U_sub_fifo_n273;
   wire FE_PHN3307_U_afifo_U_acore_U_sub_fifo_n202;
   wire FE_PHN3306_U_afifo_U_acore_U_sub_fifo_n176;
   wire FE_PHN3304_U_afifo_U_acore_U_sub_fifo_n277;
   wire FE_PHN3303_U_afifo_U_acore_U_sub_fifo_n203;
   wire FE_PHN3302_U_afifo_U_acore_U_sub_fifo_n206;
   wire FE_PHN3301_U_afifo_U_acore_U_sub_fifo_n201;
   wire FE_PHN3300_U_afifo_U_acore_U_sub_fifo_n200;
   wire FE_PHN3296_U_afifo_U_acore_U_sub_fifo_n198;
   wire FE_PHN3295_U_dfifo_U_dcore_U_sub_fifo_n450;
   wire FE_PHN3294_U_afifo_U_acore_U_sub_fifo_n249;
   wire FE_PHN3285_U_afifo_U_acore_U_sub_fifo_n269;
   wire FE_PHN3284_U_dfifo_n3;
   wire FE_PHN3281_U_rbuf_n82;
   wire FE_PHN3280_U_rbuf_n84;
   wire FE_PHN3279_U_rbuf_n85;
   wire FE_PHN3272_U_rbuf_n71;
   wire FE_PHN3271_U_ctl_n141;
   wire FE_PHN3270_U_ctl_n123;
   wire FE_PHN3269_U_ctl_n139;
   wire FE_PHN3267_U_afifo_U_acore_n142;
   wire FE_PHN3266_U_dfifo_U_dcore_n167;
   wire FE_PHN3265_U_afifo_U_acore_n144;
   wire FE_PHN3264_U_afifo_U_acore_n138;
   wire FE_PHN3263_U_afifo_U_acore_n162;
   wire FE_PHN3262_U_afifo_U_acore_n160;
   wire FE_PHN3261_U_afifo_U_acore_n33;
   wire FE_PHN3257_U_afifo_U_acore_n104;
   wire FE_PHN3254_U_afifo_U_acore_n121;
   wire FE_PHN3253_U_afifo_U_acore_n115;
   wire FE_PHN3251_U_afifo_U_acore_n147;
   wire FE_PHN3248_U_afifo_U_acore_n94;
   wire FE_PHN3246_U_dfifo_U_dcore_f_buf_data_0_;
   wire FE_PHN3243_U_afifo_U_acore_n199;
   wire FE_PHN3236_U_dfifo_U_dcore_n157;
   wire FE_PHN3226_U_dfifo_U_dcore_n155;
   wire FE_PHN3225_U_afifo_m_data_in_14_;
   wire FE_PHN3219_U_dfifo_U_dcore_n145;
   wire FE_PHN3218_U_dfifo_U_dcore_U_sub_fifo_n452;
   wire FE_PHN3214_U_dfifo_U_dcore_n148;
   wire FE_PHN3213_U_afifo_m_data_in_12_;
   wire FE_PHN3210_U_afifo_m_data_in_4_;
   wire FE_PHN3207_U_ctl_n117;
   wire FE_PHN3203_U_ctl_n120;
   wire FE_PHN3184_U_afifo_U_acore_U_sub_fifo_n287;
   wire FE_PHN3181_U_afifo_U_acore_U_sub_fifo_n322;
   wire FE_PHN3180_U_afifo_U_acore_n133;
   wire FE_PHN3179_U_afifo_U_acore_U_sub_fifo_n305;
   wire FE_PHN3178_U_afifo_U_acore_U_sub_fifo_n292;
   wire FE_PHN3177_U_afifo_U_acore_U_sub_fifo_n310;
   wire FE_PHN3176_U_afifo_U_acore_U_sub_fifo_n316;
   wire FE_PHN3175_U_afifo_U_acore_U_sub_fifo_n297;
   wire FE_PHN3174_U_afifo_U_acore_U_sub_fifo_n294;
   wire FE_PHN3173_U_afifo_U_acore_U_sub_fifo_n278;
   wire FE_PHN3172_U_afifo_U_acore_U_sub_fifo_n274;
   wire FE_PHN3171_U_afifo_U_acore_U_sub_fifo_n308;
   wire FE_PHN3163_U_afifo_U_acore_U_sub_fifo_n296;
   wire FE_PHN3161_U_afifo_U_acore_U_sub_fifo_n295;
   wire FE_PHN3159_U_afifo_U_acore_U_sub_fifo_n280;
   wire FE_PHN3158_U_afifo_U_acore_U_sub_fifo_n318;
   wire FE_PHN3157_U_afifo_U_acore_U_sub_fifo_n307;
   wire FE_PHN3155_U_ctl_n133;
   wire FE_PHN3154_U_ctl_n134;
   wire FE_PHN3152_U_ctl_n118;
   wire FE_PHN3151_U_ctl_n130;
   wire FE_PHN3150_U_ctl_n137;
   wire FE_PHN3149_U_ctl_n140;
   wire FE_PHN3148_U_ctl_n129;
   wire FE_PHN3147_U_ctl_n131;
   wire FE_PHN3146_U_ctl_n128;
   wire FE_PHN3145_U_ctl_n125;
   wire FE_PHN3144_U_ctl_n106;
   wire FE_PHN3141_U_ctl_n421;
   wire FE_PHN3132_U_dfifo_U_dcore_n139;
   wire FE_PHN3131_U_dfifo_U_dcore_n141;
   wire FE_PHN3130_U_dfifo_U_dcore_n137;
   wire FE_PHN3129_U_dfifo_U_dcore_n138;
   wire FE_PHN3128_U_dfifo_U_dcore_n135;
   wire FE_PHN3125_U_dfifo_U_dcore_n203;
   wire FE_PHN3124_U_dfifo_U_dcore_f_buf_data_6_;
   wire FE_PHN3122_U_dfifo_U_dcore_f_buf_data_19_;
   wire FE_PHN3121_U_dfifo_U_dcore_f_buf_data_7_;
   wire FE_PHN3120_U_dfifo_U_dcore_f_buf_data_3_;
   wire FE_PHN3118_U_dfifo_U_dcore_f_buf_data_15_;
   wire FE_PHN3117_U_dfifo_U_dcore_f_buf_data_17_;
   wire FE_PHN3116_U_dfifo_U_dcore_f_buf_data_22_;
   wire FE_PHN3114_U_dfifo_U_dcore_f_buf_data_9_;
   wire FE_PHN3096_U_ctl_n135;
   wire FE_PHN3095_U_ctl_n119;
   wire FE_PHN3062_U_ctl_n122;
   wire FE_PHN3042_U_ctl_n138;
   wire FE_PHN3040_U_dfifo_U_dcore_f_buf_data_30_;
   wire FE_PHN3039_U_dfifo_U_dcore_f_buf_data_2_;
   wire FE_PHN3038_U_dfifo_U_dcore_f_buf_data_5_;
   wire FE_PHN3037_U_dfifo_U_dcore_f_buf_data_31_;
   wire FE_PHN3036_U_dfifo_U_dcore_f_buf_data_4_;
   wire FE_PHN3035_U_dfifo_U_dcore_f_buf_data_28_;
   wire FE_PHN3032_U_afifo_n_new_req;
   wire FE_PHN3027_U_rbuf_n63;
   wire FE_PHN3026_U_rbuf_n64;
   wire FE_PHN3025_U_rbuf_n83;
   wire FE_PHN3024_U_rbuf_n65;
   wire FE_PHN3023_U_rbuf_n72;
   wire FE_PHN3022_U_rbuf_n59;
   wire FE_PHN3021_U_rbuf_n77;
   wire FE_PHN3020_U_rbuf_n60;
   wire FE_PHN3019_U_rbuf_n80;
   wire FE_PHN3017_U_rbuf_n76;
   wire FE_PHN3016_U_rbuf_n81;
   wire FE_PHN3015_U_rbuf_n74;
   wire FE_PHN3014_U_ctl_n124;
   wire FE_PHN3008_U_rbuf_n56;
   wire FE_PHN3007_U_rbuf_n67;
   wire FE_PHN3006_U_rbuf_n61;
   wire FE_PHN3005_U_rbuf_n70;
   wire FE_PHN3004_U_rbuf_n57;
   wire FE_PHN3003_U_rbuf_n58;
   wire FE_PHN3002_hiu_terminate;
   wire FE_PHN2999_U_rbuf_n73;
   wire FE_PHN2998_U_rbuf_n86;
   wire FE_PHN2997_U_rbuf_n79;
   wire FE_PHN2996_U_rbuf_n75;
   wire FE_PHN2979_U_afifo_U_acore_U_sub_fifo_count_0_;
   wire FE_PHN2963_U_ctl_n132;
   wire FE_PHN2957_U_rbuf_n62;
   wire FE_PHN2949_U_rbuf_n78;
   wire FE_PHN2940_U_rbuf_n55;
   wire FE_PHN2938_U_rbuf_n69;
   wire FE_PHN2937_U_rbuf_n66;
   wire FE_PHN2934_U_rbuf_n68;
   wire FE_PHN2933_U_ctl_n127;
   wire FE_PHN2930_U_rbuf_n89;
   wire FE_PHN2924_m_rb_overflow;
   wire FE_PHN2923_U_ctl_n212;
   wire FE_PHN2917_hsel_reg;
   wire FE_PHN2914_U_ctl_n382;
   wire FE_PHN2913_U_ctl_n422;
   wire FE_PHN2908_m_af_push1_n;
   wire FE_PHN2904_U_ctl_f_burst_done;
   wire FE_PHN2704_U_afifo_n20;
   wire FE_PHN2677_U_afifo_n19;
   wire FE_PHN2656_U_afifo_n18;
   wire FE_PHN2638_U_afifo_n159;
   wire FE_PHN2575_U_afifo_n166;
   wire FE_PHN2567_U_afifo_n165;
   wire FE_PHN2565_U_afifo_n191;
   wire FE_PHN2558_U_afifo_n160;
   wire FE_PHN2434_U_afifo_n158;
   wire FE_PHN2433_U_afifo_n164;
   wire FE_PHN2421_U_dfifo_U_dcore_U_sub_fifo_n448;
   wire FE_PHN2375_U_dfifo_U_dcore_U_sub_fifo_n272;
   wire FE_PHN2374_U_dfifo_U_dcore_U_sub_fifo_n271;
   wire FE_PHN2372_U_dfifo_U_dcore_U_sub_fifo_n303;
   wire FE_PHN2371_U_dfifo_U_dcore_U_sub_fifo_n306;
   wire FE_PHN2370_U_dfifo_U_dcore_U_sub_fifo_n294;
   wire FE_PHN2369_U_dfifo_U_dcore_U_sub_fifo_n260;
   wire FE_PHN2368_U_dfifo_U_dcore_U_sub_fifo_n295;
   wire FE_PHN2367_U_dfifo_U_dcore_U_sub_fifo_n309;
   wire FE_PHN2366_U_dfifo_U_dcore_U_sub_fifo_n278;
   wire FE_PHN2365_U_dfifo_U_dcore_U_sub_fifo_n305;
   wire FE_PHN2363_U_dfifo_U_dcore_U_sub_fifo_n275;
   wire FE_PHN2362_U_afifo_U_acore_U_sub_fifo_n248;
   wire FE_PHN2361_U_dfifo_U_dcore_U_sub_fifo_n269;
   wire FE_PHN2360_U_dfifo_U_dcore_U_sub_fifo_n270;
   wire FE_PHN2359_U_afifo_U_acore_U_sub_fifo_n197;
   wire FE_PHN2358_U_dfifo_U_dcore_U_sub_fifo_n283;
   wire FE_PHN2357_U_dfifo_U_dcore_U_sub_fifo_n268;
   wire FE_PHN2356_U_dfifo_U_dcore_U_sub_fifo_n307;
   wire FE_PHN2354_U_dfifo_U_dcore_U_sub_fifo_n292;
   wire FE_PHN2353_U_dfifo_U_dcore_U_sub_fifo_n257;
   wire FE_PHN2352_U_dfifo_U_dcore_U_sub_fifo_n253;
   wire FE_PHN2351_U_afifo_U_acore_U_sub_fifo_n208;
   wire FE_PHN2350_U_dfifo_U_dcore_U_sub_fifo_n279;
   wire FE_PHN2349_U_dfifo_U_dcore_U_sub_fifo_n265;
   wire FE_PHN2345_U_dfifo_U_dcore_U_sub_fifo_n290;
   wire FE_PHN2344_U_dfifo_U_dcore_U_sub_fifo_n258;
   wire FE_PHN2343_U_afifo_U_acore_U_sub_fifo_n205;
   wire FE_PHN2342_U_dfifo_U_dcore_U_sub_fifo_n255;
   wire FE_PHN2341_U_dfifo_U_dcore_U_sub_fifo_n254;
   wire FE_PHN2340_U_dfifo_U_dcore_U_sub_fifo_n274;
   wire FE_PHN2339_U_dfifo_U_dcore_U_sub_fifo_n267;
   wire FE_PHN2338_U_dfifo_U_dcore_U_sub_fifo_n277;
   wire FE_PHN2337_U_dfifo_U_dcore_U_sub_fifo_n286;
   wire FE_PHN2336_U_dfifo_U_dcore_U_sub_fifo_n276;
   wire FE_PHN2335_U_dfifo_U_dcore_U_sub_fifo_n262;
   wire FE_PHN2334_U_dfifo_U_dcore_U_sub_fifo_n246;
   wire FE_PHN2332_U_dfifo_U_dcore_U_sub_fifo_n249;
   wire FE_PHN2331_U_dfifo_U_dcore_U_sub_fifo_n248;
   wire FE_PHN2329_U_dfifo_U_dcore_U_sub_fifo_n282;
   wire FE_PHN2328_U_afifo_U_acore_U_sub_fifo_n301;
   wire FE_PHN2327_U_dfifo_U_dcore_U_sub_fifo_n299;
   wire FE_PHN2326_U_dfifo_U_dcore_U_sub_fifo_n256;
   wire FE_PHN2325_U_dfifo_U_dcore_U_sub_fifo_n263;
   wire FE_PHN2324_U_afifo_U_acore_U_sub_fifo_n265;
   wire FE_PHN2323_U_dfifo_U_dcore_U_sub_fifo_n250;
   wire FE_PHN2322_U_dfifo_U_dcore_U_sub_fifo_n302;
   wire FE_PHN2321_U_afifo_U_acore_U_sub_fifo_n257;
   wire FE_PHN2320_U_dfifo_U_dcore_U_sub_fifo_n243;
   wire FE_PHN2319_U_dfifo_U_dcore_U_sub_fifo_n261;
   wire FE_PHN2318_U_dfifo_U_dcore_U_sub_fifo_n259;
   wire FE_PHN2317_U_dfifo_U_dcore_U_sub_fifo_n284;
   wire FE_PHN2316_U_afifo_U_acore_U_sub_fifo_n302;
   wire FE_PHN2315_U_afifo_U_acore_U_sub_fifo_n279;
   wire FE_PHN2314_U_dfifo_U_dcore_U_sub_fifo_n289;
   wire FE_PHN2313_U_dfifo_U_dcore_U_sub_fifo_n287;
   wire FE_PHN2312_U_afifo_U_acore_U_sub_fifo_n306;
   wire FE_PHN2311_U_dfifo_U_dcore_U_sub_fifo_n298;
   wire FE_PHN2310_U_dfifo_U_dcore_U_sub_fifo_n266;
   wire FE_PHN2309_U_dfifo_U_dcore_U_sub_fifo_n245;
   wire FE_PHN2308_U_afifo_U_acore_U_sub_fifo_n259;
   wire FE_PHN2307_U_dfifo_U_dcore_U_sub_fifo_n310;
   wire FE_PHN2306_U_dfifo_U_dcore_U_sub_fifo_n300;
   wire FE_PHN2305_U_dfifo_U_dcore_U_sub_fifo_n244;
   wire FE_PHN2304_U_dfifo_U_dcore_U_sub_fifo_n273;
   wire FE_PHN2303_U_dfifo_U_dcore_U_sub_fifo_n301;
   wire FE_PHN2301_U_dfifo_U_dcore_U_sub_fifo_n296;
   wire FE_PHN2299_U_dfifo_U_dcore_U_sub_fifo_n304;
   wire FE_PHN2298_U_dfifo_U_dcore_U_sub_fifo_n293;
   wire FE_PHN2297_U_dfifo_U_dcore_U_sub_fifo_n308;
   wire FE_PHN2296_U_dfifo_U_dcore_U_sub_fifo_n247;
   wire FE_PHN2295_U_afifo_U_acore_U_sub_fifo_n173;
   wire FE_PHN2293_U_dfifo_U_dcore_U_sub_fifo_n252;
   wire FE_PHN2292_U_afifo_U_acore_U_sub_fifo_n180;
   wire FE_PHN2291_U_dfifo_U_dcore_U_sub_fifo_n280;
   wire FE_PHN2290_U_afifo_U_acore_U_sub_fifo_n210;
   wire FE_PHN2289_U_dfifo_U_dcore_U_sub_fifo_n288;
   wire FE_PHN2288_U_dfifo_U_dcore_U_sub_fifo_n251;
   wire FE_PHN2287_U_afifo_U_acore_U_sub_fifo_n194;
   wire FE_PHN2285_U_dfifo_U_dcore_U_sub_fifo_n281;
   wire FE_PHN2284_U_dfifo_U_dcore_U_sub_fifo_n291;
   wire FE_PHN2283_U_dfifo_U_dcore_U_sub_fifo_n297;
   wire FE_PHN2282_U_afifo_U_acore_U_sub_fifo_n224;
   wire FE_PHN2281_U_afifo_U_acore_U_sub_fifo_n213;
   wire FE_PHN2280_U_dfifo_U_dcore_U_sub_fifo_n285;
   wire FE_PHN2279_U_afifo_U_acore_U_sub_fifo_n211;
   wire FE_PHN2278_U_afifo_U_acore_U_sub_fifo_n177;
   wire FE_PHN2277_U_afifo_U_acore_U_sub_fifo_n226;
   wire FE_PHN2276_U_afifo_U_acore_U_sub_fifo_n253;
   wire FE_PHN2275_U_afifo_U_acore_U_sub_fifo_n200;
   wire FE_PHN2274_U_afifo_U_acore_U_sub_fifo_n243;
   wire FE_PHN2273_U_afifo_U_acore_U_sub_fifo_n245;
   wire FE_PHN2272_U_afifo_U_acore_U_sub_fifo_n215;
   wire FE_PHN2271_U_afifo_U_acore_U_sub_fifo_n300;
   wire FE_PHN2269_U_afifo_U_acore_U_sub_fifo_n252;
   wire FE_PHN2268_U_afifo_U_acore_U_sub_fifo_n256;
   wire FE_PHN2267_U_afifo_U_acore_U_sub_fifo_n249;
   wire FE_PHN2266_U_afifo_U_acore_U_sub_fifo_n203;
   wire FE_PHN2265_U_afifo_U_acore_U_sub_fifo_n319;
   wire FE_PHN2264_U_afifo_U_acore_U_sub_fifo_n179;
   wire FE_PHN2263_U_afifo_U_acore_U_sub_fifo_n191;
   wire FE_PHN2262_U_afifo_U_acore_U_sub_fifo_n183;
   wire FE_PHN2261_U_afifo_U_acore_U_sub_fifo_n283;
   wire FE_PHN2260_U_afifo_U_acore_U_sub_fifo_n227;
   wire FE_PHN2259_U_afifo_U_acore_U_sub_fifo_n289;
   wire FE_PHN2258_U_afifo_U_acore_U_sub_fifo_n198;
   wire FE_PHN2257_U_afifo_U_acore_U_sub_fifo_n284;
   wire FE_PHN2256_U_afifo_U_acore_U_sub_fifo_n237;
   wire FE_PHN2255_U_afifo_U_acore_U_sub_fifo_n228;
   wire FE_PHN2253_U_afifo_U_acore_U_sub_fifo_n186;
   wire FE_PHN2252_U_afifo_U_acore_U_sub_fifo_n246;
   wire FE_PHN2251_U_afifo_U_acore_U_sub_fifo_n199;
   wire FE_PHN2250_U_afifo_U_acore_U_sub_fifo_n234;
   wire FE_PHN2249_U_afifo_U_acore_U_sub_fifo_n258;
   wire FE_PHN2248_U_afifo_U_acore_U_sub_fifo_n189;
   wire FE_PHN2247_U_afifo_U_acore_U_sub_fifo_n204;
   wire FE_PHN2246_U_afifo_U_acore_U_sub_fifo_n254;
   wire FE_PHN2244_U_afifo_U_acore_U_sub_fifo_n276;
   wire FE_PHN2243_U_afifo_U_acore_U_sub_fifo_n241;
   wire FE_PHN2242_U_afifo_U_acore_U_sub_fifo_n185;
   wire FE_PHN2239_U_afifo_U_acore_U_sub_fifo_n235;
   wire FE_PHN2238_U_afifo_U_acore_U_sub_fifo_n286;
   wire FE_PHN2237_U_afifo_U_acore_U_sub_fifo_n231;
   wire FE_PHN2236_U_afifo_U_acore_U_sub_fifo_n192;
   wire FE_PHN2235_U_dfifo_U_dcore_U_sub_fifo_n396;
   wire FE_PHN2234_U_afifo_U_acore_U_sub_fifo_n181;
   wire FE_PHN2231_U_afifo_U_acore_U_sub_fifo_n182;
   wire FE_PHN2230_U_afifo_U_acore_U_sub_fifo_n232;
   wire FE_PHN2229_U_dfifo_U_dcore_U_sub_fifo_n374;
   wire FE_PHN2228_U_afifo_U_acore_U_sub_fifo_n290;
   wire FE_PHN2227_U_afifo_U_acore_U_sub_fifo_n190;
   wire FE_PHN2226_U_afifo_U_acore_U_sub_fifo_n288;
   wire FE_PHN2222_U_dfifo_U_dcore_U_sub_fifo_n376;
   wire FE_PHN2221_U_dfifo_U_dcore_U_sub_fifo_n350;
   wire FE_PHN2220_U_dfifo_U_dcore_U_sub_fifo_n430;
   wire FE_PHN2218_U_dfifo_U_dcore_U_sub_fifo_n422;
   wire FE_PHN2217_U_dfifo_U_dcore_U_sub_fifo_n381;
   wire FE_PHN2216_U_dfifo_U_dcore_U_sub_fifo_n337;
   wire FE_PHN2214_U_dfifo_U_dcore_U_sub_fifo_n388;
   wire FE_PHN2213_U_dfifo_U_dcore_U_sub_fifo_n427;
   wire FE_PHN2211_U_dfifo_U_dcore_U_sub_fifo_n386;
   wire FE_PHN2209_U_dfifo_U_dcore_U_sub_fifo_n368;
   wire FE_PHN2208_U_dfifo_U_dcore_U_sub_fifo_n445;
   wire FE_PHN2207_U_dfifo_U_dcore_U_sub_fifo_n387;
   wire FE_PHN2206_U_dfifo_U_dcore_U_sub_fifo_n432;
   wire FE_PHN2205_U_dfifo_U_dcore_U_sub_fifo_n314;
   wire FE_PHN2204_U_dfifo_U_dcore_U_sub_fifo_n394;
   wire FE_PHN2203_U_dfifo_U_dcore_U_sub_fifo_n435;
   wire FE_PHN2202_U_dfifo_U_dcore_U_sub_fifo_n373;
   wire FE_PHN2201_U_dfifo_U_dcore_U_sub_fifo_n434;
   wire FE_PHN2199_U_dfifo_U_dcore_U_sub_fifo_n423;
   wire FE_PHN2198_U_dfifo_U_dcore_U_sub_fifo_n433;
   wire FE_PHN2197_U_dfifo_U_dcore_U_sub_fifo_n426;
   wire FE_PHN2195_U_dfifo_U_dcore_U_sub_fifo_n428;
   wire FE_PHN2194_U_dfifo_U_dcore_U_sub_fifo_n437;
   wire FE_PHN2193_U_dfifo_U_dcore_U_sub_fifo_n421;
   wire FE_PHN2192_U_dfifo_U_dcore_U_sub_fifo_n384;
   wire FE_PHN2191_U_dfifo_U_dcore_U_sub_fifo_n436;
   wire FE_PHN2190_U_dfifo_U_dcore_U_sub_fifo_n379;
   wire FE_PHN2188_U_dfifo_U_dcore_U_sub_fifo_n385;
   wire FE_PHN2186_U_dfifo_U_dcore_U_sub_fifo_n431;
   wire FE_PHN2185_U_dfifo_U_dcore_U_sub_fifo_n380;
   wire FE_PHN2184_U_dfifo_U_dcore_U_sub_fifo_n366;
   wire FE_PHN2183_U_dfifo_U_dcore_U_sub_fifo_n429;
   wire FE_PHN2182_U_dfifo_U_dcore_U_sub_fifo_n365;
   wire FE_PHN2178_U_dfifo_U_dcore_U_sub_fifo_n382;
   wire FE_PHN2177_U_dfifo_U_dcore_U_sub_fifo_n424;
   wire FE_PHN2176_U_dfifo_U_dcore_U_sub_fifo_n389;
   wire FE_PHN2175_U_dfifo_U_dcore_U_sub_fifo_n317;
   wire FE_PHN2174_U_dfifo_U_dcore_U_sub_fifo_n390;
   wire FE_PHN2173_U_dfifo_U_dcore_U_sub_fifo_n391;
   wire FE_PHN2172_U_dfifo_U_dcore_U_sub_fifo_n425;
   wire FE_PHN2171_U_dfifo_U_dcore_U_sub_fifo_n419;
   wire FE_PHN2170_U_dfifo_U_dcore_U_sub_fifo_n383;
   wire FE_PHN2169_U_dfifo_U_dcore_U_sub_fifo_n392;
   wire FE_PHN2168_U_dfifo_U_dcore_U_sub_fifo_n393;
   wire FE_PHN2167_U_dfifo_U_dcore_U_sub_fifo_n321;
   wire FE_PHN2165_U_dfifo_U_dcore_U_sub_fifo_n413;
   wire FE_PHN2162_U_dfifo_U_dcore_U_sub_fifo_n395;
   wire FE_PHN2161_U_afifo_f_data2_7_;
   wire FE_PHN2160_U_dfifo_U_dcore_U_sub_fifo_n313;
   wire FE_PHN2159_U_dfifo_U_dcore_U_sub_fifo_n363;
   wire FE_PHN2158_U_dfifo_U_dcore_U_sub_fifo_n401;
   wire FE_PHN2155_U_dfifo_U_dcore_U_sub_fifo_n420;
   wire FE_PHN2153_U_dfifo_U_dcore_U_sub_fifo_n416;
   wire FE_PHN2152_U_dfifo_U_dcore_U_sub_fifo_n333;
   wire FE_PHN2151_U_dfifo_U_dcore_U_sub_fifo_n361;
   wire FE_PHN2147_U_dfifo_U_dcore_U_sub_fifo_n443;
   wire FE_PHN2144_U_dfifo_U_dcore_U_sub_fifo_n326;
   wire FE_PHN2142_U_dfifo_U_dcore_U_sub_fifo_n315;
   wire FE_PHN2139_U_dfifo_U_dcore_U_sub_fifo_n405;
   wire FE_PHN2138_U_dfifo_U_dcore_U_sub_fifo_n403;
   wire FE_PHN2137_U_dfifo_U_dcore_U_sub_fifo_n322;
   wire FE_PHN2136_U_dfifo_U_dcore_U_sub_fifo_n411;
   wire FE_PHN2135_U_dfifo_U_dcore_U_sub_fifo_n402;
   wire FE_PHN2134_U_dfifo_U_dcore_U_sub_fifo_n325;
   wire FE_PHN2133_U_afifo_n3;
   wire FE_PHN2132_U_dfifo_U_dcore_U_sub_fifo_n400;
   wire FE_PHN2131_U_dfifo_U_dcore_U_sub_fifo_n328;
   wire FE_PHN2130_U_dfifo_U_dcore_U_sub_fifo_n438;
   wire FE_PHN2129_U_dfifo_U_dcore_U_sub_fifo_n342;
   wire FE_PHN2128_U_dfifo_U_dcore_U_sub_fifo_n320;
   wire FE_PHN2127_U_dfifo_U_dcore_U_sub_fifo_n414;
   wire FE_PHN2126_U_dfifo_U_dcore_U_sub_fifo_n319;
   wire FE_PHN2124_U_dfifo_U_dcore_U_sub_fifo_n312;
   wire FE_PHN2123_U_dfifo_U_dcore_U_sub_fifo_n323;
   wire FE_PHN2122_U_dfifo_U_dcore_U_sub_fifo_n406;
   wire FE_PHN2121_U_dfifo_U_dcore_U_sub_fifo_n412;
   wire FE_PHN2119_U_dfifo_U_dcore_U_sub_fifo_n444;
   wire FE_PHN2118_U_dfifo_U_dcore_U_sub_fifo_n441;
   wire FE_PHN2117_U_dfifo_U_dcore_U_sub_fifo_n409;
   wire FE_PHN2116_U_dfifo_U_dcore_U_sub_fifo_n408;
   wire FE_PHN2115_U_dfifo_U_dcore_U_sub_fifo_n369;
   wire FE_PHN2113_U_dfifo_U_dcore_U_sub_fifo_n311;
   wire FE_PHN2112_U_dfifo_U_dcore_U_sub_fifo_n404;
   wire FE_PHN2111_U_dfifo_U_dcore_U_sub_fifo_n439;
   wire FE_PHN2110_U_dfifo_U_dcore_U_sub_fifo_n372;
   wire FE_PHN2108_U_dfifo_U_dcore_U_sub_fifo_n316;
   wire FE_PHN2026_U_afifo_U_acore_U_sub_fifo_n298;
   wire FE_PHN2024_U_afifo_U_acore_U_sub_fifo_n223;
   wire FE_PHN2023_U_dfifo_U_dcore_U_sub_fifo_n264;
   wire FE_PHN2022_U_afifo_U_acore_U_sub_fifo_n275;
   wire FE_PHN2021_U_afifo_U_acore_U_sub_fifo_n250;
   wire FE_PHN2020_U_afifo_U_acore_U_sub_fifo_n218;
   wire FE_PHN2019_U_afifo_U_acore_U_sub_fifo_n176;
   wire FE_PHN2018_U_afifo_U_acore_U_sub_fifo_n196;
   wire FE_PHN2017_U_afifo_U_acore_U_sub_fifo_n175;
   wire FE_PHN2016_U_afifo_U_acore_U_sub_fifo_n311;
   wire FE_PHN2015_U_afifo_U_acore_U_sub_fifo_n174;
   wire FE_PHN2014_U_afifo_U_acore_U_sub_fifo_n309;
   wire FE_PHN2013_U_afifo_U_acore_U_sub_fifo_n230;
   wire FE_PHN2012_U_afifo_U_acore_U_sub_fifo_n207;
   wire FE_PHN2011_U_afifo_U_acore_U_sub_fifo_n261;
   wire FE_PHN2010_U_afifo_U_acore_U_sub_fifo_n247;
   wire FE_PHN2009_U_afifo_U_acore_U_sub_fifo_n193;
   wire FE_PHN2008_U_afifo_U_acore_U_sub_fifo_n178;
   wire FE_PHN2007_U_afifo_U_acore_U_sub_fifo_n202;
   wire FE_PHN2006_U_afifo_U_acore_U_sub_fifo_n201;
   wire FE_PHN2005_U_afifo_U_acore_U_sub_fifo_n244;
   wire FE_PHN2004_U_dfifo_U_dcore_U_sub_fifo_n378;
   wire FE_PHN2003_U_afifo_U_acore_U_sub_fifo_n293;
   wire FE_PHN2002_U_afifo_U_acore_U_sub_fifo_n313;
   wire FE_PHN2001_U_afifo_U_acore_U_sub_fifo_n195;
   wire FE_PHN2000_U_afifo_U_acore_U_sub_fifo_n263;
   wire FE_PHN1999_U_afifo_U_acore_U_sub_fifo_n229;
   wire FE_PHN1998_U_afifo_U_acore_U_sub_fifo_n299;
   wire FE_PHN1997_U_dfifo_U_dcore_U_sub_fifo_n375;
   wire FE_PHN1996_U_afifo_U_acore_U_sub_fifo_n217;
   wire FE_PHN1995_U_afifo_U_acore_U_sub_fifo_n251;
   wire FE_PHN1994_U_afifo_U_acore_U_sub_fifo_n206;
   wire FE_PHN1993_U_afifo_U_acore_U_sub_fifo_n225;
   wire FE_PHN1992_U_afifo_U_acore_U_sub_fifo_n303;
   wire FE_PHN1991_U_afifo_U_acore_U_sub_fifo_n260;
   wire FE_PHN1990_U_dfifo_U_dcore_U_sub_fifo_n377;
   wire FE_PHN1989_U_afifo_U_acore_U_sub_fifo_n233;
   wire FE_PHN1988_U_afifo_U_acore_U_sub_fifo_n187;
   wire FE_PHN1987_U_afifo_U_acore_U_sub_fifo_n184;
   wire FE_PHN1986_U_afifo_U_acore_U_sub_fifo_n255;
   wire FE_PHN1985_U_afifo_U_acore_U_sub_fifo_n285;
   wire FE_PHN1984_U_afifo_U_acore_U_sub_fifo_n291;
   wire FE_PHN1982_U_afifo_U_acore_U_sub_fifo_n242;
   wire FE_PHN1981_U_afifo_U_acore_U_sub_fifo_n281;
   wire FE_PHN1980_U_afifo_U_acore_U_sub_fifo_n236;
   wire FE_PHN1979_U_afifo_U_acore_U_sub_fifo_n239;
   wire FE_PHN1977_U_afifo_U_acore_U_sub_fifo_n304;
   wire FE_PHN1976_U_afifo_U_acore_U_sub_fifo_n240;
   wire FE_PHN1975_U_afifo_U_acore_U_sub_fifo_n188;
   wire FE_PHN1974_U_afifo_U_acore_U_sub_fifo_n220;
   wire FE_PHN1973_U_afifo_U_acore_U_sub_fifo_n238;
   wire FE_PHN1972_U_afifo_U_acore_U_sub_fifo_n320;
   wire FE_PHN1971_U_afifo_U_acore_U_sub_fifo_n282;
   wire FE_PHN1969_U_dfifo_U_dcore_U_sub_fifo_n349;
   wire FE_PHN1968_U_dfifo_U_dcore_U_sub_fifo_n364;
   wire FE_PHN1966_U_afifo_U_acore_U_sub_fifo_n267;
   wire FE_PHN1965_U_dfifo_U_dcore_U_sub_fifo_n352;
   wire FE_PHN1964_U_dfifo_U_dcore_U_sub_fifo_n330;
   wire FE_PHN1963_U_dfifo_U_dcore_U_sub_fifo_n360;
   wire FE_PHN1962_U_afifo_U_acore_U_sub_fifo_n272;
   wire FE_PHN1961_U_dfifo_U_dcore_U_sub_fifo_n346;
   wire FE_PHN1960_U_dfifo_U_dcore_U_sub_fifo_n351;
   wire FE_PHN1959_U_afifo_U_acore_U_sub_fifo_n266;
   wire FE_PHN1958_U_dfifo_U_dcore_U_sub_fifo_n367;
   wire FE_PHN1957_U_dfifo_U_dcore_U_sub_fifo_n347;
   wire FE_PHN1956_U_dfifo_U_dcore_U_sub_fifo_n407;
   wire FE_PHN1955_U_dfifo_U_dcore_U_sub_fifo_n358;
   wire FE_PHN1954_U_dfifo_U_dcore_U_sub_fifo_n398;
   wire FE_PHN1953_U_dfifo_U_dcore_U_sub_fifo_n415;
   wire FE_PHN1952_U_dfifo_U_dcore_U_sub_fifo_n348;
   wire FE_PHN1951_U_dfifo_U_dcore_U_sub_fifo_n318;
   wire FE_PHN1950_U_afifo_U_acore_U_sub_fifo_n269;
   wire FE_PHN1949_U_dfifo_U_dcore_U_sub_fifo_n345;
   wire FE_PHN1948_U_afifo_U_acore_U_sub_fifo_n270;
   wire FE_PHN1947_U_dfifo_U_dcore_U_sub_fifo_n397;
   wire FE_PHN1946_U_dfifo_U_dcore_U_sub_fifo_n362;
   wire FE_PHN1945_U_dfifo_U_dcore_U_sub_fifo_n355;
   wire FE_PHN1944_U_dfifo_U_dcore_U_sub_fifo_n399;
   wire FE_PHN1943_U_dfifo_U_dcore_U_sub_fifo_n357;
   wire FE_PHN1942_U_dfifo_U_dcore_U_sub_fifo_n371;
   wire FE_PHN1941_U_dfifo_U_dcore_U_sub_fifo_n353;
   wire FE_PHN1940_U_dfifo_U_dcore_U_sub_fifo_n341;
   wire FE_PHN1939_U_dfifo_U_dcore_U_sub_fifo_n327;
   wire FE_PHN1938_U_dfifo_U_dcore_U_sub_fifo_n417;
   wire FE_PHN1937_U_dfifo_U_dcore_U_sub_fifo_n340;
   wire FE_PHN1936_U_dfifo_U_dcore_U_sub_fifo_n324;
   wire FE_PHN1935_U_dfifo_U_dcore_U_sub_fifo_n440;
   wire FE_PHN1933_U_dfifo_U_dcore_U_sub_fifo_n343;
   wire FE_PHN1932_U_dfifo_U_dcore_U_sub_fifo_n334;
   wire FE_PHN1931_U_dfifo_U_dcore_U_sub_fifo_n442;
   wire FE_PHN1930_U_dfifo_U_dcore_U_sub_fifo_n418;
   wire FE_PHN1929_U_dfifo_U_dcore_U_sub_fifo_n446;
   wire FE_PHN1928_U_dfifo_U_dcore_U_sub_fifo_n359;
   wire FE_PHN1927_U_dfifo_U_dcore_U_sub_fifo_n356;
   wire FE_PHN1926_U_dfifo_U_dcore_U_sub_fifo_n410;
   wire FE_PHN1925_U_dfifo_U_dcore_U_sub_fifo_n331;
   wire FE_PHN1924_U_dfifo_U_dcore_U_sub_fifo_n370;
   wire FE_PHN1923_U_dfifo_U_dcore_U_sub_fifo_n335;
   wire FE_PHN1922_U_dfifo_U_dcore_U_sub_fifo_n354;
   wire FE_PHN1907_U_afifo_m_data_in_7_;
   wire FE_PHN1904_U_ctl_n141;
   wire FE_PHN1886_U_afifo_f_data2_38_;
   wire FE_PHN1885_U_afifo_f_data2_44_;
   wire FE_PHN1884_U_afifo_f_data2_42_;
   wire FE_PHN1883_U_afifo_f_data2_31_;
   wire FE_PHN1882_U_afifo_f_data2_18_;
   wire FE_PHN1881_U_afifo_f_data2_5_;
   wire FE_PHN1880_U_afifo_f_data2_20_;
   wire FE_PHN1879_U_afifo_f_data2_0_;
   wire FE_PHN1878_U_afifo_f_data2_37_;
   wire FE_PHN1877_U_afifo_f_data2_6_;
   wire FE_PHN1876_U_afifo_f_data2_24_;
   wire FE_PHN1874_U_afifo_f_data2_23_;
   wire FE_PHN1873_U_afifo_f_data2_26_;
   wire FE_PHN1872_U_afifo_f_data2_43_;
   wire FE_PHN1871_U_afifo_f_data2_39_;
   wire FE_PHN1870_U_afifo_f_data2_35_;
   wire FE_PHN1869_U_afifo_f_data2_40_;
   wire FE_PHN1867_U_afifo_f_data2_27_;
   wire FE_PHN1866_U_afifo_f_data2_29_;
   wire FE_PHN1865_U_afifo_f_data2_25_;
   wire FE_PHN1864_U_afifo_f_data2_22_;
   wire FE_PHN1863_U_afifo_f_data2_32_;
   wire FE_PHN1862_U_afifo_f_data2_2_;
   wire FE_PHN1861_U_afifo_f_data2_30_;
   wire FE_PHN1860_U_afifo_f_data2_19_;
   wire FE_PHN1859_U_afifo_f_data2_36_;
   wire FE_PHN1858_U_afifo_f_data2_28_;
   wire FE_PHN1857_U_afifo_f_data2_34_;
   wire FE_PHN1856_U_afifo_f_data2_33_;
   wire FE_PHN1853_U_afifo_f_data2_21_;
   wire FE_PHN1852_U_afifo_U_acore_n100;
   wire FE_PHN1851_U_afifo_U_acore_n96;
   wire FE_PHN1850_U_afifo_U_acore_n98;
   wire FE_PHN1849_U_afifo_U_acore_n207;
   wire FE_PHN1847_U_afifo_U_acore_n181;
   wire FE_PHN1844_U_afifo_U_acore_n201;
   wire FE_PHN1843_U_afifo_U_acore_U_sub_fifo_n126;
   wire FE_PHN1842_U_dfifo_U_dcore_U_sub_fifo_n451;
   wire FE_PHN1841_U_afifo_U_acore_n184;
   wire FE_PHN1840_U_afifo_U_acore_n194;
   wire FE_PHN1839_U_afifo_U_acore_n203;
   wire FE_PHN1838_n37;
   wire FE_PHN1837_U_afifo_U_acore_n102;
   wire FE_PHN1836_U_afifo_U_acore_n210;
   wire FE_PHN1835_U_afifo_U_acore_n197;
   wire FE_PHN1834_U_afifo_U_acore_n177;
   wire FE_PHN1833_U_afifo_U_acore_U_sub_fifo_n133;
   wire FE_PHN1832_U_afifo_U_acore_U_sub_fifo_n129;
   wire FE_PHN1831_U_afifo_U_acore_U_sub_fifo_n115;
   wire FE_PHN1830_U_afifo_U_acore_U_sub_fifo_n148;
   wire FE_PHN1829_U_afifo_U_acore_U_sub_fifo_n273;
   wire FE_PHN1828_U_afifo_U_acore_U_sub_fifo_n130;
   wire FE_PHN1827_U_afifo_U_acore_U_sub_fifo_n125;
   wire FE_PHN1826_U_afifo_U_acore_U_sub_fifo_n134;
   wire FE_PHN1825_U_afifo_U_acore_U_sub_fifo_n106;
   wire FE_PHN1824_U_afifo_U_acore_U_sub_fifo_n314;
   wire FE_PHN1823_U_afifo_U_acore_U_sub_fifo_n264;
   wire FE_PHN1822_U_afifo_U_acore_U_sub_fifo_n122;
   wire FE_PHN1821_U_afifo_U_acore_U_sub_fifo_n136;
   wire FE_PHN1820_U_afifo_U_acore_U_sub_fifo_n139;
   wire FE_PHN1819_U_afifo_U_acore_U_sub_fifo_n219;
   wire FE_PHN1818_U_afifo_m_data_in_27_;
   wire FE_PHN1817_U_afifo_f_data2_41_;
   wire FE_PHN1816_U_afifo_U_acore_U_sub_fifo_n102;
   wire FE_PHN1815_U_afifo_U_acore_U_sub_fifo_n143;
   wire FE_PHN1814_U_afifo_U_acore_U_sub_fifo_n138;
   wire FE_PHN1813_U_afifo_U_acore_U_sub_fifo_n216;
   wire FE_PHN1812_U_afifo_U_acore_U_sub_fifo_n123;
   wire FE_PHN1811_U_afifo_U_acore_U_sub_fifo_n214;
   wire FE_PHN1810_U_afifo_U_acore_U_sub_fifo_n121;
   wire FE_PHN1808_U_afifo_U_acore_U_sub_fifo_n140;
   wire FE_PHN1807_U_afifo_U_acore_U_sub_fifo_n317;
   wire FE_PHN1806_U_afifo_U_acore_U_sub_fifo_n128;
   wire FE_PHN1805_U_afifo_U_acore_U_sub_fifo_n127;
   wire FE_PHN1804_U_afifo_U_acore_U_sub_fifo_n146;
   wire FE_PHN1803_U_afifo_U_acore_U_sub_fifo_n277;
   wire FE_PHN1802_U_dfifo_U_dcore_U_sub_fifo_n80;
   wire FE_PHN1801_U_afifo_U_acore_U_sub_fifo_n108;
   wire FE_PHN1800_U_afifo_U_acore_U_sub_fifo_n145;
   wire FE_PHN1799_U_afifo_U_acore_U_sub_fifo_n135;
   wire FE_PHN1798_n27;
   wire FE_PHN1797_U_afifo_U_acore_U_sub_fifo_n131;
   wire FE_PHN1796_U_afifo_U_acore_U_sub_fifo_n120;
   wire FE_PHN1795_U_dfifo_U_dcore_U_sub_fifo_n82;
   wire FE_PHN1794_U_afifo_U_acore_U_sub_fifo_n222;
   wire FE_PHN1793_U_afifo_U_acore_U_sub_fifo_n104;
   wire FE_PHN1792_U_afifo_U_acore_U_sub_fifo_n124;
   wire FE_PHN1791_U_dfifo_U_dcore_U_sub_fifo_n55;
   wire FE_PHN1790_U_dfifo_U_dcore_U_sub_fifo_n79;
   wire FE_PHN1789_U_afifo_m_data_in_28_;
   wire FE_PHN1788_U_dfifo_U_dcore_U_sub_fifo_n81;
   wire FE_PHN1787_U_dfifo_U_dcore_U_sub_fifo_n63;
   wire FE_PHN1786_U_afifo_m_data_in_19_;
   wire FE_PHN1785_U_dfifo_U_dcore_U_sub_fifo_n62;
   wire FE_PHN1784_U_afifo_U_acore_U_sub_fifo_n268;
   wire FE_PHN1783_U_afifo_m_data_in_33_;
   wire FE_PHN1782_U_dfifo_U_dcore_U_sub_fifo_n73;
   wire FE_PHN1781_U_dfifo_U_dcore_U_sub_fifo_n69;
   wire FE_PHN1780_U_dfifo_U_dcore_U_sub_fifo_n329;
   wire FE_PHN1779_U_dfifo_U_dcore_U_sub_fifo_n78;
   wire FE_PHN1778_U_dfifo_U_dcore_U_sub_fifo_n65;
   wire FE_PHN1777_n25;
   wire FE_PHN1776_U_dfifo_U_dcore_U_sub_fifo_n71;
   wire FE_PHN1775_U_dfifo_U_dcore_U_sub_fifo_n70;
   wire FE_PHN1774_U_dfifo_U_dcore_U_sub_fifo_n59;
   wire FE_PHN1773_U_dfifo_U_dcore_U_sub_fifo_n64;
   wire FE_PHN1772_U_dfifo_U_dcore_U_sub_fifo_n72;
   wire FE_PHN1771_U_dfifo_U_dcore_U_sub_fifo_n60;
   wire FE_PHN1770_U_dfifo_U_dcore_U_sub_fifo_n338;
   wire FE_PHN1769_U_afifo_m_data_in_20_;
   wire FE_PHN1768_U_dfifo_U_dcore_U_sub_fifo_n61;
   wire FE_PHN1767_U_dfifo_U_dcore_U_sub_fifo_n58;
   wire FE_PHN1766_U_dfifo_U_dcore_U_sub_fifo_n68;
   wire FE_PHN1765_U_dfifo_U_dcore_U_sub_fifo_n66;
   wire FE_PHN1764_U_dfifo_U_dcore_U_sub_fifo_n67;
   wire FE_PHN1763_U_afifo_m_data_in_31_;
   wire FE_PHN1762_n39;
   wire FE_PHN1761_U_dfifo_U_dcore_U_sub_fifo_n344;
   wire FE_PHN1760_U_dfifo_U_dcore_U_sub_fifo_n76;
   wire FE_PHN1758_U_dfifo_U_dcore_U_sub_fifo_n332;
   wire FE_PHN1757_U_afifo_f_core_ready;
   wire FE_PHN1756_U_dfifo_U_dcore_U_sub_fifo_n339;
   wire FE_PHN1755_U_dfifo_U_dcore_U_sub_fifo_n74;
   wire FE_PHN1754_U_dfifo_U_dcore_U_sub_fifo_n75;
   wire FE_PHN1753_U_dfifo_U_dcore_U_sub_fifo_n77;
   wire FE_PHN1752_U_dfifo_U_dcore_U_sub_fifo_n336;
   wire FE_PHN1750_U_afifo_m_data_in_30_;
   wire FE_PHN1749_U_afifo_m_data_in_21_;
   wire FE_PHN1691_U_afifo_n10;
   wire FE_PHN1689_n29;
   wire FE_PHN1688_U_afifo_m_data_in_24_;
   wire FE_PHN1687_U_afifo_m_data_in_2_;
   wire FE_PHN1686_U_afifo_m_data_in_43_;
   wire FE_PHN1685_U_afifo_m_data_in_23_;
   wire FE_PHN1684_U_ctl_n120;
   wire FE_PHN1681_U_ctl_n117;
   wire FE_PHN1680_U_afifo_m_data_in_49_;
   wire FE_PHN1679_U_rbuf_n82;
   wire FE_PHN1678_U_rbuf_n84;
   wire FE_PHN1677_U_rbuf_n85;
   wire FE_PHN1676_U_rbuf_n71;
   wire FE_PHN1675_U_ctl_n421;
   wire FE_PHN1660_U_dfifo_U_dcore_n_empty;
   wire FE_PHN1650_U_dfifo_U_dcore_n169;
   wire FE_PHN1635_U_afifo_U_acore_U_sub_fifo_n323;
   wire FE_PHN1630_U_dfifo_U_dcore_n145;
   wire FE_PHN1622_U_afifo_m_data_in_15_;
   wire FE_PHN1621_U_afifo_m_data_in_17_;
   wire FE_PHN1620_U_afifo_m_data_in_16_;
   wire FE_PHN1619_U_afifo_n14;
   wire FE_PHN1618_U_afifo_m_data_in_14_;
   wire FE_PHN1616_U_afifo_m_data_in_48_;
   wire FE_PHN1611_U_ctl_n137;
   wire FE_PHN1609_U_ctl_n140;
   wire FE_PHN1607_U_afifo_n5;
   wire FE_PHN1605_U_ctl_n118;
   wire FE_PHN1604_U_ctl_n106;
   wire FE_PHN1595_U_dfifo_U_dcore_U_sub_fifo_count_0_;
   wire FE_PHN1592_U_afifo_U_acore_U_sub_fifo_out_ptr_0_;
   wire FE_PHN1591_U_dfifo_U_dcore_U_sub_fifo_n242;
   wire FE_PHN1584_U_dfifo_U_dcore_U_sub_fifo_n18;
   wire FE_PHN1579_U_dfifo_U_dcore_n168;
   wire FE_PHN1564_U_afifo_U_acore_n186;
   wire FE_PHN1563_U_afifo_U_acore_n192;
   wire FE_PHN1562_U_dfifo_U_dcore_n186;
   wire FE_PHN1561_U_afifo_U_acore_n205;
   wire FE_PHN1560_U_afifo_U_acore_n175;
   wire FE_PHN1558_U_afifo_U_acore_n190;
   wire FE_PHN1556_U_dfifo_U_dcore_U_sub_fifo_n83;
   wire FE_PHN1554_U_afifo_U_acore_n179;
   wire FE_PHN1553_U_afifo_U_acore_U_sub_fifo_n209;
   wire FE_PHN1552_U_afifo_U_acore_n80;
   wire FE_PHN1550_U_dfifo_U_dcore_n193;
   wire FE_PHN1547_U_dfifo_U_dcore_n194;
   wire FE_PHN1546_U_dfifo_U_dcore_U_sub_fifo_n125;
   wire FE_PHN1545_U_dfifo_U_dcore_U_sub_fifo_n123;
   wire FE_PHN1544_U_dfifo_U_dcore_n201;
   wire FE_PHN1543_U_dfifo_U_dcore_U_sub_fifo_n120;
   wire FE_PHN1542_U_dfifo_U_dcore_U_sub_fifo_n122;
   wire FE_PHN1541_U_dfifo_U_dcore_U_sub_fifo_n118;
   wire FE_PHN1540_U_dfifo_U_dcore_U_sub_fifo_n124;
   wire FE_PHN1539_U_dfifo_U_dcore_U_sub_fifo_n119;
   wire FE_PHN1527_U_afifo_n152;
   wire FE_PHN1525_n17;
   wire FE_PHN1515_U_afifo_m_data_in_29_;
   wire FE_PHN1513_U_afifo_m_data_in_38_;
   wire FE_PHN1511_U_ctl_n130;
   wire FE_PHN1510_U_ctl_n128;
   wire FE_PHN1509_U_ctl_n129;
   wire FE_PHN1507_U_ctl_n131;
   wire FE_PHN1506_U_ctl_n394;
   wire FE_PHN1505_U_ctl_n119;
   wire FE_PHN1498_U_dfifo_U_dcore_n203;
   wire FE_PHN1474_U_afifo_U_acore_U_sub_fifo_n315;
   wire FE_PHN1471_U_afifo_U_acore_U_sub_fifo_n324;
   wire FE_PHN1467_U_dfifo_U_dcore_n188;
   wire FE_PHN1466_U_dfifo_U_dcore_n187;
   wire FE_PHN1465_U_dfifo_U_dcore_n192;
   wire FE_PHN1464_U_dfifo_U_dcore_n191;
   wire FE_PHN1460_U_dfifo_U_dcore_U_sub_fifo_n447;
   wire FE_PHN1459_U_dfifo_U_dcore_n189;
   wire FE_PHN1458_U_dfifo_U_dcore_n190;
   wire FE_PHN1454_U_dfifo_U_dcore_n197;
   wire FE_PHN1453_U_dfifo_U_dcore_n196;
   wire FE_PHN1452_U_dfifo_U_dcore_n195;
   wire FE_PHN1451_U_dfifo_U_dcore_n198;
   wire FE_PHN1446_U_dfifo_U_dcore_n173;
   wire FE_PHN1443_U_dfifo_U_dcore_n182;
   wire FE_PHN1442_U_dfifo_U_dcore_n172;
   wire FE_PHN1441_U_dfifo_U_dcore_n181;
   wire FE_PHN1440_U_dfifo_U_dcore_n174;
   wire FE_PHN1439_U_dfifo_U_dcore_n171;
   wire FE_PHN1438_U_dfifo_U_dcore_n176;
   wire FE_PHN1437_U_dfifo_U_dcore_n175;
   wire FE_PHN1436_U_dfifo_U_dcore_n179;
   wire FE_PHN1435_U_dfifo_U_dcore_n184;
   wire FE_PHN1434_U_dfifo_U_dcore_n183;
   wire FE_PHN1432_n13;
   wire FE_PHN1423_U_dfifo_U_dcore_m_sf_full;
   wire FE_PHN1422_U_dfifo_U_dcore_U_sub_fifo_count_1_;
   wire FE_PHN1417_U_dfifo_U_dcore_f_buf_data_1_;
   wire FE_PHN1408_U_afifo_U_acore_n173;
   wire FE_PHN1406_U_afifo_U_acore_n76;
   wire FE_PHN1405_U_afifo_U_acore_n90;
   wire FE_PHN1404_U_afifo_U_acore_n92;
   wire FE_PHN1374_U_afifo_m_data_in_12_;
   wire FE_PHN1373_U_afifo_m_data_in_42_;
   wire FE_PHN1370_U_ctl_n122;
   wire FE_PHN1368_U_ctl_n136;
   wire FE_PHN1342_U_ctl_n101;
   wire FE_PHN1332_U_afifo_U_acore_n141;
   wire FE_PHN1330_U_afifo_U_acore_n142;
   wire FE_PHN1327_U_afifo_U_acore_n144;
   wire FE_PHN1325_U_afifo_U_acore_n138;
   wire FE_PHN1324_U_afifo_U_acore_n139;
   wire FE_PHN1319_U_afifo_U_acore_n134;
   wire FE_PHN1318_U_afifo_U_acore_n140;
   wire FE_PHN1317_U_afifo_U_acore_n136;
   wire FE_PHN1316_U_afifo_U_acore_n135;
   wire FE_PHN1314_U_afifo_U_acore_n133;
   wire FE_PHN1313_U_afifo_U_acore_n148;
   wire FE_PHN1312_U_afifo_U_acore_n105;
   wire FE_PHN1309_U_afifo_U_acore_n121;
   wire FE_PHN1308_U_afifo_U_acore_n137;
   wire FE_PHN1307_U_afifo_U_acore_n110;
   wire FE_PHN1305_U_afifo_U_acore_n151;
   wire FE_PHN1304_U_afifo_U_acore_n115;
   wire FE_PHN1302_U_afifo_U_acore_n118;
   wire FE_PHN1301_U_afifo_U_acore_n147;
   wire FE_PHN1298_U_afifo_U_acore_n111;
   wire FE_PHN1297_U_afifo_U_acore_n114;
   wire FE_PHN1296_U_afifo_U_acore_n152;
   wire FE_PHN1293_U_afifo_U_acore_n112;
   wire FE_PHN1290_U_afifo_U_acore_n149;
   wire FE_PHN1289_U_afifo_U_acore_n109;
   wire FE_PHN1286_U_afifo_U_acore_n108;
   wire FE_PHN1285_U_afifo_U_acore_n117;
   wire FE_PHN1284_U_afifo_U_acore_n146;
   wire FE_PHN1282_U_afifo_U_acore_n154;
   wire FE_PHN1281_U_afifo_U_acore_n130;
   wire FE_PHN1280_U_afifo_U_acore_n107;
   wire FE_PHN1278_U_afifo_U_acore_n106;
   wire FE_PHN1277_U_afifo_U_acore_n113;
   wire FE_PHN1276_U_afifo_U_acore_n150;
   wire FE_PHN1274_U_afifo_U_acore_n126;
   wire FE_PHN1273_U_afifo_U_acore_n128;
   wire FE_PHN1272_U_afifo_U_acore_n116;
   wire FE_PHN1270_U_afifo_U_acore_n131;
   wire FE_PHN1267_U_afifo_U_acore_n127;
   wire FE_PHN1266_U_afifo_U_acore_n120;
   wire FE_PHN1265_U_afifo_U_acore_n145;
   wire FE_PHN1264_U_afifo_U_acore_n132;
   wire FE_PHN1263_U_afifo_U_acore_n124;
   wire FE_PHN1261_U_afifo_U_acore_n129;
   wire FE_PHN1260_U_afifo_U_acore_n123;
   wire FE_PHN1259_U_afifo_U_acore_n122;
   wire FE_PHN1258_U_afifo_U_acore_n125;
   wire FE_PHN1257_U_afifo_U_acore_n119;
   wire FE_PHN1250_U_dfifo_U_dcore_n200;
   wire FE_PHN1248_U_dfifo_U_dcore_n199;
   wire FE_PHN1246_U_dfifo_U_dcore_n170;
   wire FE_PHN1245_U_dfifo_U_dcore_n177;
   wire FE_PHN1244_U_dfifo_U_dcore_n185;
   wire FE_PHN1239_U_afifo_m_data_in_5_;
   wire FE_PHN1238_U_afifo_m_data_in_4_;
   wire FE_PHN1233_U_ctl_n125;
   wire FE_PHN1232_U_ctl_n124;
   wire FE_PHN1231_U_rbuf_n88;
   wire FE_PHN1229_U_ctl_n138;
   wire FE_PHN1226_U_ctl_n102;
   wire FE_PHN1225_U_ctl_n104;
   wire FE_PHN1223_U_afifo_U_acore_U_sub_fifo_n171;
   wire FE_PHN1197_U_afifo_U_acore_n72;
   wire FE_PHN1194_U_afifo_U_acore_n74;
   wire FE_PHN1193_U_afifo_U_acore_n88;
   wire FE_PHN1192_U_afifo_U_acore_n68;
   wire FE_PHN1191_U_afifo_U_acore_n78;
   wire FE_PHN1190_U_afifo_U_acore_n84;
   wire FE_PHN1189_U_afifo_U_acore_n167;
   wire FE_PHN1188_U_afifo_U_acore_n86;
   wire FE_PHN1187_U_afifo_U_acore_n82;
   wire FE_PHN1186_U_afifo_U_acore_n70;
   wire FE_PHN1184_U_dfifo_U_dcore_U_sub_fifo_n452;
   wire FE_PHN1182_U_dfifo_U_dcore_n143;
   wire FE_PHN1181_U_dfifo_U_dcore_n149;
   wire FE_PHN1180_U_dfifo_U_dcore_n146;
   wire FE_PHN1179_U_dfifo_U_dcore_n142;
   wire FE_PHN1178_U_afifo_m_data_in_32_;
   wire FE_PHN1162_U_ctl_n139;
   wire FE_PHN1132_U_dfifo_n3;
   wire FE_PHN1125_U_dfifo_U_dcore_n180;
   wire FE_PHN1115_U_rbuf_n86;
   wire FE_PHN1114_U_rbuf_n79;
   wire FE_PHN1113_U_afifo_n49;
   wire FE_PHN1112_U_rbuf_n75;
   wire FE_PHN1111_U_rbuf_n83;
   wire FE_PHN1110_U_rbuf_n80;
   wire FE_PHN1109_U_rbuf_n72;
   wire FE_PHN1108_U_rbuf_n77;
   wire FE_PHN1107_U_ctl_n134;
   wire FE_PHN1106_U_ctl_n133;
   wire FE_PHN1105_U_rbuf_n74;
   wire FE_PHN1104_U_rbuf_n78;
   wire FE_PHN1102_U_ctl_n103;
   wire FE_PHN1100_U_afifo_U_acore_U_sub_fifo_n325;
   wire FE_PHN1084_U_dfifo_U_dcore_n154;
   wire FE_PHN1079_U_ctl_n400;
   wire FE_PHN1075_U_rbuf_n63;
   wire FE_PHN1074_U_rbuf_n64;
   wire FE_PHN1073_U_rbuf_n59;
   wire FE_PHN1072_U_rbuf_n65;
   wire FE_PHN1071_U_rbuf_n67;
   wire FE_PHN1070_U_rbuf_n60;
   wire FE_PHN1069_U_rbuf_n56;
   wire FE_PHN1068_U_rbuf_n61;
   wire FE_PHN1067_U_rbuf_n57;
   wire FE_PHN1066_U_rbuf_n70;
   wire FE_PHN1065_U_rbuf_n58;
   wire FE_PHN1049_U_afifo_U_acore_U_sub_fifo_n11;
   wire FE_PHN1039_U_rbuf_n73;
   wire FE_PHN1036_U_ctl_f_hiu_terminate;
   wire FE_PHN1027_U_afifo_n2;
   wire FE_PHN1022_U_dfifo_U_dcore_n137;
   wire FE_PHN1021_U_dfifo_U_dcore_n138;
   wire FE_PHN1019_U_dfifo_U_dcore_n141;
   wire FE_PHN1018_U_dfifo_U_dcore_n134;
   wire FE_PHN1011_U_ctl_n135;
   wire FE_PHN1002_U_ctl_n100;
   wire FE_PHN999_U_ctl_fr_wr_bcnt_0_;
   wire FE_PHN993_U_afifo_U_acore_U_sub_fifo_n149;
   wire FE_PHN975_U_ctl_n132;
   wire FE_PHN962_U_afifo_U_acore_n_afull;
   wire FE_PHN956_U_dfifo_U_dcore_n147;
   wire FE_PHN954_U_dfifo_U_dcore_n150;
   wire FE_PHN950_U_afifo_n185;
   wire FE_PHN947_U_rbuf_n62;
   wire FE_PHN930_U_rbuf_n76;
   wire FE_PHN929_U_rbuf_n81;
   wire FE_PHN923_U_dfifo_U_dcore_n167;
   wire FE_PHN920_U_dfifo_U_dcore_n158;
   wire FE_PHN919_U_dfifo_U_dcore_n165;
   wire FE_PHN915_U_dfifo_U_dcore_n161;
   wire FE_PHN914_U_dfifo_U_dcore_n164;
   wire FE_PHN913_U_dfifo_U_dcore_n159;
   wire FE_PHN912_U_dfifo_U_dcore_n162;
   wire FE_PHN911_U_dfifo_U_dcore_n160;
   wire FE_PHN910_U_dfifo_U_dcore_n153;
   wire FE_PHN909_U_dfifo_U_dcore_n152;
   wire FE_PHN908_U_dfifo_U_dcore_n163;
   wire FE_PHN903_U_dfifo_U_dcore_n166;
   wire FE_PHN890_U_dfifo_U_dcore_n178;
   wire FE_PHN888_U_ctl_n150;
   wire FE_PHN885_U_ctl_n123;
   wire FE_PHN876_U_rbuf_n68;
   wire FE_PHN872_U_rbuf_n66;
   wire FE_PHN868_U_afifo_U_acore_U_sub_fifo_n172;
   wire FE_PHN867_U_afifo_U_acore_U_sub_fifo_count_1_;
   wire FE_PHN861_U_dfifo_U_dcore_n144;
   wire FE_PHN860_U_dfifo_U_dcore_n148;
   wire FE_PHN858_U_dfifo_U_dcore_n140;
   wire FE_PHN857_U_dfifo_U_dcore_n135;
   wire FE_PHN848_U_ctl_n127;
   wire FE_PHN828_U_rbuf_n69;
   wire FE_PHN827_U_rbuf_n55;
   wire FE_PHN817_U_afifo_U_acore_n2;
   wire FE_PHN815_U_afifo_U_acore_n11;
   wire FE_PHN812_U_dfifo_U_dcore_n151;
   wire FE_PHN811_U_dfifo_U_dcore_n156;
   wire FE_PHN810_U_dfifo_U_dcore_n155;
   wire FE_PHN809_U_dfifo_U_dcore_n157;
   wire FE_PHN808_U_afifo_n65;
   wire FE_PHN798_U_afifo_n259;
   wire FE_PHN795_U_ctl_n180;
   wire FE_PHN789_U_dfifo_U_dcore_U_sub_fifo_n450;
   wire FE_PHN785_U_dfifo_U_dcore_n136;
   wire FE_PHN784_U_dfifo_U_dcore_n139;
   wire FE_PHN782_U_rbuf_n89;
   wire FE_PHN761_U_afifo_U_acore_f_push_req_n;
   wire FE_PHN750_U_afifo_U_acore_n_obuf_empty;
   wire FE_PHN747_U_ctl_n335;
   wire FE_PHN744_U_ctl_n105;
   wire FE_PHN736_m_rb_overflow;
   wire FE_PHN714_miu_burst_done;
   wire FE_PHN708_U_ctl_n418;
   wire FE_PHN700_U_ctl_n297;
   wire FE_PHN699_U_ctl_n382;
   wire FE_PHN695_hsel_reg;
   wire FE_PHN687_U_ctl_n422;
   wire FE_PHN682_U_ctl_n295;
   wire FE_PHN676_hiu_terminate;
   wire FE_PHN673_m_af_push1_n;
   wire FE_OFN296_n64;
   wire FE_OFN295_n61;
   wire FE_OFN294_n60;
   wire FE_OFN292_n56;
   wire FE_OFN291_n55;
   wire FE_OFN290_n53;
   wire FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8;
   wire FE_OFN288_U_dfifo_U_dcore_U_sub_fifo_n9;
   wire FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10;
   wire FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14;
   wire FE_OFN281_U_dfifo_U_dcore_U_sub_fifo_n15;
   wire FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16;
   wire FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231;
   wire FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232;
   wire FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234;
   wire FE_OFN271_U_dfifo_U_dcore_U_sub_fifo_n560;
   wire FE_OFN267_U_dfifo_U_dcore_U_sub_fifo_n562;
   wire FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605;
   wire FE_OFN264_U_afifo_U_acore_U_sub_fifo_n152;
   wire FE_OFN263_U_afifo_U_acore_U_sub_fifo_n161;
   wire FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161;
   wire FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163;
   wire FE_OFN260_U_afifo_U_acore_U_sub_fifo_n212;
   wire FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369;
   wire FE_OFN258_U_dfifo_U_dcore_n1;
   wire FE_OFN256_U_dfifo_U_dcore_n2;
   wire FE_OFN255_U_dfifo_U_dcore_n3;
   wire FE_OFN252_U_dfifo_U_dcore_n127;
   wire FE_OFN250_U_afifo_U_acore_n1;
   wire FE_OFN247_U_afifo_U_acore_n211;
   wire FE_OFN244_U_rbuf_n180;
   wire FE_OFN237_U_afifo_n54;
   wire FE_OFN236_U_afifo_n93;
   wire FE_OFN225_hiu_data_26_;
   wire FE_OFN210_hwrite_s;
   wire FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169;
   wire FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369;
   wire FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1;
   wire FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162;
   wire FE_OFN197_U_afifo_U_acore_n38;
   wire FE_OFN196_HRESETn;
   wire FE_OFN193_HRESETn;
   wire FE_OFN176_HRESETn;
   wire FE_OFN171_HRESETn;
   wire FE_OFN170_HRESETn;
   wire FE_OFN169_HRESETn;
   wire FE_OFN168_HRESETn;
   wire FE_OFN157_HRESETn;
   wire FE_OFN156_HRESETn;
   wire FE_OFN153_HRESETn;
   wire FE_OFN150_HRESETn;
   wire FE_OFN149_HRESETn;
   wire FE_OFN143_HRESETn;
   wire FE_OFN136_HRESETn;
   wire FE_OFN69_HRESETn;
   wire FE_OFN67_HRESETn;
   wire FE_OFN62_HRESETn;
   wire FE_OFN58_HRESETn;
   wire FE_OFN54_HRESETn;
   wire FE_OFN47_HRESETn;
   wire FE_OFN32_HRESETn;
   wire FE_OFN26_U_afifo_U_acore_n38;
   wire FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162;
   wire FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1;
   wire FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169;
   wire m_af_push1_n;
   wire m_af_data1_in_13_;
   wire m_af_data1_in_11_;
   wire m_af_data1_in_5_;
   wire m_af_data1_in_4_;
   wire m_af_data1_in_2_;
   wire m_af_data1_in_0_;
   wire m_af_ready;
   wire m_af_new_req;
   wire m_af_dummy_req;
   wire m_df_push_n;
   wire m_df_ready;
   wire m_df_wr_term;
   wire m_two_to_one;
   wire m_rb_start;
   wire m_rb_pop_n;
   wire m_rb_sel_buf;
   wire m_double;
   wire m_rb_ready;
   wire m_rb_overflow;
   wire U_afifo_n259;
   wire U_afifo_n258;
   wire U_afifo_n257;
   wire U_afifo_n256;
   wire U_afifo_n255;
   wire U_afifo_n250;
   wire U_afifo_n248;
   wire U_afifo_n246;
   wire U_afifo_n245;
   wire U_afifo_n244;
   wire U_afifo_n243;
   wire U_afifo_n242;
   wire U_afifo_n241;
   wire U_afifo_n240;
   wire U_afifo_n239;
   wire U_afifo_n238;
   wire U_afifo_n237;
   wire U_afifo_n236;
   wire U_afifo_n235;
   wire U_afifo_n234;
   wire U_afifo_n233;
   wire U_afifo_n232;
   wire U_afifo_n231;
   wire U_afifo_n230;
   wire U_afifo_n229;
   wire U_afifo_n228;
   wire U_afifo_n227;
   wire U_afifo_n226;
   wire U_afifo_n225;
   wire U_afifo_n224;
   wire U_afifo_n223;
   wire U_afifo_n222;
   wire U_afifo_n221;
   wire U_afifo_n220;
   wire U_afifo_n219;
   wire U_afifo_n218;
   wire U_afifo_n217;
   wire U_afifo_n216;
   wire U_afifo_n215;
   wire U_afifo_n214;
   wire U_afifo_n213;
   wire U_afifo_n212;
   wire U_afifo_n211;
   wire U_afifo_n210;
   wire U_afifo_n209;
   wire U_afifo_n208;
   wire U_afifo_n207;
   wire U_afifo_n206;
   wire U_afifo_n205;
   wire U_afifo_n204;
   wire U_afifo_n203;
   wire U_afifo_n202;
   wire U_afifo_n201;
   wire U_afifo_n200;
   wire U_afifo_n198;
   wire U_afifo_n192;
   wire U_afifo_n191;
   wire U_afifo_n188;
   wire U_afifo_n187;
   wire U_afifo_n186;
   wire U_afifo_n185;
   wire U_afifo_n184;
   wire U_afifo_n183;
   wire U_afifo_n182;
   wire U_afifo_n181;
   wire U_afifo_n180;
   wire U_afifo_n179;
   wire U_afifo_n178;
   wire U_afifo_n173;
   wire U_afifo_n171;
   wire U_afifo_n169;
   wire U_afifo_n168;
   wire U_afifo_n167;
   wire U_afifo_n166;
   wire U_afifo_n165;
   wire U_afifo_n164;
   wire U_afifo_n163;
   wire U_afifo_n162;
   wire U_afifo_n161;
   wire U_afifo_n160;
   wire U_afifo_n159;
   wire U_afifo_n158;
   wire U_afifo_n157;
   wire U_afifo_n156;
   wire U_afifo_n155;
   wire U_afifo_n154;
   wire U_afifo_n153;
   wire U_afifo_n152;
   wire U_afifo_n151;
   wire U_afifo_n147;
   wire U_afifo_n140;
   wire U_afifo_n138;
   wire U_afifo_n137;
   wire U_afifo_n99;
   wire U_afifo_n98;
   wire U_afifo_n85;
   wire U_afifo_n84;
   wire U_afifo_n76;
   wire U_afifo_n75;
   wire U_afifo_n54;
   wire U_afifo_n49;
   wire U_afifo_n15;
   wire U_afifo_n14;
   wire U_afifo_n13;
   wire U_afifo_n11;
   wire U_afifo_n10;
   wire U_afifo_n9;
   wire U_afifo_n7;
   wire U_afifo_n5;
   wire U_afifo_n1;
   wire U_afifo_n65;
   wire U_afifo_n55;
   wire U_afifo_n52;
   wire U_afifo_n51;
   wire U_afifo_n48;
   wire U_afifo_n47;
   wire U_afifo_n46;
   wire U_afifo_n45;
   wire U_afifo_n44;
   wire U_afifo_n43;
   wire U_afifo_n42;
   wire U_afifo_n41;
   wire U_afifo_n40;
   wire U_afifo_n39;
   wire U_afifo_n38;
   wire U_afifo_n37;
   wire U_afifo_n36;
   wire U_afifo_n35;
   wire U_afifo_n34;
   wire U_afifo_n33;
   wire U_afifo_n32;
   wire U_afifo_n31;
   wire U_afifo_n30;
   wire U_afifo_n29;
   wire U_afifo_n28;
   wire U_afifo_n27;
   wire U_afifo_n26;
   wire U_afifo_n25;
   wire U_afifo_n24;
   wire U_afifo_n23;
   wire U_afifo_n22;
   wire U_afifo_n21;
   wire U_afifo_n20;
   wire U_afifo_n19;
   wire U_afifo_n18;
   wire U_afifo_n17;
   wire U_afifo_n16;
   wire U_afifo_n12;
   wire U_afifo_n8;
   wire U_afifo_n6;
   wire U_afifo_n4;
   wire U_afifo_n3;
   wire U_afifo_n2;
   wire U_afifo_n_new_req;
   wire U_afifo_f_clr_pers;
   wire U_afifo_f_core_ready;
   wire U_afifo_f_data2_0_;
   wire U_afifo_f_data2_2_;
   wire U_afifo_f_data2_4_;
   wire U_afifo_f_data2_5_;
   wire U_afifo_f_data2_6_;
   wire U_afifo_f_data2_7_;
   wire U_afifo_f_data2_8_;
   wire U_afifo_f_data2_12_;
   wire U_afifo_f_data2_13_;
   wire U_afifo_f_data2_14_;
   wire U_afifo_f_data2_15_;
   wire U_afifo_f_data2_16_;
   wire U_afifo_f_data2_17_;
   wire U_afifo_f_data2_18_;
   wire U_afifo_f_data2_19_;
   wire U_afifo_f_data2_20_;
   wire U_afifo_f_data2_21_;
   wire U_afifo_f_data2_22_;
   wire U_afifo_f_data2_23_;
   wire U_afifo_f_data2_24_;
   wire U_afifo_f_data2_25_;
   wire U_afifo_f_data2_26_;
   wire U_afifo_f_data2_27_;
   wire U_afifo_f_data2_28_;
   wire U_afifo_f_data2_29_;
   wire U_afifo_f_data2_30_;
   wire U_afifo_f_data2_31_;
   wire U_afifo_f_data2_32_;
   wire U_afifo_f_data2_33_;
   wire U_afifo_f_data2_34_;
   wire U_afifo_f_data2_35_;
   wire U_afifo_f_data2_36_;
   wire U_afifo_f_data2_37_;
   wire U_afifo_f_data2_38_;
   wire U_afifo_f_data2_39_;
   wire U_afifo_f_data2_40_;
   wire U_afifo_f_data2_41_;
   wire U_afifo_f_data2_42_;
   wire U_afifo_f_data2_43_;
   wire U_afifo_f_data2_44_;
   wire U_afifo_f_data2_47_;
   wire U_afifo_f_data2_48_;
   wire U_afifo_f_push2_pending;
   wire U_afifo_m_data_out_0_;
   wire U_afifo_m_data_out_3;
   wire U_afifo_m_data_out_49;
   wire U_afifo_m_full;
   wire U_afifo_m_afull;
   wire U_afifo_m_aempty;
   wire U_afifo_m_empty;
   wire U_afifo_m_pop_n;
   wire U_dfifo_n4;
   wire U_dfifo_n2;
   wire U_dfifo_n5;
   wire U_dfifo_n3;
   wire U_dfifo_f_1st_half;
   wire U_dfifo_m_full;
   wire U_dfifo_m_afull;
   wire U_dfifo_m_aempty;
   wire U_dfifo_m_empty;
   wire U_dfifo_m_data_out_0_;
   wire U_dfifo_m_data_out_1_;
   wire U_rbuf_n198;
   wire U_rbuf_n197;
   wire U_rbuf_n196;
   wire U_rbuf_n195;
   wire U_rbuf_n194;
   wire U_rbuf_n193;
   wire U_rbuf_n192;
   wire U_rbuf_n191;
   wire U_rbuf_n190;
   wire U_rbuf_n189;
   wire U_rbuf_n188;
   wire U_rbuf_n187;
   wire U_rbuf_n186;
   wire U_rbuf_n185;
   wire U_rbuf_n184;
   wire U_rbuf_n183;
   wire U_rbuf_n182;
   wire U_rbuf_n181;
   wire U_rbuf_n180;
   wire U_rbuf_n179;
   wire U_rbuf_n178;
   wire U_rbuf_n177;
   wire U_rbuf_n176;
   wire U_rbuf_n175;
   wire U_rbuf_n174;
   wire U_rbuf_n173;
   wire U_rbuf_n172;
   wire U_rbuf_n171;
   wire U_rbuf_n170;
   wire U_rbuf_n169;
   wire U_rbuf_n168;
   wire U_rbuf_n167;
   wire U_rbuf_n166;
   wire U_rbuf_n165;
   wire U_rbuf_n164;
   wire U_rbuf_n163;
   wire U_rbuf_n162;
   wire U_rbuf_n161;
   wire U_rbuf_n160;
   wire U_rbuf_n159;
   wire U_rbuf_n158;
   wire U_rbuf_n157;
   wire U_rbuf_n156;
   wire U_rbuf_n154;
   wire U_rbuf_n151;
   wire U_rbuf_n149;
   wire U_rbuf_n148;
   wire U_rbuf_n146;
   wire U_rbuf_n145;
   wire U_rbuf_n143;
   wire U_rbuf_n142;
   wire U_rbuf_n141;
   wire U_rbuf_n140;
   wire U_rbuf_n139;
   wire U_rbuf_n138;
   wire U_rbuf_n137;
   wire U_rbuf_n136;
   wire U_rbuf_n135;
   wire U_rbuf_n134;
   wire U_rbuf_n133;
   wire U_rbuf_n132;
   wire U_rbuf_n131;
   wire U_rbuf_n130;
   wire U_rbuf_n129;
   wire U_rbuf_n128;
   wire U_rbuf_n127;
   wire U_rbuf_n126;
   wire U_rbuf_n125;
   wire U_rbuf_n124;
   wire U_rbuf_n123;
   wire U_rbuf_n120;
   wire U_rbuf_n116;
   wire U_rbuf_n115;
   wire U_rbuf_n114;
   wire U_rbuf_n113;
   wire U_rbuf_n112;
   wire U_rbuf_n111;
   wire U_rbuf_n110;
   wire U_rbuf_n109;
   wire U_rbuf_n108;
   wire U_rbuf_n107;
   wire U_rbuf_n106;
   wire U_rbuf_n105;
   wire U_rbuf_n104;
   wire U_rbuf_n103;
   wire U_rbuf_n102;
   wire U_rbuf_n101;
   wire U_rbuf_n100;
   wire U_rbuf_n99;
   wire U_rbuf_n98;
   wire U_rbuf_n97;
   wire U_rbuf_n96;
   wire U_rbuf_n95;
   wire U_rbuf_n94;
   wire U_rbuf_n93;
   wire U_rbuf_n92;
   wire U_rbuf_n91;
   wire U_rbuf_n90;
   wire U_rbuf_n54;
   wire U_rbuf_n53;
   wire U_rbuf_n52;
   wire U_rbuf_n51;
   wire U_rbuf_n50;
   wire U_rbuf_n49;
   wire U_rbuf_n48;
   wire U_rbuf_n47;
   wire U_rbuf_n46;
   wire U_rbuf_n45;
   wire U_rbuf_n44;
   wire U_rbuf_n43;
   wire U_rbuf_n42;
   wire U_rbuf_n41;
   wire U_rbuf_n40;
   wire U_rbuf_n39;
   wire U_rbuf_n38;
   wire U_rbuf_n35;
   wire U_rbuf_n34;
   wire U_rbuf_n33;
   wire U_rbuf_n32;
   wire U_rbuf_n31;
   wire U_rbuf_n30;
   wire U_rbuf_n29;
   wire U_rbuf_n28;
   wire U_rbuf_n27;
   wire U_rbuf_n26;
   wire U_rbuf_n25;
   wire U_rbuf_n24;
   wire U_rbuf_n23;
   wire U_rbuf_n22;
   wire U_rbuf_n21;
   wire U_rbuf_n20;
   wire U_rbuf_n19;
   wire U_rbuf_n18;
   wire U_rbuf_n17;
   wire U_rbuf_n16;
   wire U_rbuf_n15;
   wire U_rbuf_n9;
   wire U_rbuf_n8;
   wire U_rbuf_n7;
   wire U_rbuf_n6;
   wire U_rbuf_n4;
   wire U_rbuf_n3;
   wire U_rbuf_n89;
   wire U_rbuf_n88;
   wire U_rbuf_n86;
   wire U_rbuf_n85;
   wire U_rbuf_n84;
   wire U_rbuf_n83;
   wire U_rbuf_n82;
   wire U_rbuf_n81;
   wire U_rbuf_n80;
   wire U_rbuf_n79;
   wire U_rbuf_n78;
   wire U_rbuf_n77;
   wire U_rbuf_n76;
   wire U_rbuf_n75;
   wire U_rbuf_n74;
   wire U_rbuf_n73;
   wire U_rbuf_n72;
   wire U_rbuf_n71;
   wire U_rbuf_n70;
   wire U_rbuf_n69;
   wire U_rbuf_n68;
   wire U_rbuf_n67;
   wire U_rbuf_n66;
   wire U_rbuf_n65;
   wire U_rbuf_n64;
   wire U_rbuf_n63;
   wire U_rbuf_n62;
   wire U_rbuf_n61;
   wire U_rbuf_n60;
   wire U_rbuf_n59;
   wire U_rbuf_n58;
   wire U_rbuf_n57;
   wire U_rbuf_n56;
   wire U_rbuf_n55;
   wire U_rbuf_f_top_data_0_;
   wire U_rbuf_f_top_data_1_;
   wire U_rbuf_f_top_data_2_;
   wire U_rbuf_f_top_data_3_;
   wire U_rbuf_f_top_data_4_;
   wire U_rbuf_f_top_data_5_;
   wire U_rbuf_f_top_data_6_;
   wire U_rbuf_f_top_data_7_;
   wire U_rbuf_f_top_data_8_;
   wire U_rbuf_f_top_data_9_;
   wire U_rbuf_f_top_data_10_;
   wire U_rbuf_f_top_data_11_;
   wire U_rbuf_f_top_data_12_;
   wire U_rbuf_f_top_data_13_;
   wire U_rbuf_f_top_data_14_;
   wire U_rbuf_f_top_data_15_;
   wire U_rbuf_f_1st_half;
   wire U_rbuf_f_rbuf_state_0_;
   wire U_rbuf_f_rbuf_state_1_;
   wire U_ctl_n422;
   wire U_ctl_n421;
   wire U_ctl_n420;
   wire U_ctl_n419;
   wire U_ctl_n418;
   wire U_ctl_n417;
   wire U_ctl_n416;
   wire U_ctl_n415;
   wire U_ctl_n414;
   wire U_ctl_n413;
   wire U_ctl_n412;
   wire U_ctl_n411;
   wire U_ctl_n410;
   wire U_ctl_n409;
   wire U_ctl_n408;
   wire U_ctl_n407;
   wire U_ctl_n406;
   wire U_ctl_n405;
   wire U_ctl_n404;
   wire U_ctl_n403;
   wire U_ctl_n402;
   wire U_ctl_n401;
   wire U_ctl_n400;
   wire U_ctl_n398;
   wire U_ctl_n395;
   wire U_ctl_n394;
   wire U_ctl_n392;
   wire U_ctl_n391;
   wire U_ctl_n390;
   wire U_ctl_n389;
   wire U_ctl_n388;
   wire U_ctl_n387;
   wire U_ctl_n386;
   wire U_ctl_n385;
   wire U_ctl_n384;
   wire U_ctl_n383;
   wire U_ctl_n382;
   wire U_ctl_n380;
   wire U_ctl_n379;
   wire U_ctl_n378;
   wire U_ctl_n376;
   wire U_ctl_n375;
   wire U_ctl_n374;
   wire U_ctl_n373;
   wire U_ctl_n372;
   wire U_ctl_n371;
   wire U_ctl_n370;
   wire U_ctl_n369;
   wire U_ctl_n368;
   wire U_ctl_n367;
   wire U_ctl_n366;
   wire U_ctl_n365;
   wire U_ctl_n364;
   wire U_ctl_n363;
   wire U_ctl_n362;
   wire U_ctl_n361;
   wire U_ctl_n360;
   wire U_ctl_n359;
   wire U_ctl_n358;
   wire U_ctl_n357;
   wire U_ctl_n356;
   wire U_ctl_n355;
   wire U_ctl_n354;
   wire U_ctl_n353;
   wire U_ctl_n352;
   wire U_ctl_n351;
   wire U_ctl_n350;
   wire U_ctl_n349;
   wire U_ctl_n348;
   wire U_ctl_n347;
   wire U_ctl_n346;
   wire U_ctl_n345;
   wire U_ctl_n343;
   wire U_ctl_n342;
   wire U_ctl_n341;
   wire U_ctl_n340;
   wire U_ctl_n339;
   wire U_ctl_n337;
   wire U_ctl_n336;
   wire U_ctl_n335;
   wire U_ctl_n331;
   wire U_ctl_n330;
   wire U_ctl_n329;
   wire U_ctl_n328;
   wire U_ctl_n327;
   wire U_ctl_n326;
   wire U_ctl_n325;
   wire U_ctl_n324;
   wire U_ctl_n323;
   wire U_ctl_n318;
   wire U_ctl_n317;
   wire U_ctl_n316;
   wire U_ctl_n315;
   wire U_ctl_n314;
   wire U_ctl_n313;
   wire U_ctl_n312;
   wire U_ctl_n311;
   wire U_ctl_n310;
   wire U_ctl_n309;
   wire U_ctl_n308;
   wire U_ctl_n307;
   wire U_ctl_n306;
   wire U_ctl_n305;
   wire U_ctl_n304;
   wire U_ctl_n301;
   wire U_ctl_n297;
   wire U_ctl_n296;
   wire U_ctl_n295;
   wire U_ctl_n294;
   wire U_ctl_n293;
   wire U_ctl_n292;
   wire U_ctl_n290;
   wire U_ctl_n289;
   wire U_ctl_n288;
   wire U_ctl_n276;
   wire U_ctl_n269;
   wire U_ctl_n267;
   wire U_ctl_n252;
   wire U_ctl_n251;
   wire U_ctl_n250;
   wire U_ctl_n248;
   wire U_ctl_n235;
   wire U_ctl_n230;
   wire U_ctl_n227;
   wire U_ctl_n225;
   wire U_ctl_n222;
   wire U_ctl_n221;
   wire U_ctl_n220;
   wire U_ctl_n214;
   wire U_ctl_n212;
   wire U_ctl_n211;
   wire U_ctl_n210;
   wire U_ctl_n209;
   wire U_ctl_n208;
   wire U_ctl_n202;
   wire U_ctl_n201;
   wire U_ctl_n200;
   wire U_ctl_n199;
   wire U_ctl_n198;
   wire U_ctl_n197;
   wire U_ctl_n196;
   wire U_ctl_n195;
   wire U_ctl_n194;
   wire U_ctl_n193;
   wire U_ctl_n187;
   wire U_ctl_n186;
   wire U_ctl_n183;
   wire U_ctl_n180;
   wire U_ctl_n174;
   wire U_ctl_n173;
   wire U_ctl_n171;
   wire U_ctl_n170;
   wire U_ctl_n169;
   wire U_ctl_n168;
   wire U_ctl_n167;
   wire U_ctl_n166;
   wire U_ctl_n160;
   wire U_ctl_n158;
   wire U_ctl_n156;
   wire U_ctl_n154;
   wire U_ctl_n151;
   wire U_ctl_n150;
   wire U_ctl_n148;
   wire U_ctl_n147;
   wire U_ctl_n146;
   wire U_ctl_n145;
   wire U_ctl_n144;
   wire U_ctl_n143;
   wire U_ctl_n142;
   wire U_ctl_n126;
   wire U_ctl_n99;
   wire U_ctl_n98;
   wire U_ctl_n97;
   wire U_ctl_n96;
   wire U_ctl_n95;
   wire U_ctl_n92;
   wire U_ctl_n91;
   wire U_ctl_n89;
   wire U_ctl_n88;
   wire U_ctl_n87;
   wire U_ctl_n85;
   wire U_ctl_n63;
   wire U_ctl_n58;
   wire U_ctl_n57;
   wire U_ctl_n56;
   wire U_ctl_n55;
   wire U_ctl_n54;
   wire U_ctl_n50;
   wire U_ctl_n47;
   wire U_ctl_n45;
   wire U_ctl_n44;
   wire U_ctl_n43;
   wire U_ctl_n42;
   wire U_ctl_n41;
   wire U_ctl_n40;
   wire U_ctl_n39;
   wire U_ctl_n38;
   wire U_ctl_n36;
   wire U_ctl_n35;
   wire U_ctl_n30;
   wire U_ctl_n29;
   wire U_ctl_n28;
   wire U_ctl_n21;
   wire U_ctl_n20;
   wire U_ctl_n19;
   wire U_ctl_n16;
   wire U_ctl_n15;
   wire U_ctl_n14;
   wire U_ctl_n13;
   wire U_ctl_n11;
   wire U_ctl_n6;
   wire U_ctl_n3;
   wire U_ctl_DP_OP_140_125_8947_n1;
   wire U_ctl_DP_OP_140_125_8947_n2;
   wire U_ctl_DP_OP_140_125_8947_n3;
   wire U_ctl_DP_OP_140_125_8947_n4;
   wire U_ctl_DP_OP_140_125_8947_n5;
   wire U_ctl_DP_OP_140_125_8947_n6;
   wire U_ctl_DP_OP_140_125_8947_n7;
   wire U_ctl_DP_OP_140_125_8947_n8;
   wire U_ctl_DP_OP_140_125_8947_n9;
   wire U_ctl_DP_OP_140_125_8947_n10;
   wire U_ctl_DP_OP_140_125_8947_n11;
   wire U_ctl_DP_OP_140_125_8947_n12;
   wire U_ctl_DP_OP_140_125_8947_n13;
   wire U_ctl_DP_OP_140_125_8947_n14;
   wire U_ctl_DP_OP_140_125_8947_n15;
   wire U_ctl_DP_OP_140_125_8947_n16;
   wire U_ctl_DP_OP_140_125_8947_n17;
   wire U_ctl_DP_OP_140_125_8947_n18;
   wire U_ctl_DP_OP_140_125_8947_n19;
   wire U_ctl_DP_OP_140_125_8947_n20;
   wire U_ctl_DP_OP_140_125_8947_n22;
   wire U_ctl_DP_OP_140_125_8947_n23;
   wire U_ctl_DP_OP_140_125_8947_n24;
   wire U_ctl_DP_OP_140_125_8947_n30;
   wire U_ctl_DP_OP_140_125_8947_n31;
   wire U_ctl_DP_OP_140_125_8947_n32;
   wire U_ctl_DP_OP_140_125_8947_n33;
   wire U_ctl_DP_OP_140_125_8947_n34;
   wire U_ctl_DP_OP_140_125_8947_n35;
   wire U_ctl_DP_OP_140_125_8947_I2;
   wire U_ctl_n299;
   wire U_ctl_n141;
   wire U_ctl_n140;
   wire U_ctl_n139;
   wire U_ctl_n138;
   wire U_ctl_n137;
   wire U_ctl_n136;
   wire U_ctl_n135;
   wire U_ctl_n134;
   wire U_ctl_n133;
   wire U_ctl_n132;
   wire U_ctl_n131;
   wire U_ctl_n130;
   wire U_ctl_n129;
   wire U_ctl_n128;
   wire U_ctl_n127;
   wire U_ctl_n125;
   wire U_ctl_n124;
   wire U_ctl_n123;
   wire U_ctl_n122;
   wire U_ctl_n120;
   wire U_ctl_n119;
   wire U_ctl_n118;
   wire U_ctl_n117;
   wire U_ctl_n116;
   wire U_ctl_n106;
   wire U_ctl_n105;
   wire U_ctl_n104;
   wire U_ctl_n103;
   wire U_ctl_n102;
   wire U_ctl_n101;
   wire U_ctl_n100;
   wire U_ctl_C64_DATA2_5;
   wire U_ctl_C64_DATA2_0;
   wire U_ctl_f_burst_done;
   wire U_ctl_f_burst_done2;
   wire U_ctl_n_sel_buf;
   wire U_ctl_N288;
   wire U_ctl_N287;
   wire U_ctl_N286;
   wire U_ctl_N285;
   wire U_ctl_N284;
   wire U_ctl_f_hiu_terminate;
   wire U_ctl_fr_wr_bcnt_0_;
   wire U_ctl_fr_wr_bcnt_1_;
   wire U_ctl_fr_wr_bcnt_2_;
   wire U_ctl_fr_wr_bcnt_3_;
   wire U_ctl_fr_wr_bcnt_4_;
   wire U_ctl_fr_wr_bcnt_5_;
   wire U_ctl_N237;
   wire U_ctl_fr_prv_1wrap_tm;
   wire U_ctl_fr_prv_1wrap;
   wire U_ctl_N236;
   wire U_ctl_f_bh_state_0_;
   wire U_ctl_f_bh_state_1_;
   wire U_ctl_f_bh_state_2_;
   wire U_ctl_fd_rd_ready;
   wire U_ctl_fd_amba_bcnt_0_;
   wire U_ctl_fd_amba_bcnt_1_;
   wire U_ctl_fd_amba_bcnt_2_;
   wire U_ctl_fd_amba_bcnt_3_;
   wire U_ctl_N89;
   wire U_ctl_fd_rd_bz;
   wire U_ctl_fd_haddr_1_;
   wire U_ctl_fd_narrow_trans;
   wire U_ctl_fd_non_single;
   wire U_ctl_fd_incr;
   wire U_ctl_fd_miu_data_width_0_;
   wire U_ctl_fd_miu_data_width_1_;
   wire U_ctl_fd_miu_col_width_0_;
   wire U_ctl_fd_miu_col_width_1_;
   wire U_ctl_fd_miu_col_width_2_;
   wire U_ctl_fd_miu_col_width_3_;
   wire U_ctl_f_data_width_0_;
   wire U_ctl_fd_wr_width;
   wire U_afifo_U_acore_n211;
   wire U_afifo_U_acore_n210;
   wire U_afifo_U_acore_n209;
   wire U_afifo_U_acore_n208;
   wire U_afifo_U_acore_n207;
   wire U_afifo_U_acore_n206;
   wire U_afifo_U_acore_n205;
   wire U_afifo_U_acore_n204;
   wire U_afifo_U_acore_n203;
   wire U_afifo_U_acore_n202;
   wire U_afifo_U_acore_n201;
   wire U_afifo_U_acore_n200;
   wire U_afifo_U_acore_n199;
   wire U_afifo_U_acore_n198;
   wire U_afifo_U_acore_n197;
   wire U_afifo_U_acore_n196;
   wire U_afifo_U_acore_n195;
   wire U_afifo_U_acore_n194;
   wire U_afifo_U_acore_n193;
   wire U_afifo_U_acore_n192;
   wire U_afifo_U_acore_n191;
   wire U_afifo_U_acore_n190;
   wire U_afifo_U_acore_n189;
   wire U_afifo_U_acore_n188;
   wire U_afifo_U_acore_n187;
   wire U_afifo_U_acore_n186;
   wire U_afifo_U_acore_n185;
   wire U_afifo_U_acore_n184;
   wire U_afifo_U_acore_n183;
   wire U_afifo_U_acore_n182;
   wire U_afifo_U_acore_n181;
   wire U_afifo_U_acore_n180;
   wire U_afifo_U_acore_n179;
   wire U_afifo_U_acore_n178;
   wire U_afifo_U_acore_n177;
   wire U_afifo_U_acore_n176;
   wire U_afifo_U_acore_n175;
   wire U_afifo_U_acore_n174;
   wire U_afifo_U_acore_n173;
   wire U_afifo_U_acore_n172;
   wire U_afifo_U_acore_n171;
   wire U_afifo_U_acore_n170;
   wire U_afifo_U_acore_n169;
   wire U_afifo_U_acore_n168;
   wire U_afifo_U_acore_n167;
   wire U_afifo_U_acore_n164;
   wire U_afifo_U_acore_n163;
   wire U_afifo_U_acore_n162;
   wire U_afifo_U_acore_n161;
   wire U_afifo_U_acore_n160;
   wire U_afifo_U_acore_n159;
   wire U_afifo_U_acore_n158;
   wire U_afifo_U_acore_n157;
   wire U_afifo_U_acore_n156;
   wire U_afifo_U_acore_n155;
   wire U_afifo_U_acore_n153;
   wire U_afifo_U_acore_n143;
   wire U_afifo_U_acore_n104;
   wire U_afifo_U_acore_n103;
   wire U_afifo_U_acore_n102;
   wire U_afifo_U_acore_n101;
   wire U_afifo_U_acore_n100;
   wire U_afifo_U_acore_n99;
   wire U_afifo_U_acore_n98;
   wire U_afifo_U_acore_n97;
   wire U_afifo_U_acore_n96;
   wire U_afifo_U_acore_n95;
   wire U_afifo_U_acore_n94;
   wire U_afifo_U_acore_n93;
   wire U_afifo_U_acore_n92;
   wire U_afifo_U_acore_n91;
   wire U_afifo_U_acore_n90;
   wire U_afifo_U_acore_n89;
   wire U_afifo_U_acore_n88;
   wire U_afifo_U_acore_n87;
   wire U_afifo_U_acore_n86;
   wire U_afifo_U_acore_n85;
   wire U_afifo_U_acore_n84;
   wire U_afifo_U_acore_n83;
   wire U_afifo_U_acore_n82;
   wire U_afifo_U_acore_n81;
   wire U_afifo_U_acore_n80;
   wire U_afifo_U_acore_n79;
   wire U_afifo_U_acore_n78;
   wire U_afifo_U_acore_n77;
   wire U_afifo_U_acore_n76;
   wire U_afifo_U_acore_n75;
   wire U_afifo_U_acore_n74;
   wire U_afifo_U_acore_n73;
   wire U_afifo_U_acore_n72;
   wire U_afifo_U_acore_n71;
   wire U_afifo_U_acore_n70;
   wire U_afifo_U_acore_n69;
   wire U_afifo_U_acore_n68;
   wire U_afifo_U_acore_n67;
   wire U_afifo_U_acore_n66;
   wire U_afifo_U_acore_n65;
   wire U_afifo_U_acore_n64;
   wire U_afifo_U_acore_n63;
   wire U_afifo_U_acore_n62;
   wire U_afifo_U_acore_n61;
   wire U_afifo_U_acore_n60;
   wire U_afifo_U_acore_n59;
   wire U_afifo_U_acore_n58;
   wire U_afifo_U_acore_n57;
   wire U_afifo_U_acore_n56;
   wire U_afifo_U_acore_n55;
   wire U_afifo_U_acore_n54;
   wire U_afifo_U_acore_n53;
   wire U_afifo_U_acore_n51;
   wire U_afifo_U_acore_n49;
   wire U_afifo_U_acore_n48;
   wire U_afifo_U_acore_n47;
   wire U_afifo_U_acore_n46;
   wire U_afifo_U_acore_n45;
   wire U_afifo_U_acore_n44;
   wire U_afifo_U_acore_n43;
   wire U_afifo_U_acore_n40;
   wire U_afifo_U_acore_n39;
   wire U_afifo_U_acore_n38;
   wire U_afifo_U_acore_n34;
   wire U_afifo_U_acore_n33;
   wire U_afifo_U_acore_n32;
   wire U_afifo_U_acore_n31;
   wire U_afifo_U_acore_n30;
   wire U_afifo_U_acore_n29;
   wire U_afifo_U_acore_n28;
   wire U_afifo_U_acore_n27;
   wire U_afifo_U_acore_n26;
   wire U_afifo_U_acore_n25;
   wire U_afifo_U_acore_n24;
   wire U_afifo_U_acore_n23;
   wire U_afifo_U_acore_n22;
   wire U_afifo_U_acore_n21;
   wire U_afifo_U_acore_n20;
   wire U_afifo_U_acore_n19;
   wire U_afifo_U_acore_n18;
   wire U_afifo_U_acore_n17;
   wire U_afifo_U_acore_n16;
   wire U_afifo_U_acore_n15;
   wire U_afifo_U_acore_n14;
   wire U_afifo_U_acore_n13;
   wire U_afifo_U_acore_n12;
   wire U_afifo_U_acore_n11;
   wire U_afifo_U_acore_n10;
   wire U_afifo_U_acore_n9;
   wire U_afifo_U_acore_n8;
   wire U_afifo_U_acore_n7;
   wire U_afifo_U_acore_n6;
   wire U_afifo_U_acore_n5;
   wire U_afifo_U_acore_n4;
   wire U_afifo_U_acore_n3;
   wire U_afifo_U_acore_n2;
   wire U_afifo_U_acore_n1;
   wire U_afifo_U_acore_n166;
   wire U_afifo_U_acore_n165;
   wire U_afifo_U_acore_n154;
   wire U_afifo_U_acore_n152;
   wire U_afifo_U_acore_n151;
   wire U_afifo_U_acore_n150;
   wire U_afifo_U_acore_n149;
   wire U_afifo_U_acore_n148;
   wire U_afifo_U_acore_n147;
   wire U_afifo_U_acore_n146;
   wire U_afifo_U_acore_n145;
   wire U_afifo_U_acore_n144;
   wire U_afifo_U_acore_n142;
   wire U_afifo_U_acore_n141;
   wire U_afifo_U_acore_n140;
   wire U_afifo_U_acore_n139;
   wire U_afifo_U_acore_n138;
   wire U_afifo_U_acore_n137;
   wire U_afifo_U_acore_n136;
   wire U_afifo_U_acore_n135;
   wire U_afifo_U_acore_n134;
   wire U_afifo_U_acore_n133;
   wire U_afifo_U_acore_n132;
   wire U_afifo_U_acore_n131;
   wire U_afifo_U_acore_n130;
   wire U_afifo_U_acore_n129;
   wire U_afifo_U_acore_n128;
   wire U_afifo_U_acore_n127;
   wire U_afifo_U_acore_n126;
   wire U_afifo_U_acore_n125;
   wire U_afifo_U_acore_n124;
   wire U_afifo_U_acore_n123;
   wire U_afifo_U_acore_n122;
   wire U_afifo_U_acore_n121;
   wire U_afifo_U_acore_n120;
   wire U_afifo_U_acore_n119;
   wire U_afifo_U_acore_n118;
   wire U_afifo_U_acore_n117;
   wire U_afifo_U_acore_n116;
   wire U_afifo_U_acore_n115;
   wire U_afifo_U_acore_n114;
   wire U_afifo_U_acore_n113;
   wire U_afifo_U_acore_n112;
   wire U_afifo_U_acore_n111;
   wire U_afifo_U_acore_n110;
   wire U_afifo_U_acore_n109;
   wire U_afifo_U_acore_n108;
   wire U_afifo_U_acore_n107;
   wire U_afifo_U_acore_n106;
   wire U_afifo_U_acore_n105;
   wire U_afifo_U_acore_n_afull;
   wire U_afifo_U_acore_f_afull;
   wire U_afifo_U_acore_n_obuf_empty;
   wire U_afifo_U_acore_f_obuf_0_;
   wire U_afifo_U_acore_f_obuf_2_;
   wire U_afifo_U_acore_f_obuf_3_;
   wire U_afifo_U_acore_f_obuf_4_;
   wire U_afifo_U_acore_f_obuf_5_;
   wire U_afifo_U_acore_f_obuf_6_;
   wire U_afifo_U_acore_f_obuf_7_;
   wire U_afifo_U_acore_f_obuf_8_;
   wire U_afifo_U_acore_f_obuf_9_;
   wire U_afifo_U_acore_f_obuf_11_;
   wire U_afifo_U_acore_f_obuf_12_;
   wire U_afifo_U_acore_f_obuf_13_;
   wire U_afifo_U_acore_f_obuf_14_;
   wire U_afifo_U_acore_f_obuf_15_;
   wire U_afifo_U_acore_f_obuf_16_;
   wire U_afifo_U_acore_f_obuf_17_;
   wire U_afifo_U_acore_f_obuf_18_;
   wire U_afifo_U_acore_f_obuf_19_;
   wire U_afifo_U_acore_f_obuf_20_;
   wire U_afifo_U_acore_f_obuf_21_;
   wire U_afifo_U_acore_f_obuf_22_;
   wire U_afifo_U_acore_f_obuf_23_;
   wire U_afifo_U_acore_f_obuf_24_;
   wire U_afifo_U_acore_f_obuf_25_;
   wire U_afifo_U_acore_f_obuf_26_;
   wire U_afifo_U_acore_f_obuf_27_;
   wire U_afifo_U_acore_f_obuf_28_;
   wire U_afifo_U_acore_f_obuf_29_;
   wire U_afifo_U_acore_f_obuf_30_;
   wire U_afifo_U_acore_f_obuf_31_;
   wire U_afifo_U_acore_f_obuf_32_;
   wire U_afifo_U_acore_f_obuf_33_;
   wire U_afifo_U_acore_f_obuf_34_;
   wire U_afifo_U_acore_f_obuf_35_;
   wire U_afifo_U_acore_f_obuf_36_;
   wire U_afifo_U_acore_f_obuf_37_;
   wire U_afifo_U_acore_f_obuf_38_;
   wire U_afifo_U_acore_f_obuf_39_;
   wire U_afifo_U_acore_f_obuf_40_;
   wire U_afifo_U_acore_f_obuf_41_;
   wire U_afifo_U_acore_f_obuf_42_;
   wire U_afifo_U_acore_f_obuf_43_;
   wire U_afifo_U_acore_f_obuf_44_;
   wire U_afifo_U_acore_f_obuf_45_;
   wire U_afifo_U_acore_f_obuf_46_;
   wire U_afifo_U_acore_f_obuf_47_;
   wire U_afifo_U_acore_f_obuf_48_;
   wire U_afifo_U_acore_f_obuf_49_;
   wire U_afifo_U_acore_f_push_req_n;
   wire U_afifo_U_acore_m_sf_full;
   wire U_afifo_U_acore_f_ibuf_2_;
   wire U_afifo_U_acore_f_ibuf_18_;
   wire U_afifo_U_acore_f_ibuf_30_;
   wire U_afifo_U_acore_f_ibuf_31_;
   wire U_afifo_U_acore_f_ibuf_32_;
   wire U_afifo_U_acore_f_ibuf_33_;
   wire U_afifo_U_acore_f_ibuf_34_;
   wire U_afifo_U_acore_f_ibuf_35_;
   wire U_afifo_U_acore_f_ibuf_36_;
   wire U_afifo_U_acore_f_ibuf_37_;
   wire U_afifo_U_acore_f_ibuf_38_;
   wire U_afifo_U_acore_f_ibuf_39_;
   wire U_afifo_U_acore_f_ibuf_40_;
   wire U_afifo_U_acore_f_ibuf_41_;
   wire U_dfifo_U_dcore_n234;
   wire U_dfifo_U_dcore_n233;
   wire U_dfifo_U_dcore_n232;
   wire U_dfifo_U_dcore_n231;
   wire U_dfifo_U_dcore_n230;
   wire U_dfifo_U_dcore_n229;
   wire U_dfifo_U_dcore_n228;
   wire U_dfifo_U_dcore_n227;
   wire U_dfifo_U_dcore_n226;
   wire U_dfifo_U_dcore_n225;
   wire U_dfifo_U_dcore_n224;
   wire U_dfifo_U_dcore_n223;
   wire U_dfifo_U_dcore_n222;
   wire U_dfifo_U_dcore_n221;
   wire U_dfifo_U_dcore_n220;
   wire U_dfifo_U_dcore_n219;
   wire U_dfifo_U_dcore_n218;
   wire U_dfifo_U_dcore_n217;
   wire U_dfifo_U_dcore_n216;
   wire U_dfifo_U_dcore_n215;
   wire U_dfifo_U_dcore_n214;
   wire U_dfifo_U_dcore_n213;
   wire U_dfifo_U_dcore_n212;
   wire U_dfifo_U_dcore_n211;
   wire U_dfifo_U_dcore_n210;
   wire U_dfifo_U_dcore_n207;
   wire U_dfifo_U_dcore_n206;
   wire U_dfifo_U_dcore_n205;
   wire U_dfifo_U_dcore_n204;
   wire U_dfifo_U_dcore_n202;
   wire U_dfifo_U_dcore_n133;
   wire U_dfifo_U_dcore_n132;
   wire U_dfifo_U_dcore_n131;
   wire U_dfifo_U_dcore_n130;
   wire U_dfifo_U_dcore_n129;
   wire U_dfifo_U_dcore_n128;
   wire U_dfifo_U_dcore_n127;
   wire U_dfifo_U_dcore_n126;
   wire U_dfifo_U_dcore_n125;
   wire U_dfifo_U_dcore_n124;
   wire U_dfifo_U_dcore_n123;
   wire U_dfifo_U_dcore_n122;
   wire U_dfifo_U_dcore_n121;
   wire U_dfifo_U_dcore_n120;
   wire U_dfifo_U_dcore_n119;
   wire U_dfifo_U_dcore_n118;
   wire U_dfifo_U_dcore_n117;
   wire U_dfifo_U_dcore_n116;
   wire U_dfifo_U_dcore_n115;
   wire U_dfifo_U_dcore_n114;
   wire U_dfifo_U_dcore_n113;
   wire U_dfifo_U_dcore_n112;
   wire U_dfifo_U_dcore_n111;
   wire U_dfifo_U_dcore_n110;
   wire U_dfifo_U_dcore_n109;
   wire U_dfifo_U_dcore_n108;
   wire U_dfifo_U_dcore_n107;
   wire U_dfifo_U_dcore_n106;
   wire U_dfifo_U_dcore_n105;
   wire U_dfifo_U_dcore_n104;
   wire U_dfifo_U_dcore_n103;
   wire U_dfifo_U_dcore_n102;
   wire U_dfifo_U_dcore_n101;
   wire U_dfifo_U_dcore_n100;
   wire U_dfifo_U_dcore_n99;
   wire U_dfifo_U_dcore_n98;
   wire U_dfifo_U_dcore_n97;
   wire U_dfifo_U_dcore_n96;
   wire U_dfifo_U_dcore_n95;
   wire U_dfifo_U_dcore_n94;
   wire U_dfifo_U_dcore_n93;
   wire U_dfifo_U_dcore_n92;
   wire U_dfifo_U_dcore_n91;
   wire U_dfifo_U_dcore_n90;
   wire U_dfifo_U_dcore_n89;
   wire U_dfifo_U_dcore_n88;
   wire U_dfifo_U_dcore_n87;
   wire U_dfifo_U_dcore_n86;
   wire U_dfifo_U_dcore_n85;
   wire U_dfifo_U_dcore_n84;
   wire U_dfifo_U_dcore_n83;
   wire U_dfifo_U_dcore_n82;
   wire U_dfifo_U_dcore_n81;
   wire U_dfifo_U_dcore_n80;
   wire U_dfifo_U_dcore_n79;
   wire U_dfifo_U_dcore_n78;
   wire U_dfifo_U_dcore_n77;
   wire U_dfifo_U_dcore_n76;
   wire U_dfifo_U_dcore_n75;
   wire U_dfifo_U_dcore_n74;
   wire U_dfifo_U_dcore_n73;
   wire U_dfifo_U_dcore_n72;
   wire U_dfifo_U_dcore_n71;
   wire U_dfifo_U_dcore_n70;
   wire U_dfifo_U_dcore_n69;
   wire U_dfifo_U_dcore_n68;
   wire U_dfifo_U_dcore_n67;
   wire U_dfifo_U_dcore_n66;
   wire U_dfifo_U_dcore_n65;
   wire U_dfifo_U_dcore_n64;
   wire U_dfifo_U_dcore_n63;
   wire U_dfifo_U_dcore_n62;
   wire U_dfifo_U_dcore_n61;
   wire U_dfifo_U_dcore_n60;
   wire U_dfifo_U_dcore_n59;
   wire U_dfifo_U_dcore_n58;
   wire U_dfifo_U_dcore_n57;
   wire U_dfifo_U_dcore_n56;
   wire U_dfifo_U_dcore_n55;
   wire U_dfifo_U_dcore_n54;
   wire U_dfifo_U_dcore_n53;
   wire U_dfifo_U_dcore_n52;
   wire U_dfifo_U_dcore_n51;
   wire U_dfifo_U_dcore_n50;
   wire U_dfifo_U_dcore_n49;
   wire U_dfifo_U_dcore_n48;
   wire U_dfifo_U_dcore_n47;
   wire U_dfifo_U_dcore_n46;
   wire U_dfifo_U_dcore_n45;
   wire U_dfifo_U_dcore_n44;
   wire U_dfifo_U_dcore_n43;
   wire U_dfifo_U_dcore_n42;
   wire U_dfifo_U_dcore_n41;
   wire U_dfifo_U_dcore_n40;
   wire U_dfifo_U_dcore_n39;
   wire U_dfifo_U_dcore_n38;
   wire U_dfifo_U_dcore_n37;
   wire U_dfifo_U_dcore_n36;
   wire U_dfifo_U_dcore_n35;
   wire U_dfifo_U_dcore_n34;
   wire U_dfifo_U_dcore_n33;
   wire U_dfifo_U_dcore_n32;
   wire U_dfifo_U_dcore_n31;
   wire U_dfifo_U_dcore_n30;
   wire U_dfifo_U_dcore_n29;
   wire U_dfifo_U_dcore_n28;
   wire U_dfifo_U_dcore_n27;
   wire U_dfifo_U_dcore_n26;
   wire U_dfifo_U_dcore_n25;
   wire U_dfifo_U_dcore_n24;
   wire U_dfifo_U_dcore_n23;
   wire U_dfifo_U_dcore_n22;
   wire U_dfifo_U_dcore_n21;
   wire U_dfifo_U_dcore_n20;
   wire U_dfifo_U_dcore_n19;
   wire U_dfifo_U_dcore_n18;
   wire U_dfifo_U_dcore_n17;
   wire U_dfifo_U_dcore_n16;
   wire U_dfifo_U_dcore_n15;
   wire U_dfifo_U_dcore_n14;
   wire U_dfifo_U_dcore_n13;
   wire U_dfifo_U_dcore_n12;
   wire U_dfifo_U_dcore_n11;
   wire U_dfifo_U_dcore_n10;
   wire U_dfifo_U_dcore_n9;
   wire U_dfifo_U_dcore_n8;
   wire U_dfifo_U_dcore_n7;
   wire U_dfifo_U_dcore_n6;
   wire U_dfifo_U_dcore_n5;
   wire U_dfifo_U_dcore_n4;
   wire U_dfifo_U_dcore_n3;
   wire U_dfifo_U_dcore_n2;
   wire U_dfifo_U_dcore_n1;
   wire U_dfifo_U_dcore_n209;
   wire U_dfifo_U_dcore_n208;
   wire U_dfifo_U_dcore_n203;
   wire U_dfifo_U_dcore_n201;
   wire U_dfifo_U_dcore_n200;
   wire U_dfifo_U_dcore_n199;
   wire U_dfifo_U_dcore_n198;
   wire U_dfifo_U_dcore_n197;
   wire U_dfifo_U_dcore_n196;
   wire U_dfifo_U_dcore_n195;
   wire U_dfifo_U_dcore_n194;
   wire U_dfifo_U_dcore_n193;
   wire U_dfifo_U_dcore_n192;
   wire U_dfifo_U_dcore_n191;
   wire U_dfifo_U_dcore_n190;
   wire U_dfifo_U_dcore_n189;
   wire U_dfifo_U_dcore_n188;
   wire U_dfifo_U_dcore_n187;
   wire U_dfifo_U_dcore_n186;
   wire U_dfifo_U_dcore_n185;
   wire U_dfifo_U_dcore_n184;
   wire U_dfifo_U_dcore_n183;
   wire U_dfifo_U_dcore_n182;
   wire U_dfifo_U_dcore_n181;
   wire U_dfifo_U_dcore_n180;
   wire U_dfifo_U_dcore_n179;
   wire U_dfifo_U_dcore_n178;
   wire U_dfifo_U_dcore_n177;
   wire U_dfifo_U_dcore_n176;
   wire U_dfifo_U_dcore_n175;
   wire U_dfifo_U_dcore_n174;
   wire U_dfifo_U_dcore_n173;
   wire U_dfifo_U_dcore_n172;
   wire U_dfifo_U_dcore_n171;
   wire U_dfifo_U_dcore_n170;
   wire U_dfifo_U_dcore_n169;
   wire U_dfifo_U_dcore_n168;
   wire U_dfifo_U_dcore_n167;
   wire U_dfifo_U_dcore_n166;
   wire U_dfifo_U_dcore_n165;
   wire U_dfifo_U_dcore_n164;
   wire U_dfifo_U_dcore_n163;
   wire U_dfifo_U_dcore_n162;
   wire U_dfifo_U_dcore_n161;
   wire U_dfifo_U_dcore_n160;
   wire U_dfifo_U_dcore_n159;
   wire U_dfifo_U_dcore_n158;
   wire U_dfifo_U_dcore_n157;
   wire U_dfifo_U_dcore_n156;
   wire U_dfifo_U_dcore_n155;
   wire U_dfifo_U_dcore_n154;
   wire U_dfifo_U_dcore_n153;
   wire U_dfifo_U_dcore_n152;
   wire U_dfifo_U_dcore_n151;
   wire U_dfifo_U_dcore_n150;
   wire U_dfifo_U_dcore_n149;
   wire U_dfifo_U_dcore_n148;
   wire U_dfifo_U_dcore_n147;
   wire U_dfifo_U_dcore_n146;
   wire U_dfifo_U_dcore_n145;
   wire U_dfifo_U_dcore_n144;
   wire U_dfifo_U_dcore_n143;
   wire U_dfifo_U_dcore_n142;
   wire U_dfifo_U_dcore_n141;
   wire U_dfifo_U_dcore_n140;
   wire U_dfifo_U_dcore_n139;
   wire U_dfifo_U_dcore_n138;
   wire U_dfifo_U_dcore_n137;
   wire U_dfifo_U_dcore_n136;
   wire U_dfifo_U_dcore_n135;
   wire U_dfifo_U_dcore_n134;
   wire U_dfifo_U_dcore_n_empty;
   wire U_dfifo_U_dcore_f_buf_has_data;
   wire U_dfifo_U_dcore_m_sf_full;
   wire U_dfifo_U_dcore_m_sf_afull;
   wire U_dfifo_U_dcore_m_sf_empty;
   wire U_dfifo_U_dcore_f_buf_data_0_;
   wire U_dfifo_U_dcore_f_buf_data_1_;
   wire U_dfifo_U_dcore_f_buf_data_2_;
   wire U_dfifo_U_dcore_f_buf_data_3_;
   wire U_dfifo_U_dcore_f_buf_data_4_;
   wire U_dfifo_U_dcore_f_buf_data_5_;
   wire U_dfifo_U_dcore_f_buf_data_6_;
   wire U_dfifo_U_dcore_f_buf_data_7_;
   wire U_dfifo_U_dcore_f_buf_data_8_;
   wire U_dfifo_U_dcore_f_buf_data_9_;
   wire U_dfifo_U_dcore_f_buf_data_10_;
   wire U_dfifo_U_dcore_f_buf_data_11_;
   wire U_dfifo_U_dcore_f_buf_data_12_;
   wire U_dfifo_U_dcore_f_buf_data_13_;
   wire U_dfifo_U_dcore_f_buf_data_14_;
   wire U_dfifo_U_dcore_f_buf_data_15_;
   wire U_dfifo_U_dcore_f_buf_data_16_;
   wire U_dfifo_U_dcore_f_buf_data_17_;
   wire U_dfifo_U_dcore_f_buf_data_18_;
   wire U_dfifo_U_dcore_f_buf_data_19_;
   wire U_dfifo_U_dcore_f_buf_data_20_;
   wire U_dfifo_U_dcore_f_buf_data_21_;
   wire U_dfifo_U_dcore_f_buf_data_22_;
   wire U_dfifo_U_dcore_f_buf_data_23_;
   wire U_dfifo_U_dcore_f_buf_data_24_;
   wire U_dfifo_U_dcore_f_buf_data_25_;
   wire U_dfifo_U_dcore_f_buf_data_26_;
   wire U_dfifo_U_dcore_f_buf_data_27_;
   wire U_dfifo_U_dcore_f_buf_data_28_;
   wire U_dfifo_U_dcore_f_buf_data_29_;
   wire U_dfifo_U_dcore_f_buf_data_30_;
   wire U_dfifo_U_dcore_f_buf_data_31_;
   wire U_dfifo_U_dcore_f_buf_data_32_;
   wire U_dfifo_U_dcore_f_buf_data_33_;
   wire U_afifo_U_acore_U_sub_fifo_n373;
   wire U_afifo_U_acore_U_sub_fifo_n372;
   wire U_afifo_U_acore_U_sub_fifo_n371;
   wire U_afifo_U_acore_U_sub_fifo_n370;
   wire U_afifo_U_acore_U_sub_fifo_n369;
   wire U_afifo_U_acore_U_sub_fifo_n212;
   wire U_afifo_U_acore_U_sub_fifo_n169;
   wire U_afifo_U_acore_U_sub_fifo_n167;
   wire U_afifo_U_acore_U_sub_fifo_n166;
   wire U_afifo_U_acore_U_sub_fifo_n165;
   wire U_afifo_U_acore_U_sub_fifo_n163;
   wire U_afifo_U_acore_U_sub_fifo_n162;
   wire U_afifo_U_acore_U_sub_fifo_n161;
   wire U_afifo_U_acore_U_sub_fifo_n160;
   wire U_afifo_U_acore_U_sub_fifo_n159;
   wire U_afifo_U_acore_U_sub_fifo_n158;
   wire U_afifo_U_acore_U_sub_fifo_n153;
   wire U_afifo_U_acore_U_sub_fifo_n152;
   wire U_afifo_U_acore_U_sub_fifo_n151;
   wire U_afifo_U_acore_U_sub_fifo_n150;
   wire U_afifo_U_acore_U_sub_fifo_n149;
   wire U_afifo_U_acore_U_sub_fifo_n148;
   wire U_afifo_U_acore_U_sub_fifo_n147;
   wire U_afifo_U_acore_U_sub_fifo_n146;
   wire U_afifo_U_acore_U_sub_fifo_n145;
   wire U_afifo_U_acore_U_sub_fifo_n144;
   wire U_afifo_U_acore_U_sub_fifo_n143;
   wire U_afifo_U_acore_U_sub_fifo_n142;
   wire U_afifo_U_acore_U_sub_fifo_n141;
   wire U_afifo_U_acore_U_sub_fifo_n140;
   wire U_afifo_U_acore_U_sub_fifo_n139;
   wire U_afifo_U_acore_U_sub_fifo_n138;
   wire U_afifo_U_acore_U_sub_fifo_n137;
   wire U_afifo_U_acore_U_sub_fifo_n136;
   wire U_afifo_U_acore_U_sub_fifo_n135;
   wire U_afifo_U_acore_U_sub_fifo_n134;
   wire U_afifo_U_acore_U_sub_fifo_n133;
   wire U_afifo_U_acore_U_sub_fifo_n132;
   wire U_afifo_U_acore_U_sub_fifo_n131;
   wire U_afifo_U_acore_U_sub_fifo_n130;
   wire U_afifo_U_acore_U_sub_fifo_n129;
   wire U_afifo_U_acore_U_sub_fifo_n128;
   wire U_afifo_U_acore_U_sub_fifo_n127;
   wire U_afifo_U_acore_U_sub_fifo_n126;
   wire U_afifo_U_acore_U_sub_fifo_n125;
   wire U_afifo_U_acore_U_sub_fifo_n124;
   wire U_afifo_U_acore_U_sub_fifo_n123;
   wire U_afifo_U_acore_U_sub_fifo_n122;
   wire U_afifo_U_acore_U_sub_fifo_n121;
   wire U_afifo_U_acore_U_sub_fifo_n120;
   wire U_afifo_U_acore_U_sub_fifo_n119;
   wire U_afifo_U_acore_U_sub_fifo_n118;
   wire U_afifo_U_acore_U_sub_fifo_n117;
   wire U_afifo_U_acore_U_sub_fifo_n116;
   wire U_afifo_U_acore_U_sub_fifo_n115;
   wire U_afifo_U_acore_U_sub_fifo_n114;
   wire U_afifo_U_acore_U_sub_fifo_n113;
   wire U_afifo_U_acore_U_sub_fifo_n112;
   wire U_afifo_U_acore_U_sub_fifo_n111;
   wire U_afifo_U_acore_U_sub_fifo_n110;
   wire U_afifo_U_acore_U_sub_fifo_n109;
   wire U_afifo_U_acore_U_sub_fifo_n108;
   wire U_afifo_U_acore_U_sub_fifo_n107;
   wire U_afifo_U_acore_U_sub_fifo_n106;
   wire U_afifo_U_acore_U_sub_fifo_n105;
   wire U_afifo_U_acore_U_sub_fifo_n104;
   wire U_afifo_U_acore_U_sub_fifo_n103;
   wire U_afifo_U_acore_U_sub_fifo_n102;
   wire U_afifo_U_acore_U_sub_fifo_n101;
   wire U_afifo_U_acore_U_sub_fifo_n100;
   wire U_afifo_U_acore_U_sub_fifo_n99;
   wire U_afifo_U_acore_U_sub_fifo_n98;
   wire U_afifo_U_acore_U_sub_fifo_n97;
   wire U_afifo_U_acore_U_sub_fifo_n96;
   wire U_afifo_U_acore_U_sub_fifo_n95;
   wire U_afifo_U_acore_U_sub_fifo_n94;
   wire U_afifo_U_acore_U_sub_fifo_n93;
   wire U_afifo_U_acore_U_sub_fifo_n92;
   wire U_afifo_U_acore_U_sub_fifo_n91;
   wire U_afifo_U_acore_U_sub_fifo_n90;
   wire U_afifo_U_acore_U_sub_fifo_n89;
   wire U_afifo_U_acore_U_sub_fifo_n88;
   wire U_afifo_U_acore_U_sub_fifo_n87;
   wire U_afifo_U_acore_U_sub_fifo_n86;
   wire U_afifo_U_acore_U_sub_fifo_n85;
   wire U_afifo_U_acore_U_sub_fifo_n84;
   wire U_afifo_U_acore_U_sub_fifo_n83;
   wire U_afifo_U_acore_U_sub_fifo_n82;
   wire U_afifo_U_acore_U_sub_fifo_n81;
   wire U_afifo_U_acore_U_sub_fifo_n80;
   wire U_afifo_U_acore_U_sub_fifo_n79;
   wire U_afifo_U_acore_U_sub_fifo_n78;
   wire U_afifo_U_acore_U_sub_fifo_n77;
   wire U_afifo_U_acore_U_sub_fifo_n76;
   wire U_afifo_U_acore_U_sub_fifo_n75;
   wire U_afifo_U_acore_U_sub_fifo_n74;
   wire U_afifo_U_acore_U_sub_fifo_n73;
   wire U_afifo_U_acore_U_sub_fifo_n72;
   wire U_afifo_U_acore_U_sub_fifo_n71;
   wire U_afifo_U_acore_U_sub_fifo_n70;
   wire U_afifo_U_acore_U_sub_fifo_n69;
   wire U_afifo_U_acore_U_sub_fifo_n68;
   wire U_afifo_U_acore_U_sub_fifo_n67;
   wire U_afifo_U_acore_U_sub_fifo_n66;
   wire U_afifo_U_acore_U_sub_fifo_n65;
   wire U_afifo_U_acore_U_sub_fifo_n64;
   wire U_afifo_U_acore_U_sub_fifo_n63;
   wire U_afifo_U_acore_U_sub_fifo_n62;
   wire U_afifo_U_acore_U_sub_fifo_n61;
   wire U_afifo_U_acore_U_sub_fifo_n60;
   wire U_afifo_U_acore_U_sub_fifo_n59;
   wire U_afifo_U_acore_U_sub_fifo_n58;
   wire U_afifo_U_acore_U_sub_fifo_n57;
   wire U_afifo_U_acore_U_sub_fifo_n56;
   wire U_afifo_U_acore_U_sub_fifo_n55;
   wire U_afifo_U_acore_U_sub_fifo_n54;
   wire U_afifo_U_acore_U_sub_fifo_n53;
   wire U_afifo_U_acore_U_sub_fifo_n52;
   wire U_afifo_U_acore_U_sub_fifo_n51;
   wire U_afifo_U_acore_U_sub_fifo_n50;
   wire U_afifo_U_acore_U_sub_fifo_n49;
   wire U_afifo_U_acore_U_sub_fifo_n48;
   wire U_afifo_U_acore_U_sub_fifo_n47;
   wire U_afifo_U_acore_U_sub_fifo_n46;
   wire U_afifo_U_acore_U_sub_fifo_n45;
   wire U_afifo_U_acore_U_sub_fifo_n44;
   wire U_afifo_U_acore_U_sub_fifo_n43;
   wire U_afifo_U_acore_U_sub_fifo_n42;
   wire U_afifo_U_acore_U_sub_fifo_n41;
   wire U_afifo_U_acore_U_sub_fifo_n40;
   wire U_afifo_U_acore_U_sub_fifo_n39;
   wire U_afifo_U_acore_U_sub_fifo_n38;
   wire U_afifo_U_acore_U_sub_fifo_n37;
   wire U_afifo_U_acore_U_sub_fifo_n36;
   wire U_afifo_U_acore_U_sub_fifo_n35;
   wire U_afifo_U_acore_U_sub_fifo_n34;
   wire U_afifo_U_acore_U_sub_fifo_n33;
   wire U_afifo_U_acore_U_sub_fifo_n32;
   wire U_afifo_U_acore_U_sub_fifo_n31;
   wire U_afifo_U_acore_U_sub_fifo_n30;
   wire U_afifo_U_acore_U_sub_fifo_n29;
   wire U_afifo_U_acore_U_sub_fifo_n28;
   wire U_afifo_U_acore_U_sub_fifo_n27;
   wire U_afifo_U_acore_U_sub_fifo_n26;
   wire U_afifo_U_acore_U_sub_fifo_n25;
   wire U_afifo_U_acore_U_sub_fifo_n24;
   wire U_afifo_U_acore_U_sub_fifo_n23;
   wire U_afifo_U_acore_U_sub_fifo_n22;
   wire U_afifo_U_acore_U_sub_fifo_n21;
   wire U_afifo_U_acore_U_sub_fifo_n20;
   wire U_afifo_U_acore_U_sub_fifo_n19;
   wire U_afifo_U_acore_U_sub_fifo_n18;
   wire U_afifo_U_acore_U_sub_fifo_n17;
   wire U_afifo_U_acore_U_sub_fifo_n16;
   wire U_afifo_U_acore_U_sub_fifo_n15;
   wire U_afifo_U_acore_U_sub_fifo_n14;
   wire U_afifo_U_acore_U_sub_fifo_n13;
   wire U_afifo_U_acore_U_sub_fifo_n12;
   wire U_afifo_U_acore_U_sub_fifo_n11;
   wire U_afifo_U_acore_U_sub_fifo_n10;
   wire U_afifo_U_acore_U_sub_fifo_n9;
   wire U_afifo_U_acore_U_sub_fifo_n8;
   wire U_afifo_U_acore_U_sub_fifo_n7;
   wire U_afifo_U_acore_U_sub_fifo_n6;
   wire U_afifo_U_acore_U_sub_fifo_n5;
   wire U_afifo_U_acore_U_sub_fifo_n4;
   wire U_afifo_U_acore_U_sub_fifo_n3;
   wire U_afifo_U_acore_U_sub_fifo_n2;
   wire U_afifo_U_acore_U_sub_fifo_n1;
   wire U_afifo_U_acore_U_sub_fifo_n325;
   wire U_afifo_U_acore_U_sub_fifo_n324;
   wire U_afifo_U_acore_U_sub_fifo_n323;
   wire U_afifo_U_acore_U_sub_fifo_n322;
   wire U_afifo_U_acore_U_sub_fifo_n320;
   wire U_afifo_U_acore_U_sub_fifo_n319;
   wire U_afifo_U_acore_U_sub_fifo_n318;
   wire U_afifo_U_acore_U_sub_fifo_n317;
   wire U_afifo_U_acore_U_sub_fifo_n316;
   wire U_afifo_U_acore_U_sub_fifo_n315;
   wire U_afifo_U_acore_U_sub_fifo_n314;
   wire U_afifo_U_acore_U_sub_fifo_n313;
   wire U_afifo_U_acore_U_sub_fifo_n311;
   wire U_afifo_U_acore_U_sub_fifo_n310;
   wire U_afifo_U_acore_U_sub_fifo_n309;
   wire U_afifo_U_acore_U_sub_fifo_n308;
   wire U_afifo_U_acore_U_sub_fifo_n307;
   wire U_afifo_U_acore_U_sub_fifo_n306;
   wire U_afifo_U_acore_U_sub_fifo_n305;
   wire U_afifo_U_acore_U_sub_fifo_n304;
   wire U_afifo_U_acore_U_sub_fifo_n303;
   wire U_afifo_U_acore_U_sub_fifo_n302;
   wire U_afifo_U_acore_U_sub_fifo_n301;
   wire U_afifo_U_acore_U_sub_fifo_n300;
   wire U_afifo_U_acore_U_sub_fifo_n299;
   wire U_afifo_U_acore_U_sub_fifo_n298;
   wire U_afifo_U_acore_U_sub_fifo_n297;
   wire U_afifo_U_acore_U_sub_fifo_n296;
   wire U_afifo_U_acore_U_sub_fifo_n295;
   wire U_afifo_U_acore_U_sub_fifo_n294;
   wire U_afifo_U_acore_U_sub_fifo_n293;
   wire U_afifo_U_acore_U_sub_fifo_n292;
   wire U_afifo_U_acore_U_sub_fifo_n291;
   wire U_afifo_U_acore_U_sub_fifo_n290;
   wire U_afifo_U_acore_U_sub_fifo_n289;
   wire U_afifo_U_acore_U_sub_fifo_n288;
   wire U_afifo_U_acore_U_sub_fifo_n287;
   wire U_afifo_U_acore_U_sub_fifo_n286;
   wire U_afifo_U_acore_U_sub_fifo_n285;
   wire U_afifo_U_acore_U_sub_fifo_n284;
   wire U_afifo_U_acore_U_sub_fifo_n283;
   wire U_afifo_U_acore_U_sub_fifo_n282;
   wire U_afifo_U_acore_U_sub_fifo_n281;
   wire U_afifo_U_acore_U_sub_fifo_n280;
   wire U_afifo_U_acore_U_sub_fifo_n279;
   wire U_afifo_U_acore_U_sub_fifo_n278;
   wire U_afifo_U_acore_U_sub_fifo_n277;
   wire U_afifo_U_acore_U_sub_fifo_n276;
   wire U_afifo_U_acore_U_sub_fifo_n275;
   wire U_afifo_U_acore_U_sub_fifo_n274;
   wire U_afifo_U_acore_U_sub_fifo_n273;
   wire U_afifo_U_acore_U_sub_fifo_n272;
   wire U_afifo_U_acore_U_sub_fifo_n270;
   wire U_afifo_U_acore_U_sub_fifo_n269;
   wire U_afifo_U_acore_U_sub_fifo_n268;
   wire U_afifo_U_acore_U_sub_fifo_n267;
   wire U_afifo_U_acore_U_sub_fifo_n266;
   wire U_afifo_U_acore_U_sub_fifo_n265;
   wire U_afifo_U_acore_U_sub_fifo_n264;
   wire U_afifo_U_acore_U_sub_fifo_n263;
   wire U_afifo_U_acore_U_sub_fifo_n261;
   wire U_afifo_U_acore_U_sub_fifo_n260;
   wire U_afifo_U_acore_U_sub_fifo_n259;
   wire U_afifo_U_acore_U_sub_fifo_n258;
   wire U_afifo_U_acore_U_sub_fifo_n257;
   wire U_afifo_U_acore_U_sub_fifo_n256;
   wire U_afifo_U_acore_U_sub_fifo_n255;
   wire U_afifo_U_acore_U_sub_fifo_n254;
   wire U_afifo_U_acore_U_sub_fifo_n253;
   wire U_afifo_U_acore_U_sub_fifo_n252;
   wire U_afifo_U_acore_U_sub_fifo_n251;
   wire U_afifo_U_acore_U_sub_fifo_n250;
   wire U_afifo_U_acore_U_sub_fifo_n249;
   wire U_afifo_U_acore_U_sub_fifo_n248;
   wire U_afifo_U_acore_U_sub_fifo_n247;
   wire U_afifo_U_acore_U_sub_fifo_n246;
   wire U_afifo_U_acore_U_sub_fifo_n245;
   wire U_afifo_U_acore_U_sub_fifo_n244;
   wire U_afifo_U_acore_U_sub_fifo_n243;
   wire U_afifo_U_acore_U_sub_fifo_n242;
   wire U_afifo_U_acore_U_sub_fifo_n241;
   wire U_afifo_U_acore_U_sub_fifo_n240;
   wire U_afifo_U_acore_U_sub_fifo_n239;
   wire U_afifo_U_acore_U_sub_fifo_n238;
   wire U_afifo_U_acore_U_sub_fifo_n237;
   wire U_afifo_U_acore_U_sub_fifo_n236;
   wire U_afifo_U_acore_U_sub_fifo_n235;
   wire U_afifo_U_acore_U_sub_fifo_n234;
   wire U_afifo_U_acore_U_sub_fifo_n233;
   wire U_afifo_U_acore_U_sub_fifo_n232;
   wire U_afifo_U_acore_U_sub_fifo_n231;
   wire U_afifo_U_acore_U_sub_fifo_n230;
   wire U_afifo_U_acore_U_sub_fifo_n229;
   wire U_afifo_U_acore_U_sub_fifo_n228;
   wire U_afifo_U_acore_U_sub_fifo_n227;
   wire U_afifo_U_acore_U_sub_fifo_n226;
   wire U_afifo_U_acore_U_sub_fifo_n225;
   wire U_afifo_U_acore_U_sub_fifo_n224;
   wire U_afifo_U_acore_U_sub_fifo_n223;
   wire U_afifo_U_acore_U_sub_fifo_n222;
   wire U_afifo_U_acore_U_sub_fifo_n220;
   wire U_afifo_U_acore_U_sub_fifo_n219;
   wire U_afifo_U_acore_U_sub_fifo_n218;
   wire U_afifo_U_acore_U_sub_fifo_n217;
   wire U_afifo_U_acore_U_sub_fifo_n216;
   wire U_afifo_U_acore_U_sub_fifo_n215;
   wire U_afifo_U_acore_U_sub_fifo_n214;
   wire U_afifo_U_acore_U_sub_fifo_n213;
   wire U_afifo_U_acore_U_sub_fifo_n211;
   wire U_afifo_U_acore_U_sub_fifo_n210;
   wire U_afifo_U_acore_U_sub_fifo_n209;
   wire U_afifo_U_acore_U_sub_fifo_n208;
   wire U_afifo_U_acore_U_sub_fifo_n207;
   wire U_afifo_U_acore_U_sub_fifo_n206;
   wire U_afifo_U_acore_U_sub_fifo_n205;
   wire U_afifo_U_acore_U_sub_fifo_n204;
   wire U_afifo_U_acore_U_sub_fifo_n203;
   wire U_afifo_U_acore_U_sub_fifo_n202;
   wire U_afifo_U_acore_U_sub_fifo_n201;
   wire U_afifo_U_acore_U_sub_fifo_n200;
   wire U_afifo_U_acore_U_sub_fifo_n199;
   wire U_afifo_U_acore_U_sub_fifo_n198;
   wire U_afifo_U_acore_U_sub_fifo_n197;
   wire U_afifo_U_acore_U_sub_fifo_n196;
   wire U_afifo_U_acore_U_sub_fifo_n195;
   wire U_afifo_U_acore_U_sub_fifo_n194;
   wire U_afifo_U_acore_U_sub_fifo_n193;
   wire U_afifo_U_acore_U_sub_fifo_n192;
   wire U_afifo_U_acore_U_sub_fifo_n191;
   wire U_afifo_U_acore_U_sub_fifo_n190;
   wire U_afifo_U_acore_U_sub_fifo_n189;
   wire U_afifo_U_acore_U_sub_fifo_n188;
   wire U_afifo_U_acore_U_sub_fifo_n187;
   wire U_afifo_U_acore_U_sub_fifo_n186;
   wire U_afifo_U_acore_U_sub_fifo_n185;
   wire U_afifo_U_acore_U_sub_fifo_n184;
   wire U_afifo_U_acore_U_sub_fifo_n183;
   wire U_afifo_U_acore_U_sub_fifo_n182;
   wire U_afifo_U_acore_U_sub_fifo_n181;
   wire U_afifo_U_acore_U_sub_fifo_n180;
   wire U_afifo_U_acore_U_sub_fifo_n179;
   wire U_afifo_U_acore_U_sub_fifo_n178;
   wire U_afifo_U_acore_U_sub_fifo_n177;
   wire U_afifo_U_acore_U_sub_fifo_n176;
   wire U_afifo_U_acore_U_sub_fifo_n175;
   wire U_afifo_U_acore_U_sub_fifo_n174;
   wire U_afifo_U_acore_U_sub_fifo_n173;
   wire U_afifo_U_acore_U_sub_fifo_n172;
   wire U_afifo_U_acore_U_sub_fifo_n171;
   wire U_afifo_U_acore_U_sub_fifo_n170;
   wire U_afifo_U_acore_U_sub_fifo_in_ptr_1_;
   wire U_afifo_U_acore_U_sub_fifo_count_0_;
   wire U_afifo_U_acore_U_sub_fifo_count_1_;
   wire U_afifo_U_acore_U_sub_fifo_out_ptr_0_;
   wire U_afifo_U_acore_U_sub_fifo_out_ptr_1_;
   wire U_dfifo_U_dcore_U_sub_fifo_n609;
   wire U_dfifo_U_dcore_U_sub_fifo_n608;
   wire U_dfifo_U_dcore_U_sub_fifo_n607;
   wire U_dfifo_U_dcore_U_sub_fifo_n606;
   wire U_dfifo_U_dcore_U_sub_fifo_n605;
   wire U_dfifo_U_dcore_U_sub_fifo_n604;
   wire U_dfifo_U_dcore_U_sub_fifo_n603;
   wire U_dfifo_U_dcore_U_sub_fifo_n602;
   wire U_dfifo_U_dcore_U_sub_fifo_n567;
   wire U_dfifo_U_dcore_U_sub_fifo_n566;
   wire U_dfifo_U_dcore_U_sub_fifo_n565;
   wire U_dfifo_U_dcore_U_sub_fifo_n564;
   wire U_dfifo_U_dcore_U_sub_fifo_n563;
   wire U_dfifo_U_dcore_U_sub_fifo_n562;
   wire U_dfifo_U_dcore_U_sub_fifo_n561;
   wire U_dfifo_U_dcore_U_sub_fifo_n560;
   wire U_dfifo_U_dcore_U_sub_fifo_n559;
   wire U_dfifo_U_dcore_U_sub_fifo_n558;
   wire U_dfifo_U_dcore_U_sub_fifo_n557;
   wire U_dfifo_U_dcore_U_sub_fifo_n556;
   wire U_dfifo_U_dcore_U_sub_fifo_n555;
   wire U_dfifo_U_dcore_U_sub_fifo_n554;
   wire U_dfifo_U_dcore_U_sub_fifo_n553;
   wire U_dfifo_U_dcore_U_sub_fifo_n552;
   wire U_dfifo_U_dcore_U_sub_fifo_n551;
   wire U_dfifo_U_dcore_U_sub_fifo_n550;
   wire U_dfifo_U_dcore_U_sub_fifo_n549;
   wire U_dfifo_U_dcore_U_sub_fifo_n548;
   wire U_dfifo_U_dcore_U_sub_fifo_n547;
   wire U_dfifo_U_dcore_U_sub_fifo_n546;
   wire U_dfifo_U_dcore_U_sub_fifo_n545;
   wire U_dfifo_U_dcore_U_sub_fifo_n544;
   wire U_dfifo_U_dcore_U_sub_fifo_n543;
   wire U_dfifo_U_dcore_U_sub_fifo_n542;
   wire U_dfifo_U_dcore_U_sub_fifo_n541;
   wire U_dfifo_U_dcore_U_sub_fifo_n540;
   wire U_dfifo_U_dcore_U_sub_fifo_n539;
   wire U_dfifo_U_dcore_U_sub_fifo_n538;
   wire U_dfifo_U_dcore_U_sub_fifo_n537;
   wire U_dfifo_U_dcore_U_sub_fifo_n536;
   wire U_dfifo_U_dcore_U_sub_fifo_n535;
   wire U_dfifo_U_dcore_U_sub_fifo_n534;
   wire U_dfifo_U_dcore_U_sub_fifo_n533;
   wire U_dfifo_U_dcore_U_sub_fifo_n532;
   wire U_dfifo_U_dcore_U_sub_fifo_n531;
   wire U_dfifo_U_dcore_U_sub_fifo_n530;
   wire U_dfifo_U_dcore_U_sub_fifo_n529;
   wire U_dfifo_U_dcore_U_sub_fifo_n528;
   wire U_dfifo_U_dcore_U_sub_fifo_n527;
   wire U_dfifo_U_dcore_U_sub_fifo_n526;
   wire U_dfifo_U_dcore_U_sub_fifo_n525;
   wire U_dfifo_U_dcore_U_sub_fifo_n524;
   wire U_dfifo_U_dcore_U_sub_fifo_n523;
   wire U_dfifo_U_dcore_U_sub_fifo_n522;
   wire U_dfifo_U_dcore_U_sub_fifo_n521;
   wire U_dfifo_U_dcore_U_sub_fifo_n520;
   wire U_dfifo_U_dcore_U_sub_fifo_n519;
   wire U_dfifo_U_dcore_U_sub_fifo_n518;
   wire U_dfifo_U_dcore_U_sub_fifo_n517;
   wire U_dfifo_U_dcore_U_sub_fifo_n516;
   wire U_dfifo_U_dcore_U_sub_fifo_n515;
   wire U_dfifo_U_dcore_U_sub_fifo_n514;
   wire U_dfifo_U_dcore_U_sub_fifo_n513;
   wire U_dfifo_U_dcore_U_sub_fifo_n512;
   wire U_dfifo_U_dcore_U_sub_fifo_n511;
   wire U_dfifo_U_dcore_U_sub_fifo_n510;
   wire U_dfifo_U_dcore_U_sub_fifo_n509;
   wire U_dfifo_U_dcore_U_sub_fifo_n508;
   wire U_dfifo_U_dcore_U_sub_fifo_n507;
   wire U_dfifo_U_dcore_U_sub_fifo_n506;
   wire U_dfifo_U_dcore_U_sub_fifo_n505;
   wire U_dfifo_U_dcore_U_sub_fifo_n504;
   wire U_dfifo_U_dcore_U_sub_fifo_n503;
   wire U_dfifo_U_dcore_U_sub_fifo_n502;
   wire U_dfifo_U_dcore_U_sub_fifo_n501;
   wire U_dfifo_U_dcore_U_sub_fifo_n500;
   wire U_dfifo_U_dcore_U_sub_fifo_n499;
   wire U_dfifo_U_dcore_U_sub_fifo_n498;
   wire U_dfifo_U_dcore_U_sub_fifo_n497;
   wire U_dfifo_U_dcore_U_sub_fifo_n496;
   wire U_dfifo_U_dcore_U_sub_fifo_n495;
   wire U_dfifo_U_dcore_U_sub_fifo_n494;
   wire U_dfifo_U_dcore_U_sub_fifo_n493;
   wire U_dfifo_U_dcore_U_sub_fifo_n492;
   wire U_dfifo_U_dcore_U_sub_fifo_n491;
   wire U_dfifo_U_dcore_U_sub_fifo_n490;
   wire U_dfifo_U_dcore_U_sub_fifo_n489;
   wire U_dfifo_U_dcore_U_sub_fifo_n488;
   wire U_dfifo_U_dcore_U_sub_fifo_n487;
   wire U_dfifo_U_dcore_U_sub_fifo_n486;
   wire U_dfifo_U_dcore_U_sub_fifo_n485;
   wire U_dfifo_U_dcore_U_sub_fifo_n484;
   wire U_dfifo_U_dcore_U_sub_fifo_n483;
   wire U_dfifo_U_dcore_U_sub_fifo_n482;
   wire U_dfifo_U_dcore_U_sub_fifo_n481;
   wire U_dfifo_U_dcore_U_sub_fifo_n480;
   wire U_dfifo_U_dcore_U_sub_fifo_n479;
   wire U_dfifo_U_dcore_U_sub_fifo_n478;
   wire U_dfifo_U_dcore_U_sub_fifo_n477;
   wire U_dfifo_U_dcore_U_sub_fifo_n476;
   wire U_dfifo_U_dcore_U_sub_fifo_n475;
   wire U_dfifo_U_dcore_U_sub_fifo_n474;
   wire U_dfifo_U_dcore_U_sub_fifo_n473;
   wire U_dfifo_U_dcore_U_sub_fifo_n472;
   wire U_dfifo_U_dcore_U_sub_fifo_n471;
   wire U_dfifo_U_dcore_U_sub_fifo_n470;
   wire U_dfifo_U_dcore_U_sub_fifo_n469;
   wire U_dfifo_U_dcore_U_sub_fifo_n468;
   wire U_dfifo_U_dcore_U_sub_fifo_n467;
   wire U_dfifo_U_dcore_U_sub_fifo_n466;
   wire U_dfifo_U_dcore_U_sub_fifo_n465;
   wire U_dfifo_U_dcore_U_sub_fifo_n464;
   wire U_dfifo_U_dcore_U_sub_fifo_n463;
   wire U_dfifo_U_dcore_U_sub_fifo_n462;
   wire U_dfifo_U_dcore_U_sub_fifo_n461;
   wire U_dfifo_U_dcore_U_sub_fifo_n460;
   wire U_dfifo_U_dcore_U_sub_fifo_n459;
   wire U_dfifo_U_dcore_U_sub_fifo_n458;
   wire U_dfifo_U_dcore_U_sub_fifo_n456;
   wire U_dfifo_U_dcore_U_sub_fifo_n455;
   wire U_dfifo_U_dcore_U_sub_fifo_n241;
   wire U_dfifo_U_dcore_U_sub_fifo_n234;
   wire U_dfifo_U_dcore_U_sub_fifo_n233;
   wire U_dfifo_U_dcore_U_sub_fifo_n232;
   wire U_dfifo_U_dcore_U_sub_fifo_n231;
   wire U_dfifo_U_dcore_U_sub_fifo_n229;
   wire U_dfifo_U_dcore_U_sub_fifo_n228;
   wire U_dfifo_U_dcore_U_sub_fifo_n227;
   wire U_dfifo_U_dcore_U_sub_fifo_n226;
   wire U_dfifo_U_dcore_U_sub_fifo_n225;
   wire U_dfifo_U_dcore_U_sub_fifo_n224;
   wire U_dfifo_U_dcore_U_sub_fifo_n223;
   wire U_dfifo_U_dcore_U_sub_fifo_n222;
   wire U_dfifo_U_dcore_U_sub_fifo_n221;
   wire U_dfifo_U_dcore_U_sub_fifo_n220;
   wire U_dfifo_U_dcore_U_sub_fifo_n219;
   wire U_dfifo_U_dcore_U_sub_fifo_n218;
   wire U_dfifo_U_dcore_U_sub_fifo_n217;
   wire U_dfifo_U_dcore_U_sub_fifo_n216;
   wire U_dfifo_U_dcore_U_sub_fifo_n215;
   wire U_dfifo_U_dcore_U_sub_fifo_n214;
   wire U_dfifo_U_dcore_U_sub_fifo_n213;
   wire U_dfifo_U_dcore_U_sub_fifo_n212;
   wire U_dfifo_U_dcore_U_sub_fifo_n211;
   wire U_dfifo_U_dcore_U_sub_fifo_n210;
   wire U_dfifo_U_dcore_U_sub_fifo_n209;
   wire U_dfifo_U_dcore_U_sub_fifo_n208;
   wire U_dfifo_U_dcore_U_sub_fifo_n207;
   wire U_dfifo_U_dcore_U_sub_fifo_n206;
   wire U_dfifo_U_dcore_U_sub_fifo_n205;
   wire U_dfifo_U_dcore_U_sub_fifo_n204;
   wire U_dfifo_U_dcore_U_sub_fifo_n203;
   wire U_dfifo_U_dcore_U_sub_fifo_n202;
   wire U_dfifo_U_dcore_U_sub_fifo_n201;
   wire U_dfifo_U_dcore_U_sub_fifo_n200;
   wire U_dfifo_U_dcore_U_sub_fifo_n199;
   wire U_dfifo_U_dcore_U_sub_fifo_n198;
   wire U_dfifo_U_dcore_U_sub_fifo_n197;
   wire U_dfifo_U_dcore_U_sub_fifo_n196;
   wire U_dfifo_U_dcore_U_sub_fifo_n195;
   wire U_dfifo_U_dcore_U_sub_fifo_n194;
   wire U_dfifo_U_dcore_U_sub_fifo_n193;
   wire U_dfifo_U_dcore_U_sub_fifo_n192;
   wire U_dfifo_U_dcore_U_sub_fifo_n191;
   wire U_dfifo_U_dcore_U_sub_fifo_n190;
   wire U_dfifo_U_dcore_U_sub_fifo_n189;
   wire U_dfifo_U_dcore_U_sub_fifo_n188;
   wire U_dfifo_U_dcore_U_sub_fifo_n187;
   wire U_dfifo_U_dcore_U_sub_fifo_n186;
   wire U_dfifo_U_dcore_U_sub_fifo_n185;
   wire U_dfifo_U_dcore_U_sub_fifo_n184;
   wire U_dfifo_U_dcore_U_sub_fifo_n183;
   wire U_dfifo_U_dcore_U_sub_fifo_n182;
   wire U_dfifo_U_dcore_U_sub_fifo_n181;
   wire U_dfifo_U_dcore_U_sub_fifo_n180;
   wire U_dfifo_U_dcore_U_sub_fifo_n179;
   wire U_dfifo_U_dcore_U_sub_fifo_n178;
   wire U_dfifo_U_dcore_U_sub_fifo_n177;
   wire U_dfifo_U_dcore_U_sub_fifo_n176;
   wire U_dfifo_U_dcore_U_sub_fifo_n175;
   wire U_dfifo_U_dcore_U_sub_fifo_n174;
   wire U_dfifo_U_dcore_U_sub_fifo_n173;
   wire U_dfifo_U_dcore_U_sub_fifo_n172;
   wire U_dfifo_U_dcore_U_sub_fifo_n171;
   wire U_dfifo_U_dcore_U_sub_fifo_n170;
   wire U_dfifo_U_dcore_U_sub_fifo_n169;
   wire U_dfifo_U_dcore_U_sub_fifo_n168;
   wire U_dfifo_U_dcore_U_sub_fifo_n167;
   wire U_dfifo_U_dcore_U_sub_fifo_n166;
   wire U_dfifo_U_dcore_U_sub_fifo_n165;
   wire U_dfifo_U_dcore_U_sub_fifo_n164;
   wire U_dfifo_U_dcore_U_sub_fifo_n163;
   wire U_dfifo_U_dcore_U_sub_fifo_n162;
   wire U_dfifo_U_dcore_U_sub_fifo_n161;
   wire U_dfifo_U_dcore_U_sub_fifo_n160;
   wire U_dfifo_U_dcore_U_sub_fifo_n159;
   wire U_dfifo_U_dcore_U_sub_fifo_n158;
   wire U_dfifo_U_dcore_U_sub_fifo_n157;
   wire U_dfifo_U_dcore_U_sub_fifo_n156;
   wire U_dfifo_U_dcore_U_sub_fifo_n155;
   wire U_dfifo_U_dcore_U_sub_fifo_n154;
   wire U_dfifo_U_dcore_U_sub_fifo_n153;
   wire U_dfifo_U_dcore_U_sub_fifo_n152;
   wire U_dfifo_U_dcore_U_sub_fifo_n151;
   wire U_dfifo_U_dcore_U_sub_fifo_n150;
   wire U_dfifo_U_dcore_U_sub_fifo_n149;
   wire U_dfifo_U_dcore_U_sub_fifo_n148;
   wire U_dfifo_U_dcore_U_sub_fifo_n147;
   wire U_dfifo_U_dcore_U_sub_fifo_n146;
   wire U_dfifo_U_dcore_U_sub_fifo_n145;
   wire U_dfifo_U_dcore_U_sub_fifo_n144;
   wire U_dfifo_U_dcore_U_sub_fifo_n143;
   wire U_dfifo_U_dcore_U_sub_fifo_n142;
   wire U_dfifo_U_dcore_U_sub_fifo_n141;
   wire U_dfifo_U_dcore_U_sub_fifo_n140;
   wire U_dfifo_U_dcore_U_sub_fifo_n139;
   wire U_dfifo_U_dcore_U_sub_fifo_n138;
   wire U_dfifo_U_dcore_U_sub_fifo_n137;
   wire U_dfifo_U_dcore_U_sub_fifo_n136;
   wire U_dfifo_U_dcore_U_sub_fifo_n135;
   wire U_dfifo_U_dcore_U_sub_fifo_n134;
   wire U_dfifo_U_dcore_U_sub_fifo_n133;
   wire U_dfifo_U_dcore_U_sub_fifo_n132;
   wire U_dfifo_U_dcore_U_sub_fifo_n131;
   wire U_dfifo_U_dcore_U_sub_fifo_n130;
   wire U_dfifo_U_dcore_U_sub_fifo_n129;
   wire U_dfifo_U_dcore_U_sub_fifo_n128;
   wire U_dfifo_U_dcore_U_sub_fifo_n127;
   wire U_dfifo_U_dcore_U_sub_fifo_n126;
   wire U_dfifo_U_dcore_U_sub_fifo_n125;
   wire U_dfifo_U_dcore_U_sub_fifo_n124;
   wire U_dfifo_U_dcore_U_sub_fifo_n123;
   wire U_dfifo_U_dcore_U_sub_fifo_n122;
   wire U_dfifo_U_dcore_U_sub_fifo_n121;
   wire U_dfifo_U_dcore_U_sub_fifo_n120;
   wire U_dfifo_U_dcore_U_sub_fifo_n119;
   wire U_dfifo_U_dcore_U_sub_fifo_n118;
   wire U_dfifo_U_dcore_U_sub_fifo_n117;
   wire U_dfifo_U_dcore_U_sub_fifo_n116;
   wire U_dfifo_U_dcore_U_sub_fifo_n115;
   wire U_dfifo_U_dcore_U_sub_fifo_n114;
   wire U_dfifo_U_dcore_U_sub_fifo_n113;
   wire U_dfifo_U_dcore_U_sub_fifo_n112;
   wire U_dfifo_U_dcore_U_sub_fifo_n111;
   wire U_dfifo_U_dcore_U_sub_fifo_n110;
   wire U_dfifo_U_dcore_U_sub_fifo_n109;
   wire U_dfifo_U_dcore_U_sub_fifo_n108;
   wire U_dfifo_U_dcore_U_sub_fifo_n107;
   wire U_dfifo_U_dcore_U_sub_fifo_n106;
   wire U_dfifo_U_dcore_U_sub_fifo_n105;
   wire U_dfifo_U_dcore_U_sub_fifo_n104;
   wire U_dfifo_U_dcore_U_sub_fifo_n103;
   wire U_dfifo_U_dcore_U_sub_fifo_n102;
   wire U_dfifo_U_dcore_U_sub_fifo_n101;
   wire U_dfifo_U_dcore_U_sub_fifo_n100;
   wire U_dfifo_U_dcore_U_sub_fifo_n99;
   wire U_dfifo_U_dcore_U_sub_fifo_n98;
   wire U_dfifo_U_dcore_U_sub_fifo_n97;
   wire U_dfifo_U_dcore_U_sub_fifo_n96;
   wire U_dfifo_U_dcore_U_sub_fifo_n95;
   wire U_dfifo_U_dcore_U_sub_fifo_n94;
   wire U_dfifo_U_dcore_U_sub_fifo_n93;
   wire U_dfifo_U_dcore_U_sub_fifo_n92;
   wire U_dfifo_U_dcore_U_sub_fifo_n91;
   wire U_dfifo_U_dcore_U_sub_fifo_n90;
   wire U_dfifo_U_dcore_U_sub_fifo_n89;
   wire U_dfifo_U_dcore_U_sub_fifo_n88;
   wire U_dfifo_U_dcore_U_sub_fifo_n87;
   wire U_dfifo_U_dcore_U_sub_fifo_n86;
   wire U_dfifo_U_dcore_U_sub_fifo_n85;
   wire U_dfifo_U_dcore_U_sub_fifo_n84;
   wire U_dfifo_U_dcore_U_sub_fifo_n83;
   wire U_dfifo_U_dcore_U_sub_fifo_n82;
   wire U_dfifo_U_dcore_U_sub_fifo_n81;
   wire U_dfifo_U_dcore_U_sub_fifo_n80;
   wire U_dfifo_U_dcore_U_sub_fifo_n79;
   wire U_dfifo_U_dcore_U_sub_fifo_n78;
   wire U_dfifo_U_dcore_U_sub_fifo_n77;
   wire U_dfifo_U_dcore_U_sub_fifo_n76;
   wire U_dfifo_U_dcore_U_sub_fifo_n75;
   wire U_dfifo_U_dcore_U_sub_fifo_n74;
   wire U_dfifo_U_dcore_U_sub_fifo_n73;
   wire U_dfifo_U_dcore_U_sub_fifo_n72;
   wire U_dfifo_U_dcore_U_sub_fifo_n71;
   wire U_dfifo_U_dcore_U_sub_fifo_n70;
   wire U_dfifo_U_dcore_U_sub_fifo_n69;
   wire U_dfifo_U_dcore_U_sub_fifo_n68;
   wire U_dfifo_U_dcore_U_sub_fifo_n67;
   wire U_dfifo_U_dcore_U_sub_fifo_n66;
   wire U_dfifo_U_dcore_U_sub_fifo_n65;
   wire U_dfifo_U_dcore_U_sub_fifo_n64;
   wire U_dfifo_U_dcore_U_sub_fifo_n63;
   wire U_dfifo_U_dcore_U_sub_fifo_n62;
   wire U_dfifo_U_dcore_U_sub_fifo_n61;
   wire U_dfifo_U_dcore_U_sub_fifo_n60;
   wire U_dfifo_U_dcore_U_sub_fifo_n59;
   wire U_dfifo_U_dcore_U_sub_fifo_n58;
   wire U_dfifo_U_dcore_U_sub_fifo_n57;
   wire U_dfifo_U_dcore_U_sub_fifo_n56;
   wire U_dfifo_U_dcore_U_sub_fifo_n55;
   wire U_dfifo_U_dcore_U_sub_fifo_n54;
   wire U_dfifo_U_dcore_U_sub_fifo_n53;
   wire U_dfifo_U_dcore_U_sub_fifo_n52;
   wire U_dfifo_U_dcore_U_sub_fifo_n51;
   wire U_dfifo_U_dcore_U_sub_fifo_n50;
   wire U_dfifo_U_dcore_U_sub_fifo_n49;
   wire U_dfifo_U_dcore_U_sub_fifo_n48;
   wire U_dfifo_U_dcore_U_sub_fifo_n47;
   wire U_dfifo_U_dcore_U_sub_fifo_n46;
   wire U_dfifo_U_dcore_U_sub_fifo_n45;
   wire U_dfifo_U_dcore_U_sub_fifo_n44;
   wire U_dfifo_U_dcore_U_sub_fifo_n43;
   wire U_dfifo_U_dcore_U_sub_fifo_n42;
   wire U_dfifo_U_dcore_U_sub_fifo_n41;
   wire U_dfifo_U_dcore_U_sub_fifo_n40;
   wire U_dfifo_U_dcore_U_sub_fifo_n39;
   wire U_dfifo_U_dcore_U_sub_fifo_n38;
   wire U_dfifo_U_dcore_U_sub_fifo_n37;
   wire U_dfifo_U_dcore_U_sub_fifo_n36;
   wire U_dfifo_U_dcore_U_sub_fifo_n35;
   wire U_dfifo_U_dcore_U_sub_fifo_n34;
   wire U_dfifo_U_dcore_U_sub_fifo_n33;
   wire U_dfifo_U_dcore_U_sub_fifo_n32;
   wire U_dfifo_U_dcore_U_sub_fifo_n31;
   wire U_dfifo_U_dcore_U_sub_fifo_n30;
   wire U_dfifo_U_dcore_U_sub_fifo_n29;
   wire U_dfifo_U_dcore_U_sub_fifo_n28;
   wire U_dfifo_U_dcore_U_sub_fifo_n27;
   wire U_dfifo_U_dcore_U_sub_fifo_n26;
   wire U_dfifo_U_dcore_U_sub_fifo_n25;
   wire U_dfifo_U_dcore_U_sub_fifo_n24;
   wire U_dfifo_U_dcore_U_sub_fifo_n23;
   wire U_dfifo_U_dcore_U_sub_fifo_n22;
   wire U_dfifo_U_dcore_U_sub_fifo_n21;
   wire U_dfifo_U_dcore_U_sub_fifo_n20;
   wire U_dfifo_U_dcore_U_sub_fifo_n19;
   wire U_dfifo_U_dcore_U_sub_fifo_n18;
   wire U_dfifo_U_dcore_U_sub_fifo_n17;
   wire U_dfifo_U_dcore_U_sub_fifo_n16;
   wire U_dfifo_U_dcore_U_sub_fifo_n15;
   wire U_dfifo_U_dcore_U_sub_fifo_n14;
   wire U_dfifo_U_dcore_U_sub_fifo_n13;
   wire U_dfifo_U_dcore_U_sub_fifo_n12;
   wire U_dfifo_U_dcore_U_sub_fifo_n11;
   wire U_dfifo_U_dcore_U_sub_fifo_n10;
   wire U_dfifo_U_dcore_U_sub_fifo_n9;
   wire U_dfifo_U_dcore_U_sub_fifo_n8;
   wire U_dfifo_U_dcore_U_sub_fifo_n7;
   wire U_dfifo_U_dcore_U_sub_fifo_n6;
   wire U_dfifo_U_dcore_U_sub_fifo_n5;
   wire U_dfifo_U_dcore_U_sub_fifo_n4;
   wire U_dfifo_U_dcore_U_sub_fifo_n3;
   wire U_dfifo_U_dcore_U_sub_fifo_n1;
   wire U_dfifo_U_dcore_U_sub_fifo_n454;
   wire U_dfifo_U_dcore_U_sub_fifo_n453;
   wire U_dfifo_U_dcore_U_sub_fifo_n452;
   wire U_dfifo_U_dcore_U_sub_fifo_n451;
   wire U_dfifo_U_dcore_U_sub_fifo_n450;
   wire U_dfifo_U_dcore_U_sub_fifo_n449;
   wire U_dfifo_U_dcore_U_sub_fifo_n448;
   wire U_dfifo_U_dcore_U_sub_fifo_n447;
   wire U_dfifo_U_dcore_U_sub_fifo_n446;
   wire U_dfifo_U_dcore_U_sub_fifo_n445;
   wire U_dfifo_U_dcore_U_sub_fifo_n444;
   wire U_dfifo_U_dcore_U_sub_fifo_n443;
   wire U_dfifo_U_dcore_U_sub_fifo_n442;
   wire U_dfifo_U_dcore_U_sub_fifo_n441;
   wire U_dfifo_U_dcore_U_sub_fifo_n440;
   wire U_dfifo_U_dcore_U_sub_fifo_n439;
   wire U_dfifo_U_dcore_U_sub_fifo_n438;
   wire U_dfifo_U_dcore_U_sub_fifo_n437;
   wire U_dfifo_U_dcore_U_sub_fifo_n436;
   wire U_dfifo_U_dcore_U_sub_fifo_n435;
   wire U_dfifo_U_dcore_U_sub_fifo_n434;
   wire U_dfifo_U_dcore_U_sub_fifo_n433;
   wire U_dfifo_U_dcore_U_sub_fifo_n432;
   wire U_dfifo_U_dcore_U_sub_fifo_n431;
   wire U_dfifo_U_dcore_U_sub_fifo_n430;
   wire U_dfifo_U_dcore_U_sub_fifo_n429;
   wire U_dfifo_U_dcore_U_sub_fifo_n428;
   wire U_dfifo_U_dcore_U_sub_fifo_n427;
   wire U_dfifo_U_dcore_U_sub_fifo_n426;
   wire U_dfifo_U_dcore_U_sub_fifo_n425;
   wire U_dfifo_U_dcore_U_sub_fifo_n424;
   wire U_dfifo_U_dcore_U_sub_fifo_n423;
   wire U_dfifo_U_dcore_U_sub_fifo_n422;
   wire U_dfifo_U_dcore_U_sub_fifo_n421;
   wire U_dfifo_U_dcore_U_sub_fifo_n420;
   wire U_dfifo_U_dcore_U_sub_fifo_n419;
   wire U_dfifo_U_dcore_U_sub_fifo_n418;
   wire U_dfifo_U_dcore_U_sub_fifo_n417;
   wire U_dfifo_U_dcore_U_sub_fifo_n416;
   wire U_dfifo_U_dcore_U_sub_fifo_n415;
   wire U_dfifo_U_dcore_U_sub_fifo_n414;
   wire U_dfifo_U_dcore_U_sub_fifo_n413;
   wire U_dfifo_U_dcore_U_sub_fifo_n412;
   wire U_dfifo_U_dcore_U_sub_fifo_n411;
   wire U_dfifo_U_dcore_U_sub_fifo_n410;
   wire U_dfifo_U_dcore_U_sub_fifo_n409;
   wire U_dfifo_U_dcore_U_sub_fifo_n408;
   wire U_dfifo_U_dcore_U_sub_fifo_n407;
   wire U_dfifo_U_dcore_U_sub_fifo_n406;
   wire U_dfifo_U_dcore_U_sub_fifo_n405;
   wire U_dfifo_U_dcore_U_sub_fifo_n404;
   wire U_dfifo_U_dcore_U_sub_fifo_n403;
   wire U_dfifo_U_dcore_U_sub_fifo_n402;
   wire U_dfifo_U_dcore_U_sub_fifo_n401;
   wire U_dfifo_U_dcore_U_sub_fifo_n400;
   wire U_dfifo_U_dcore_U_sub_fifo_n399;
   wire U_dfifo_U_dcore_U_sub_fifo_n398;
   wire U_dfifo_U_dcore_U_sub_fifo_n397;
   wire U_dfifo_U_dcore_U_sub_fifo_n396;
   wire U_dfifo_U_dcore_U_sub_fifo_n395;
   wire U_dfifo_U_dcore_U_sub_fifo_n394;
   wire U_dfifo_U_dcore_U_sub_fifo_n393;
   wire U_dfifo_U_dcore_U_sub_fifo_n392;
   wire U_dfifo_U_dcore_U_sub_fifo_n391;
   wire U_dfifo_U_dcore_U_sub_fifo_n390;
   wire U_dfifo_U_dcore_U_sub_fifo_n389;
   wire U_dfifo_U_dcore_U_sub_fifo_n388;
   wire U_dfifo_U_dcore_U_sub_fifo_n387;
   wire U_dfifo_U_dcore_U_sub_fifo_n386;
   wire U_dfifo_U_dcore_U_sub_fifo_n385;
   wire U_dfifo_U_dcore_U_sub_fifo_n384;
   wire U_dfifo_U_dcore_U_sub_fifo_n383;
   wire U_dfifo_U_dcore_U_sub_fifo_n382;
   wire U_dfifo_U_dcore_U_sub_fifo_n381;
   wire U_dfifo_U_dcore_U_sub_fifo_n380;
   wire U_dfifo_U_dcore_U_sub_fifo_n379;
   wire U_dfifo_U_dcore_U_sub_fifo_n378;
   wire U_dfifo_U_dcore_U_sub_fifo_n377;
   wire U_dfifo_U_dcore_U_sub_fifo_n376;
   wire U_dfifo_U_dcore_U_sub_fifo_n375;
   wire U_dfifo_U_dcore_U_sub_fifo_n374;
   wire U_dfifo_U_dcore_U_sub_fifo_n373;
   wire U_dfifo_U_dcore_U_sub_fifo_n372;
   wire U_dfifo_U_dcore_U_sub_fifo_n371;
   wire U_dfifo_U_dcore_U_sub_fifo_n370;
   wire U_dfifo_U_dcore_U_sub_fifo_n369;
   wire U_dfifo_U_dcore_U_sub_fifo_n368;
   wire U_dfifo_U_dcore_U_sub_fifo_n367;
   wire U_dfifo_U_dcore_U_sub_fifo_n366;
   wire U_dfifo_U_dcore_U_sub_fifo_n365;
   wire U_dfifo_U_dcore_U_sub_fifo_n364;
   wire U_dfifo_U_dcore_U_sub_fifo_n363;
   wire U_dfifo_U_dcore_U_sub_fifo_n362;
   wire U_dfifo_U_dcore_U_sub_fifo_n361;
   wire U_dfifo_U_dcore_U_sub_fifo_n360;
   wire U_dfifo_U_dcore_U_sub_fifo_n359;
   wire U_dfifo_U_dcore_U_sub_fifo_n358;
   wire U_dfifo_U_dcore_U_sub_fifo_n357;
   wire U_dfifo_U_dcore_U_sub_fifo_n356;
   wire U_dfifo_U_dcore_U_sub_fifo_n355;
   wire U_dfifo_U_dcore_U_sub_fifo_n354;
   wire U_dfifo_U_dcore_U_sub_fifo_n353;
   wire U_dfifo_U_dcore_U_sub_fifo_n352;
   wire U_dfifo_U_dcore_U_sub_fifo_n351;
   wire U_dfifo_U_dcore_U_sub_fifo_n350;
   wire U_dfifo_U_dcore_U_sub_fifo_n349;
   wire U_dfifo_U_dcore_U_sub_fifo_n348;
   wire U_dfifo_U_dcore_U_sub_fifo_n347;
   wire U_dfifo_U_dcore_U_sub_fifo_n346;
   wire U_dfifo_U_dcore_U_sub_fifo_n345;
   wire U_dfifo_U_dcore_U_sub_fifo_n344;
   wire U_dfifo_U_dcore_U_sub_fifo_n343;
   wire U_dfifo_U_dcore_U_sub_fifo_n342;
   wire U_dfifo_U_dcore_U_sub_fifo_n341;
   wire U_dfifo_U_dcore_U_sub_fifo_n340;
   wire U_dfifo_U_dcore_U_sub_fifo_n339;
   wire U_dfifo_U_dcore_U_sub_fifo_n338;
   wire U_dfifo_U_dcore_U_sub_fifo_n337;
   wire U_dfifo_U_dcore_U_sub_fifo_n336;
   wire U_dfifo_U_dcore_U_sub_fifo_n335;
   wire U_dfifo_U_dcore_U_sub_fifo_n334;
   wire U_dfifo_U_dcore_U_sub_fifo_n333;
   wire U_dfifo_U_dcore_U_sub_fifo_n332;
   wire U_dfifo_U_dcore_U_sub_fifo_n331;
   wire U_dfifo_U_dcore_U_sub_fifo_n330;
   wire U_dfifo_U_dcore_U_sub_fifo_n329;
   wire U_dfifo_U_dcore_U_sub_fifo_n328;
   wire U_dfifo_U_dcore_U_sub_fifo_n327;
   wire U_dfifo_U_dcore_U_sub_fifo_n326;
   wire U_dfifo_U_dcore_U_sub_fifo_n325;
   wire U_dfifo_U_dcore_U_sub_fifo_n324;
   wire U_dfifo_U_dcore_U_sub_fifo_n323;
   wire U_dfifo_U_dcore_U_sub_fifo_n322;
   wire U_dfifo_U_dcore_U_sub_fifo_n321;
   wire U_dfifo_U_dcore_U_sub_fifo_n320;
   wire U_dfifo_U_dcore_U_sub_fifo_n319;
   wire U_dfifo_U_dcore_U_sub_fifo_n318;
   wire U_dfifo_U_dcore_U_sub_fifo_n317;
   wire U_dfifo_U_dcore_U_sub_fifo_n316;
   wire U_dfifo_U_dcore_U_sub_fifo_n315;
   wire U_dfifo_U_dcore_U_sub_fifo_n314;
   wire U_dfifo_U_dcore_U_sub_fifo_n313;
   wire U_dfifo_U_dcore_U_sub_fifo_n312;
   wire U_dfifo_U_dcore_U_sub_fifo_n311;
   wire U_dfifo_U_dcore_U_sub_fifo_n310;
   wire U_dfifo_U_dcore_U_sub_fifo_n309;
   wire U_dfifo_U_dcore_U_sub_fifo_n308;
   wire U_dfifo_U_dcore_U_sub_fifo_n307;
   wire U_dfifo_U_dcore_U_sub_fifo_n306;
   wire U_dfifo_U_dcore_U_sub_fifo_n305;
   wire U_dfifo_U_dcore_U_sub_fifo_n304;
   wire U_dfifo_U_dcore_U_sub_fifo_n303;
   wire U_dfifo_U_dcore_U_sub_fifo_n302;
   wire U_dfifo_U_dcore_U_sub_fifo_n301;
   wire U_dfifo_U_dcore_U_sub_fifo_n300;
   wire U_dfifo_U_dcore_U_sub_fifo_n299;
   wire U_dfifo_U_dcore_U_sub_fifo_n298;
   wire U_dfifo_U_dcore_U_sub_fifo_n297;
   wire U_dfifo_U_dcore_U_sub_fifo_n296;
   wire U_dfifo_U_dcore_U_sub_fifo_n295;
   wire U_dfifo_U_dcore_U_sub_fifo_n294;
   wire U_dfifo_U_dcore_U_sub_fifo_n293;
   wire U_dfifo_U_dcore_U_sub_fifo_n292;
   wire U_dfifo_U_dcore_U_sub_fifo_n291;
   wire U_dfifo_U_dcore_U_sub_fifo_n290;
   wire U_dfifo_U_dcore_U_sub_fifo_n289;
   wire U_dfifo_U_dcore_U_sub_fifo_n288;
   wire U_dfifo_U_dcore_U_sub_fifo_n287;
   wire U_dfifo_U_dcore_U_sub_fifo_n286;
   wire U_dfifo_U_dcore_U_sub_fifo_n285;
   wire U_dfifo_U_dcore_U_sub_fifo_n284;
   wire U_dfifo_U_dcore_U_sub_fifo_n283;
   wire U_dfifo_U_dcore_U_sub_fifo_n282;
   wire U_dfifo_U_dcore_U_sub_fifo_n281;
   wire U_dfifo_U_dcore_U_sub_fifo_n280;
   wire U_dfifo_U_dcore_U_sub_fifo_n279;
   wire U_dfifo_U_dcore_U_sub_fifo_n278;
   wire U_dfifo_U_dcore_U_sub_fifo_n277;
   wire U_dfifo_U_dcore_U_sub_fifo_n276;
   wire U_dfifo_U_dcore_U_sub_fifo_n275;
   wire U_dfifo_U_dcore_U_sub_fifo_n274;
   wire U_dfifo_U_dcore_U_sub_fifo_n273;
   wire U_dfifo_U_dcore_U_sub_fifo_n272;
   wire U_dfifo_U_dcore_U_sub_fifo_n271;
   wire U_dfifo_U_dcore_U_sub_fifo_n270;
   wire U_dfifo_U_dcore_U_sub_fifo_n269;
   wire U_dfifo_U_dcore_U_sub_fifo_n268;
   wire U_dfifo_U_dcore_U_sub_fifo_n267;
   wire U_dfifo_U_dcore_U_sub_fifo_n266;
   wire U_dfifo_U_dcore_U_sub_fifo_n265;
   wire U_dfifo_U_dcore_U_sub_fifo_n264;
   wire U_dfifo_U_dcore_U_sub_fifo_n263;
   wire U_dfifo_U_dcore_U_sub_fifo_n262;
   wire U_dfifo_U_dcore_U_sub_fifo_n261;
   wire U_dfifo_U_dcore_U_sub_fifo_n260;
   wire U_dfifo_U_dcore_U_sub_fifo_n259;
   wire U_dfifo_U_dcore_U_sub_fifo_n258;
   wire U_dfifo_U_dcore_U_sub_fifo_n257;
   wire U_dfifo_U_dcore_U_sub_fifo_n256;
   wire U_dfifo_U_dcore_U_sub_fifo_n255;
   wire U_dfifo_U_dcore_U_sub_fifo_n254;
   wire U_dfifo_U_dcore_U_sub_fifo_n253;
   wire U_dfifo_U_dcore_U_sub_fifo_n252;
   wire U_dfifo_U_dcore_U_sub_fifo_n251;
   wire U_dfifo_U_dcore_U_sub_fifo_n250;
   wire U_dfifo_U_dcore_U_sub_fifo_n249;
   wire U_dfifo_U_dcore_U_sub_fifo_n248;
   wire U_dfifo_U_dcore_U_sub_fifo_n247;
   wire U_dfifo_U_dcore_U_sub_fifo_n246;
   wire U_dfifo_U_dcore_U_sub_fifo_n245;
   wire U_dfifo_U_dcore_U_sub_fifo_n244;
   wire U_dfifo_U_dcore_U_sub_fifo_n243;
   wire U_dfifo_U_dcore_U_sub_fifo_n242;
   wire U_dfifo_U_dcore_U_sub_fifo_in_ptr_0_;
   wire U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_;
   wire U_dfifo_U_dcore_U_sub_fifo_in_ptr_2_;
   wire U_dfifo_U_dcore_U_sub_fifo_count_0_;
   wire U_dfifo_U_dcore_U_sub_fifo_count_1_;
   wire U_dfifo_U_dcore_U_sub_fifo_count_2_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__0_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__1_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__2_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__3_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__4_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__5_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__6_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__7_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__8_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__9_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__10_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__11_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__12_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__13_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__14_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__15_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__16_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__17_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__18_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__19_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__20_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__21_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__22_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__23_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__24_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__25_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__26_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__27_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__28_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__29_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__30_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__31_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__32_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_0__33_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__0_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__1_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__2_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__3_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__4_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__5_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__6_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__7_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__8_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__9_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__10_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__11_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__12_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__13_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__14_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__15_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__16_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__17_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__18_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__19_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__20_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__21_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__22_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__23_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__24_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__25_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__26_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__27_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__28_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__29_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__30_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__31_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__32_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_2__33_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__0_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__1_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__2_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__3_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__4_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__5_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__6_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__7_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__8_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__9_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__10_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__11_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__12_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__13_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__14_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__15_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__16_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__17_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__18_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__19_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__20_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__21_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__22_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__23_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__24_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__25_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__26_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__27_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__28_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__29_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__30_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__31_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__32_;
   wire U_dfifo_U_dcore_U_sub_fifo_mem_3__33_;
   wire U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_;
   wire U_dfifo_U_dcore_U_sub_fifo_out_ptr_1_;
   wire U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n48;
   wire n50;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire [16:4] m_af_data2_in;
   wire [33:0] m_df_data_in;
   wire [49:0] U_afifo_m_data_in;
   wire [15:0] U_dfifo_m_btm_data;
   wire [2:0] U_ctl_n_bh_state;
   wire [3:0] U_ctl_f_amba_bsz2;
   wire [3:0] U_ctl_f_col_width;
   wire [49:0] U_afifo_U_acore_m_sf_data_out;
   wire [33:0] U_dfifo_U_dcore_m_sf_data_out;

   CLKBUF_X1 FE_PHC5241_U_rbuf_n175 (.Z(FE_PHN5241_U_rbuf_n175), 
	.A(FE_PHN5189_U_rbuf_n175));
   CLKBUF_X1 FE_PHC5240_U_rbuf_n69 (.Z(FE_PHN5240_U_rbuf_n69), 
	.A(FE_PHN5190_U_rbuf_n69));
   CLKBUF_X1 FE_PHC5239_U_ctl_n299 (.Z(FE_PHN5239_U_ctl_n299), 
	.A(FE_PHN5203_U_ctl_n299));
   BUF_X32 FE_PHC5218_U_ctl_N89 (.Z(FE_PHN5218_U_ctl_N89), 
	.A(U_ctl_N89));
   BUF_X8 FE_PHC5203_U_ctl_n299 (.Z(FE_PHN5203_U_ctl_n299), 
	.A(U_ctl_n299));
   CLKBUF_X1 FE_PHC5191_miu_data_27_ (.Z(FE_PHN5191_miu_data_27_), 
	.A(miu_data[27]));
   CLKBUF_X1 FE_PHC5190_U_rbuf_n69 (.Z(FE_PHN5190_U_rbuf_n69), 
	.A(U_rbuf_n69));
   BUF_X8 FE_PHC5189_U_rbuf_n175 (.Z(FE_PHN5189_U_rbuf_n175), 
	.A(U_rbuf_n175));
   CLKBUF_X1 FE_PHC5181_hsel_reg (.Z(FE_PHN5181_hsel_reg), 
	.A(FE_PHN4636_hsel_reg));
   CLKBUF_X1 FE_PHC5180_U_rbuf_n63 (.Z(FE_PHN5180_U_rbuf_n63), 
	.A(FE_PHN4650_U_rbuf_n63));
   CLKBUF_X1 FE_PHC5179_U_rbuf_n72 (.Z(FE_PHN5179_U_rbuf_n72), 
	.A(U_rbuf_n72));
   CLKBUF_X1 FE_PHC5175_U_rbuf_n188 (.Z(FE_PHN5175_U_rbuf_n188), 
	.A(U_rbuf_n188));
   CLKBUF_X1 FE_PHC5165_U_afifo_U_acore_U_sub_fifo_n282 (.Z(FE_PHN5165_U_afifo_U_acore_U_sub_fifo_n282), 
	.A(FE_PHN3946_U_afifo_U_acore_U_sub_fifo_n282));
   CLKBUF_X1 FE_PHC5164_U_afifo_U_acore_U_sub_fifo_n260 (.Z(FE_PHN5164_U_afifo_U_acore_U_sub_fifo_n260), 
	.A(FE_PHN3920_U_afifo_U_acore_U_sub_fifo_n260));
   CLKBUF_X1 FE_PHC5162_U_afifo_U_acore_U_sub_fifo_n316 (.Z(FE_PHN5162_U_afifo_U_acore_U_sub_fifo_n316), 
	.A(FE_PHN3176_U_afifo_U_acore_U_sub_fifo_n316));
   CLKBUF_X1 FE_PHC5159_U_dfifo_U_dcore_U_sub_fifo_n275 (.Z(FE_PHN5159_U_dfifo_U_dcore_U_sub_fifo_n275), 
	.A(FE_PHN4157_U_dfifo_U_dcore_U_sub_fifo_n275));
   CLKBUF_X1 FE_PHC5157_U_dfifo_U_dcore_U_sub_fifo_n299 (.Z(FE_PHN5157_U_dfifo_U_dcore_U_sub_fifo_n299), 
	.A(FE_PHN4244_U_dfifo_U_dcore_U_sub_fifo_n299));
   CLKBUF_X1 FE_PHC5154_U_afifo_U_acore_U_sub_fifo_n249 (.Z(FE_PHN5154_U_afifo_U_acore_U_sub_fifo_n249), 
	.A(FE_PHN3294_U_afifo_U_acore_U_sub_fifo_n249));
   CLKBUF_X1 FE_PHC5153_U_afifo_U_acore_U_sub_fifo_n209 (.Z(FE_PHN5153_U_afifo_U_acore_U_sub_fifo_n209), 
	.A(FE_PHN3939_U_afifo_U_acore_U_sub_fifo_n209));
   CLKBUF_X2 FE_PHC5152_U_afifo_U_acore_U_sub_fifo_n294 (.Z(FE_PHN5152_U_afifo_U_acore_U_sub_fifo_n294), 
	.A(FE_PHN3174_U_afifo_U_acore_U_sub_fifo_n294));
   BUF_X1 FE_PHC5148_U_dfifo_U_dcore_U_sub_fifo_n257 (.Z(FE_PHN5148_U_dfifo_U_dcore_U_sub_fifo_n257), 
	.A(FE_PHN4236_U_dfifo_U_dcore_U_sub_fifo_n257));
   CLKBUF_X2 FE_PHC5147_U_dfifo_U_dcore_U_sub_fifo_n259 (.Z(FE_PHN5147_U_dfifo_U_dcore_U_sub_fifo_n259), 
	.A(FE_PHN4255_U_dfifo_U_dcore_U_sub_fifo_n259));
   CLKBUF_X1 FE_PHC5143_U_afifo_U_acore_U_sub_fifo_n188 (.Z(FE_PHN5143_U_afifo_U_acore_U_sub_fifo_n188), 
	.A(FE_PHN4128_U_afifo_U_acore_U_sub_fifo_n188));
   CLKBUF_X1 FE_PHC5140_U_afifo_U_acore_U_sub_fifo_n245 (.Z(FE_PHN5140_U_afifo_U_acore_U_sub_fifo_n245), 
	.A(FE_PHN3967_U_afifo_U_acore_U_sub_fifo_n245));
   CLKBUF_X1 FE_PHC5138_U_dfifo_U_dcore_U_sub_fifo_n307 (.Z(FE_PHN5138_U_dfifo_U_dcore_U_sub_fifo_n307), 
	.A(FE_PHN4194_U_dfifo_U_dcore_U_sub_fifo_n307));
   CLKBUF_X1 FE_PHC5133_U_afifo_U_acore_U_sub_fifo_n236 (.Z(FE_PHN5133_U_afifo_U_acore_U_sub_fifo_n236), 
	.A(FE_PHN3901_U_afifo_U_acore_U_sub_fifo_n236));
   CLKBUF_X1 FE_PHC5132_U_afifo_n158 (.Z(FE_PHN5132_U_afifo_n158), 
	.A(FE_PHN3897_U_afifo_n158));
   CLKBUF_X2 FE_PHC5128_U_dfifo_U_dcore_U_sub_fifo_n251 (.Z(FE_PHN5128_U_dfifo_U_dcore_U_sub_fifo_n251), 
	.A(FE_PHN4173_U_dfifo_U_dcore_U_sub_fifo_n251));
   CLKBUF_X1 FE_PHC5118_U_afifo_U_acore_U_sub_fifo_n250 (.Z(FE_PHN5118_U_afifo_U_acore_U_sub_fifo_n250), 
	.A(FE_PHN3498_U_afifo_U_acore_U_sub_fifo_n250));
   CLKBUF_X1 FE_PHC5117_U_afifo_U_acore_U_sub_fifo_n275 (.Z(FE_PHN5117_U_afifo_U_acore_U_sub_fifo_n275), 
	.A(FE_PHN4164_U_afifo_U_acore_U_sub_fifo_n275));
   CLKBUF_X1 FE_PHC5116_U_dfifo_U_dcore_U_sub_fifo_n247 (.Z(FE_PHN5116_U_dfifo_U_dcore_U_sub_fifo_n247), 
	.A(FE_PHN4184_U_dfifo_U_dcore_U_sub_fifo_n247));
   CLKBUF_X1 FE_PHC5115_U_dfifo_U_dcore_U_sub_fifo_n292 (.Z(FE_PHN5115_U_dfifo_U_dcore_U_sub_fifo_n292), 
	.A(FE_PHN4211_U_dfifo_U_dcore_U_sub_fifo_n292));
   CLKBUF_X1 FE_PHC5111_U_afifo_U_acore_U_sub_fifo_n220 (.Z(FE_PHN5111_U_afifo_U_acore_U_sub_fifo_n220), 
	.A(FE_PHN3935_U_afifo_U_acore_U_sub_fifo_n220));
   BUF_X1 FE_PHC5109_U_dfifo_U_dcore_U_sub_fifo_n310 (.Z(FE_PHN5109_U_dfifo_U_dcore_U_sub_fifo_n310), 
	.A(FE_PHN4225_U_dfifo_U_dcore_U_sub_fifo_n310));
   CLKBUF_X1 FE_PHC5103_U_afifo_U_acore_U_sub_fifo_n308 (.Z(FE_PHN5103_U_afifo_U_acore_U_sub_fifo_n308), 
	.A(FE_PHN3171_U_afifo_U_acore_U_sub_fifo_n308));
   CLKBUF_X1 FE_PHC5101_U_afifo_U_acore_U_sub_fifo_n177 (.Z(FE_PHN5101_U_afifo_U_acore_U_sub_fifo_n177), 
	.A(FE_PHN3491_U_afifo_U_acore_U_sub_fifo_n177));
   CLKBUF_X1 FE_PHC5100_U_afifo_n159 (.Z(FE_PHN5100_U_afifo_n159), 
	.A(FE_PHN4186_U_afifo_n159));
   CLKBUF_X1 FE_PHC5098_U_afifo_U_acore_U_sub_fifo_n251 (.Z(FE_PHN5098_U_afifo_U_acore_U_sub_fifo_n251), 
	.A(FE_PHN3484_U_afifo_U_acore_U_sub_fifo_n251));
   CLKBUF_X1 FE_PHC5095_U_afifo_U_acore_U_sub_fifo_n194 (.Z(FE_PHN5095_U_afifo_U_acore_U_sub_fifo_n194), 
	.A(FE_PHN3947_U_afifo_U_acore_U_sub_fifo_n194));
   CLKBUF_X1 FE_PHC5092_U_dfifo_U_dcore_U_sub_fifo_n287 (.Z(FE_PHN5092_U_dfifo_U_dcore_U_sub_fifo_n287), 
	.A(FE_PHN4095_U_dfifo_U_dcore_U_sub_fifo_n287));
   CLKBUF_X2 FE_PHC5087_U_afifo_U_acore_U_sub_fifo_n265 (.Z(FE_PHN5087_U_afifo_U_acore_U_sub_fifo_n265), 
	.A(FE_PHN4121_U_afifo_U_acore_U_sub_fifo_n265));
   BUF_X1 FE_PHC5083_U_dfifo_U_dcore_U_sub_fifo_n274 (.Z(FE_PHN5083_U_dfifo_U_dcore_U_sub_fifo_n274), 
	.A(FE_PHN4222_U_dfifo_U_dcore_U_sub_fifo_n274));
   BUF_X1 FE_PHC5082_U_dfifo_U_dcore_U_sub_fifo_n280 (.Z(FE_PHN5082_U_dfifo_U_dcore_U_sub_fifo_n280), 
	.A(FE_PHN4188_U_dfifo_U_dcore_U_sub_fifo_n280));
   CLKBUF_X2 FE_PHC5081_U_afifo_U_acore_U_sub_fifo_n309 (.Z(FE_PHN5081_U_afifo_U_acore_U_sub_fifo_n309), 
	.A(FE_PHN4223_U_afifo_U_acore_U_sub_fifo_n309));
   BUF_X1 FE_PHC5079_U_afifo_U_acore_U_sub_fifo_n231 (.Z(FE_PHN5079_U_afifo_U_acore_U_sub_fifo_n231), 
	.A(FE_PHN3936_U_afifo_U_acore_U_sub_fifo_n231));
   BUF_X1 FE_PHC5078_U_afifo_U_acore_U_sub_fifo_n246 (.Z(FE_PHN5078_U_afifo_U_acore_U_sub_fifo_n246), 
	.A(FE_PHN3881_U_afifo_U_acore_U_sub_fifo_n246));
   CLKBUF_X1 FE_PHC5075_U_afifo_U_acore_U_sub_fifo_n213 (.Z(FE_PHN5075_U_afifo_U_acore_U_sub_fifo_n213), 
	.A(FE_PHN4081_U_afifo_U_acore_U_sub_fifo_n213));
   CLKBUF_X1 FE_PHC5073_U_afifo_U_acore_U_sub_fifo_n180 (.Z(FE_PHN5073_U_afifo_U_acore_U_sub_fifo_n180), 
	.A(FE_PHN4111_U_afifo_U_acore_U_sub_fifo_n180));
   CLKBUF_X1 FE_PHC5072_U_dfifo_U_dcore_U_sub_fifo_n263 (.Z(FE_PHN5072_U_dfifo_U_dcore_U_sub_fifo_n263), 
	.A(FE_PHN4125_U_dfifo_U_dcore_U_sub_fifo_n263));
   CLKBUF_X1 FE_PHC5071_U_afifo_U_acore_U_sub_fifo_n264 (.Z(FE_PHN5071_U_afifo_U_acore_U_sub_fifo_n264), 
	.A(FE_PHN4099_U_afifo_U_acore_U_sub_fifo_n264));
   CLKBUF_X1 FE_PHC5070_U_dfifo_U_dcore_U_sub_fifo_n308 (.Z(FE_PHN5070_U_dfifo_U_dcore_U_sub_fifo_n308), 
	.A(FE_PHN4195_U_dfifo_U_dcore_U_sub_fifo_n308));
   CLKBUF_X1 FE_PHC5069_U_afifo_U_acore_U_sub_fifo_n185 (.Z(FE_PHN5069_U_afifo_U_acore_U_sub_fifo_n185), 
	.A(FE_PHN3891_U_afifo_U_acore_U_sub_fifo_n185));
   CLKBUF_X1 FE_PHC5068_U_afifo_U_acore_U_sub_fifo_n243 (.Z(FE_PHN5068_U_afifo_U_acore_U_sub_fifo_n243), 
	.A(FE_PHN3483_U_afifo_U_acore_U_sub_fifo_n243));
   CLKBUF_X1 FE_PHC5067_U_afifo_U_acore_U_sub_fifo_n307 (.Z(FE_PHN5067_U_afifo_U_acore_U_sub_fifo_n307), 
	.A(FE_PHN3157_U_afifo_U_acore_U_sub_fifo_n307));
   CLKBUF_X1 FE_PHC5063_U_afifo_U_acore_U_sub_fifo_n227 (.Z(FE_PHN5063_U_afifo_U_acore_U_sub_fifo_n227), 
	.A(FE_PHN3490_U_afifo_U_acore_U_sub_fifo_n227));
   CLKBUF_X1 FE_PHC5062_U_dfifo_U_dcore_U_sub_fifo_n297 (.Z(FE_PHN5062_U_dfifo_U_dcore_U_sub_fifo_n297), 
	.A(FE_PHN4073_U_dfifo_U_dcore_U_sub_fifo_n297));
   CLKBUF_X1 FE_PHC5058_U_afifo_U_acore_U_sub_fifo_n205 (.Z(FE_PHN5058_U_afifo_U_acore_U_sub_fifo_n205), 
	.A(FE_PHN4163_U_afifo_U_acore_U_sub_fifo_n205));
   CLKBUF_X1 FE_PHC5057_U_dfifo_U_dcore_U_sub_fifo_n285 (.Z(FE_PHN5057_U_dfifo_U_dcore_U_sub_fifo_n285), 
	.A(FE_PHN4190_U_dfifo_U_dcore_U_sub_fifo_n285));
   CLKBUF_X2 FE_PHC5054_U_dfifo_U_dcore_n153 (.Z(FE_PHN5054_U_dfifo_U_dcore_n153), 
	.A(FE_PHN4155_U_dfifo_U_dcore_n153));
   CLKBUF_X2 FE_PHC5051_U_dfifo_U_dcore_U_sub_fifo_n254 (.Z(FE_PHN5051_U_dfifo_U_dcore_U_sub_fifo_n254), 
	.A(FE_PHN4228_U_dfifo_U_dcore_U_sub_fifo_n254));
   BUF_X1 FE_PHC5048_U_afifo_U_acore_U_sub_fifo_n255 (.Z(FE_PHN5048_U_afifo_U_acore_U_sub_fifo_n255), 
	.A(FE_PHN3890_U_afifo_U_acore_U_sub_fifo_n255));
   CLKBUF_X1 FE_PHC5041_U_dfifo_U_dcore_U_sub_fifo_n178 (.Z(FE_PHN5041_U_dfifo_U_dcore_U_sub_fifo_n178), 
	.A(FE_PHN3850_U_dfifo_U_dcore_U_sub_fifo_n178));
   CLKBUF_X1 FE_PHC5040_U_afifo_U_acore_U_sub_fifo_n237 (.Z(FE_PHN5040_U_afifo_U_acore_U_sub_fifo_n237), 
	.A(FE_PHN3905_U_afifo_U_acore_U_sub_fifo_n237));
   CLKBUF_X1 FE_PHC5038_U_afifo_U_acore_U_sub_fifo_n274 (.Z(FE_PHN5038_U_afifo_U_acore_U_sub_fifo_n274), 
	.A(FE_PHN3172_U_afifo_U_acore_U_sub_fifo_n274));
   CLKBUF_X1 FE_PHC5037_U_afifo_U_acore_U_sub_fifo_n315 (.Z(FE_PHN5037_U_afifo_U_acore_U_sub_fifo_n315), 
	.A(FE_PHN4069_U_afifo_U_acore_U_sub_fifo_n315));
   CLKBUF_X1 FE_PHC5036_U_dfifo_U_dcore_U_sub_fifo_n255 (.Z(FE_PHN5036_U_dfifo_U_dcore_U_sub_fifo_n255), 
	.A(FE_PHN4210_U_dfifo_U_dcore_U_sub_fifo_n255));
   CLKBUF_X1 FE_PHC5033_U_dfifo_U_dcore_U_sub_fifo_n281 (.Z(FE_PHN5033_U_dfifo_U_dcore_U_sub_fifo_n281), 
	.A(FE_PHN4130_U_dfifo_U_dcore_U_sub_fifo_n281));
   CLKBUF_X1 FE_PHC5032_U_afifo_U_acore_U_sub_fifo_n192 (.Z(FE_PHN5032_U_afifo_U_acore_U_sub_fifo_n192), 
	.A(FE_PHN4179_U_afifo_U_acore_U_sub_fifo_n192));
   CLKBUF_X1 FE_PHC5030_U_dfifo_U_dcore_U_sub_fifo_n304 (.Z(FE_PHN5030_U_dfifo_U_dcore_U_sub_fifo_n304), 
	.A(FE_PHN4151_U_dfifo_U_dcore_U_sub_fifo_n304));
   BUF_X1 FE_PHC5024_U_afifo_n17 (.Z(FE_PHN5024_U_afifo_n17), 
	.A(FE_PHN4105_U_afifo_n17));
   BUF_X1 FE_PHC5022_U_afifo_U_acore_U_sub_fifo_n191 (.Z(FE_PHN5022_U_afifo_U_acore_U_sub_fifo_n191), 
	.A(FE_PHN4158_U_afifo_U_acore_U_sub_fifo_n191));
   CLKBUF_X2 FE_PHC5021_U_afifo_n166 (.Z(FE_PHN5021_U_afifo_n166), 
	.A(FE_PHN4079_U_afifo_n166));
   CLKBUF_X1 FE_PHC5020_U_afifo_U_acore_U_sub_fifo_n184 (.Z(FE_PHN5020_U_afifo_U_acore_U_sub_fifo_n184), 
	.A(FE_PHN4153_U_afifo_U_acore_U_sub_fifo_n184));
   BUF_X1 FE_PHC5016_U_dfifo_U_dcore_n156 (.Z(FE_PHN5016_U_dfifo_U_dcore_n156), 
	.A(FE_PHN4207_U_dfifo_U_dcore_n156));
   CLKBUF_X1 FE_PHC5009_U_afifo_U_acore_U_sub_fifo_n273 (.Z(FE_PHN5009_U_afifo_U_acore_U_sub_fifo_n273), 
	.A(FE_PHN3308_U_afifo_U_acore_U_sub_fifo_n273));
   CLKBUF_X1 FE_PHC5007_U_afifo_U_acore_U_sub_fifo_n285 (.Z(FE_PHN5007_U_afifo_U_acore_U_sub_fifo_n285), 
	.A(FE_PHN4106_U_afifo_U_acore_U_sub_fifo_n285));
   CLKBUF_X1 FE_PHC5005_U_afifo_U_acore_U_sub_fifo_n187 (.Z(FE_PHN5005_U_afifo_U_acore_U_sub_fifo_n187), 
	.A(FE_PHN4159_U_afifo_U_acore_U_sub_fifo_n187));
   CLKBUF_X1 FE_PHC5004_U_afifo_n165 (.Z(FE_PHN5004_U_afifo_n165), 
	.A(FE_PHN4025_U_afifo_n165));
   CLKBUF_X1 FE_PHC5003_U_afifo_U_acore_U_sub_fifo_n283 (.Z(FE_PHN5003_U_afifo_U_acore_U_sub_fifo_n283), 
	.A(FE_PHN4098_U_afifo_U_acore_U_sub_fifo_n283));
   BUF_X1 FE_PHC4998_U_dfifo_U_dcore_U_sub_fifo_n302 (.Z(FE_PHN4998_U_dfifo_U_dcore_U_sub_fifo_n302), 
	.A(FE_PHN4033_U_dfifo_U_dcore_U_sub_fifo_n302));
   CLKBUF_X2 FE_PHC4996_U_afifo_U_acore_U_sub_fifo_n202 (.Z(FE_PHN4996_U_afifo_U_acore_U_sub_fifo_n202), 
	.A(FE_PHN3307_U_afifo_U_acore_U_sub_fifo_n202));
   BUF_X1 FE_PHC4993_U_dfifo_U_dcore_U_sub_fifo_n279 (.Z(FE_PHN4993_U_dfifo_U_dcore_U_sub_fifo_n279), 
	.A(FE_PHN4143_U_dfifo_U_dcore_U_sub_fifo_n279));
   BUF_X1 FE_PHC4992_U_afifo_U_acore_U_sub_fifo_n235 (.Z(FE_PHN4992_U_afifo_U_acore_U_sub_fifo_n235), 
	.A(FE_PHN3895_U_afifo_U_acore_U_sub_fifo_n235));
   CLKBUF_X1 FE_PHC4987_U_afifo_U_acore_U_sub_fifo_n210 (.Z(FE_PHN4987_U_afifo_U_acore_U_sub_fifo_n210), 
	.A(FE_PHN4134_U_afifo_U_acore_U_sub_fifo_n210));
   CLKBUF_X1 FE_PHC4981_U_afifo_U_acore_U_sub_fifo_n277 (.Z(FE_PHN4981_U_afifo_U_acore_U_sub_fifo_n277), 
	.A(FE_PHN3304_U_afifo_U_acore_U_sub_fifo_n277));
   CLKBUF_X1 FE_PHC4979_U_afifo_U_acore_U_sub_fifo_n173 (.Z(FE_PHN4979_U_afifo_U_acore_U_sub_fifo_n173), 
	.A(FE_PHN3495_U_afifo_U_acore_U_sub_fifo_n173));
   CLKBUF_X1 FE_PHC4978_U_afifo_U_acore_U_sub_fifo_n247 (.Z(FE_PHN4978_U_afifo_U_acore_U_sub_fifo_n247), 
	.A(FE_PHN4049_U_afifo_U_acore_U_sub_fifo_n247));
   CLKBUF_X1 FE_PHC4975_U_dfifo_U_dcore_U_sub_fifo_n213 (.Z(FE_PHN4975_U_dfifo_U_dcore_U_sub_fifo_n213), 
	.A(FE_PHN3899_U_dfifo_U_dcore_U_sub_fifo_n213));
   BUF_X1 FE_PHC4973_U_afifo_U_acore_U_sub_fifo_n218 (.Z(FE_PHN4973_U_afifo_U_acore_U_sub_fifo_n218), 
	.A(FE_PHN4114_U_afifo_U_acore_U_sub_fifo_n218));
   BUF_X1 FE_PHC4968_U_dfifo_U_dcore_U_sub_fifo_n266 (.Z(FE_PHN4968_U_dfifo_U_dcore_U_sub_fifo_n266), 
	.A(FE_PHN4103_U_dfifo_U_dcore_U_sub_fifo_n266));
   CLKBUF_X1 FE_PHC4965_U_afifo_U_acore_U_sub_fifo_n203 (.Z(FE_PHN4965_U_afifo_U_acore_U_sub_fifo_n203), 
	.A(FE_PHN3303_U_afifo_U_acore_U_sub_fifo_n203));
   CLKBUF_X1 FE_PHC4964_U_afifo_U_acore_U_sub_fifo_n240 (.Z(FE_PHN4964_U_afifo_U_acore_U_sub_fifo_n240), 
	.A(FE_PHN3992_U_afifo_U_acore_U_sub_fifo_n240));
   CLKBUF_X1 FE_PHC4961_U_dfifo_U_dcore_U_sub_fifo_n291 (.Z(FE_PHN4961_U_dfifo_U_dcore_U_sub_fifo_n291), 
	.A(FE_PHN4156_U_dfifo_U_dcore_U_sub_fifo_n291));
   CLKBUF_X1 FE_PHC4957_U_afifo_n192 (.Z(FE_PHN4957_U_afifo_n192), 
	.A(U_afifo_n192));
   CLKBUF_X2 FE_PHC4951_U_afifo_U_acore_U_sub_fifo_n229 (.Z(FE_PHN4951_U_afifo_U_acore_U_sub_fifo_n229), 
	.A(FE_PHN3994_U_afifo_U_acore_U_sub_fifo_n229));
   BUF_X1 FE_PHC4948_U_dfifo_U_dcore_U_sub_fifo_n261 (.Z(FE_PHN4948_U_dfifo_U_dcore_U_sub_fifo_n261), 
	.A(FE_PHN4116_U_dfifo_U_dcore_U_sub_fifo_n261));
   CLKBUF_X1 FE_PHC4945_U_dfifo_U_dcore_n151 (.Z(FE_PHN4945_U_dfifo_U_dcore_n151), 
	.A(FE_PHN3873_U_dfifo_U_dcore_n151));
   CLKBUF_X1 FE_PHC4942_U_afifo_U_acore_U_sub_fifo_n258 (.Z(FE_PHN4942_U_afifo_U_acore_U_sub_fifo_n258), 
	.A(FE_PHN3979_U_afifo_U_acore_U_sub_fifo_n258));
   CLKBUF_X1 FE_PHC4939_U_dfifo_U_dcore_U_sub_fifo_n253 (.Z(FE_PHN4939_U_dfifo_U_dcore_U_sub_fifo_n253), 
	.A(FE_PHN4137_U_dfifo_U_dcore_U_sub_fifo_n253));
   CLKBUF_X1 FE_PHC4936_U_afifo_U_acore_U_sub_fifo_n222 (.Z(FE_PHN4936_U_afifo_U_acore_U_sub_fifo_n222), 
	.A(FE_PHN3990_U_afifo_U_acore_U_sub_fifo_n222));
   CLKBUF_X1 FE_PHC4929_U_dfifo_U_dcore_U_sub_fifo_n210 (.Z(FE_PHN4929_U_dfifo_U_dcore_U_sub_fifo_n210), 
	.A(FE_PHN3933_U_dfifo_U_dcore_U_sub_fifo_n210));
   BUF_X1 FE_PHC4928_U_dfifo_U_dcore_n157 (.Z(FE_PHN4928_U_dfifo_U_dcore_n157), 
	.A(FE_PHN3236_U_dfifo_U_dcore_n157));
   BUF_X1 FE_PHC4926_U_dfifo_U_dcore_n154 (.Z(FE_PHN4926_U_dfifo_U_dcore_n154), 
	.A(FE_PHN4162_U_dfifo_U_dcore_n154));
   BUF_X1 FE_PHC4925_U_dfifo_U_dcore_U_sub_fifo_n267 (.Z(FE_PHN4925_U_dfifo_U_dcore_U_sub_fifo_n267), 
	.A(FE_PHN4144_U_dfifo_U_dcore_U_sub_fifo_n267));
   CLKBUF_X1 FE_PHC4918_U_dfifo_U_dcore_U_sub_fifo_n296 (.Z(FE_PHN4918_U_dfifo_U_dcore_U_sub_fifo_n296), 
	.A(FE_PHN4131_U_dfifo_U_dcore_U_sub_fifo_n296));
   CLKBUF_X1 FE_PHC4917_U_afifo_n191 (.Z(FE_PHN4917_U_afifo_n191), 
	.A(FE_PHN4086_U_afifo_n191));
   CLKBUF_X1 FE_PHC4908_U_dfifo_U_dcore_U_sub_fifo_n216 (.Z(FE_PHN4908_U_dfifo_U_dcore_U_sub_fifo_n216), 
	.A(FE_PHN3894_U_dfifo_U_dcore_U_sub_fifo_n216));
   CLKBUF_X1 FE_PHC4903_U_dfifo_U_dcore_U_sub_fifo_n164 (.Z(FE_PHN4903_U_dfifo_U_dcore_U_sub_fifo_n164), 
	.A(FE_PHN3913_U_dfifo_U_dcore_U_sub_fifo_n164));
   CLKBUF_X1 FE_PHC4901_U_dfifo_U_dcore_n155 (.Z(FE_PHN4901_U_dfifo_U_dcore_n155), 
	.A(FE_PHN3226_U_dfifo_U_dcore_n155));
   BUF_X1 FE_PHC4899_U_afifo_U_acore_U_sub_fifo_n256 (.Z(FE_PHN4899_U_afifo_U_acore_U_sub_fifo_n256), 
	.A(FE_PHN3489_U_afifo_U_acore_U_sub_fifo_n256));
   CLKBUF_X1 FE_PHC4892_U_dfifo_U_dcore_U_sub_fifo_n202 (.Z(FE_PHN4892_U_dfifo_U_dcore_U_sub_fifo_n202), 
	.A(FE_PHN3852_U_dfifo_U_dcore_U_sub_fifo_n202));
   CLKBUF_X1 FE_PHC4889_U_dfifo_U_dcore_U_sub_fifo_n314 (.Z(FE_PHN4889_U_dfifo_U_dcore_U_sub_fifo_n314), 
	.A(FE_PHN3840_U_dfifo_U_dcore_U_sub_fifo_n314));
   CLKBUF_X1 FE_PHC4881_U_dfifo_U_dcore_U_sub_fifo_n256 (.Z(FE_PHN4881_U_dfifo_U_dcore_U_sub_fifo_n256), 
	.A(FE_PHN4062_U_dfifo_U_dcore_U_sub_fifo_n256));
   CLKBUF_X1 FE_PHC4880_U_dfifo_U_dcore_U_sub_fifo_n174 (.Z(FE_PHN4880_U_dfifo_U_dcore_U_sub_fifo_n174), 
	.A(FE_PHN3832_U_dfifo_U_dcore_U_sub_fifo_n174));
   BUF_X1 FE_PHC4879_U_dfifo_U_dcore_U_sub_fifo_n176 (.Z(FE_PHN4879_U_dfifo_U_dcore_U_sub_fifo_n176), 
	.A(FE_PHN3812_U_dfifo_U_dcore_U_sub_fifo_n176));
   CLKBUF_X1 FE_PHC4877_U_afifo_U_acore_U_sub_fifo_n320 (.Z(FE_PHN4877_U_afifo_U_acore_U_sub_fifo_n320), 
	.A(FE_PHN4037_U_afifo_U_acore_U_sub_fifo_n320));
   CLKBUF_X1 FE_PHC4875_U_dfifo_U_dcore_U_sub_fifo_n172 (.Z(FE_PHN4875_U_dfifo_U_dcore_U_sub_fifo_n172), 
	.A(FE_PHN3807_U_dfifo_U_dcore_U_sub_fifo_n172));
   CLKBUF_X1 FE_PHC4872_U_dfifo_U_dcore_U_sub_fifo_n163 (.Z(FE_PHN4872_U_dfifo_U_dcore_U_sub_fifo_n163), 
	.A(FE_PHN3859_U_dfifo_U_dcore_U_sub_fifo_n163));
   CLKBUF_X1 FE_PHC4858_U_afifo_U_acore_U_sub_fifo_n214 (.Z(FE_PHN4858_U_afifo_U_acore_U_sub_fifo_n214), 
	.A(FE_PHN4087_U_afifo_U_acore_U_sub_fifo_n214));
   CLKBUF_X1 FE_PHC4856_U_dfifo_U_dcore_U_sub_fifo_n413 (.Z(FE_PHN4856_U_dfifo_U_dcore_U_sub_fifo_n413), 
	.A(FE_PHN3822_U_dfifo_U_dcore_U_sub_fifo_n413));
   CLKBUF_X1 FE_PHC4852_U_dfifo_U_dcore_U_sub_fifo_n207 (.Z(FE_PHN4852_U_dfifo_U_dcore_U_sub_fifo_n207), 
	.A(FE_PHN3841_U_dfifo_U_dcore_U_sub_fifo_n207));
   CLKBUF_X1 FE_PHC4848_U_dfifo_U_dcore_U_sub_fifo_n179 (.Z(FE_PHN4848_U_dfifo_U_dcore_U_sub_fifo_n179), 
	.A(FE_PHN4064_U_dfifo_U_dcore_U_sub_fifo_n179));
   CLKBUF_X1 FE_PHC4846_U_dfifo_U_dcore_U_sub_fifo_n166 (.Z(FE_PHN4846_U_dfifo_U_dcore_U_sub_fifo_n166), 
	.A(FE_PHN3848_U_dfifo_U_dcore_U_sub_fifo_n166));
   CLKBUF_X1 FE_PHC4843_U_dfifo_U_dcore_U_sub_fifo_n298 (.Z(FE_PHN4843_U_dfifo_U_dcore_U_sub_fifo_n298), 
	.A(FE_PHN4008_U_dfifo_U_dcore_U_sub_fifo_n298));
   CLKBUF_X1 FE_PHC4837_U_dfifo_U_dcore_U_sub_fifo_n214 (.Z(FE_PHN4837_U_dfifo_U_dcore_U_sub_fifo_n214), 
	.A(FE_PHN3861_U_dfifo_U_dcore_U_sub_fifo_n214));
   CLKBUF_X1 FE_PHC4836_U_dfifo_U_dcore_U_sub_fifo_n212 (.Z(FE_PHN4836_U_dfifo_U_dcore_U_sub_fifo_n212), 
	.A(FE_PHN3815_U_dfifo_U_dcore_U_sub_fifo_n212));
   CLKBUF_X1 FE_PHC4832_U_dfifo_U_dcore_U_sub_fifo_n338 (.Z(FE_PHN4832_U_dfifo_U_dcore_U_sub_fifo_n338), 
	.A(FE_PHN3790_U_dfifo_U_dcore_U_sub_fifo_n338));
   CLKBUF_X1 FE_PHC4826_U_dfifo_U_dcore_U_sub_fifo_n169 (.Z(FE_PHN4826_U_dfifo_U_dcore_U_sub_fifo_n169), 
	.A(FE_PHN3835_U_dfifo_U_dcore_U_sub_fifo_n169));
   CLKBUF_X1 FE_PHC4825_U_dfifo_U_dcore_U_sub_fifo_n168 (.Z(FE_PHN4825_U_dfifo_U_dcore_U_sub_fifo_n168), 
	.A(FE_PHN3824_U_dfifo_U_dcore_U_sub_fifo_n168));
   CLKBUF_X1 FE_PHC4824_U_dfifo_U_dcore_U_sub_fifo_n445 (.Z(FE_PHN4824_U_dfifo_U_dcore_U_sub_fifo_n445), 
	.A(FE_PHN3825_U_dfifo_U_dcore_U_sub_fifo_n445));
   CLKBUF_X1 FE_PHC4819_U_afifo_U_acore_U_sub_fifo_n267 (.Z(FE_PHN4819_U_afifo_U_acore_U_sub_fifo_n267), 
	.A(FE_PHN3817_U_afifo_U_acore_U_sub_fifo_n267));
   CLKBUF_X1 FE_PHC4817_U_dfifo_U_dcore_U_sub_fifo_n218 (.Z(FE_PHN4817_U_dfifo_U_dcore_U_sub_fifo_n218), 
	.A(FE_PHN3860_U_dfifo_U_dcore_U_sub_fifo_n218));
   CLKBUF_X1 FE_PHC4816_U_dfifo_U_dcore_U_sub_fifo_n209 (.Z(FE_PHN4816_U_dfifo_U_dcore_U_sub_fifo_n209), 
	.A(FE_PHN3858_U_dfifo_U_dcore_U_sub_fifo_n209));
   BUF_X1 FE_PHC4812_U_dfifo_U_dcore_U_sub_fifo_n450 (.Z(FE_PHN4812_U_dfifo_U_dcore_U_sub_fifo_n450), 
	.A(FE_PHN3295_U_dfifo_U_dcore_U_sub_fifo_n450));
   CLKBUF_X1 FE_PHC4811_U_dfifo_U_dcore_U_sub_fifo_n165 (.Z(FE_PHN4811_U_dfifo_U_dcore_U_sub_fifo_n165), 
	.A(FE_PHN3819_U_dfifo_U_dcore_U_sub_fifo_n165));
   CLKBUF_X1 FE_PHC4806_U_dfifo_U_dcore_U_sub_fifo_n401 (.Z(FE_PHN4806_U_dfifo_U_dcore_U_sub_fifo_n401), 
	.A(FE_PHN3791_U_dfifo_U_dcore_U_sub_fifo_n401));
   CLKBUF_X1 FE_PHC4803_U_dfifo_U_dcore_U_sub_fifo_n170 (.Z(FE_PHN4803_U_dfifo_U_dcore_U_sub_fifo_n170), 
	.A(FE_PHN3932_U_dfifo_U_dcore_U_sub_fifo_n170));
   CLKBUF_X1 FE_PHC4800_U_dfifo_U_dcore_U_sub_fifo_n173 (.Z(FE_PHN4800_U_dfifo_U_dcore_U_sub_fifo_n173), 
	.A(FE_PHN3818_U_dfifo_U_dcore_U_sub_fifo_n173));
   CLKBUF_X1 FE_PHC4799_U_dfifo_U_dcore_U_sub_fifo_n175 (.Z(FE_PHN4799_U_dfifo_U_dcore_U_sub_fifo_n175), 
	.A(FE_PHN3849_U_dfifo_U_dcore_U_sub_fifo_n175));
   CLKBUF_X1 FE_PHC4793_U_afifo_U_acore_U_sub_fifo_n266 (.Z(FE_PHN4793_U_afifo_U_acore_U_sub_fifo_n266), 
	.A(FE_PHN3795_U_afifo_U_acore_U_sub_fifo_n266));
   CLKBUF_X1 FE_PHC4791_U_dfifo_U_dcore_U_sub_fifo_n205 (.Z(FE_PHN4791_U_dfifo_U_dcore_U_sub_fifo_n205), 
	.A(FE_PHN3964_U_dfifo_U_dcore_U_sub_fifo_n205));
   CLKBUF_X1 FE_PHC4789_U_afifo_U_acore_U_sub_fifo_n296 (.Z(FE_PHN4789_U_afifo_U_acore_U_sub_fifo_n296), 
	.A(FE_PHN3163_U_afifo_U_acore_U_sub_fifo_n296));
   CLKBUF_X1 FE_PHC4786_U_dfifo_U_dcore_U_sub_fifo_n211 (.Z(FE_PHN4786_U_dfifo_U_dcore_U_sub_fifo_n211), 
	.A(FE_PHN3846_U_dfifo_U_dcore_U_sub_fifo_n211));
   CLKBUF_X1 FE_PHC4780_U_dfifo_U_dcore_n145 (.Z(FE_PHN4780_U_dfifo_U_dcore_n145), 
	.A(FE_PHN3219_U_dfifo_U_dcore_n145));
   CLKBUF_X1 FE_PHC4773_U_dfifo_U_dcore_U_sub_fifo_n215 (.Z(FE_PHN4773_U_dfifo_U_dcore_U_sub_fifo_n215), 
	.A(FE_PHN3855_U_dfifo_U_dcore_U_sub_fifo_n215));
   CLKBUF_X1 FE_PHC4771_U_dfifo_U_dcore_U_sub_fifo_n219 (.Z(FE_PHN4771_U_dfifo_U_dcore_U_sub_fifo_n219), 
	.A(FE_PHN3854_U_dfifo_U_dcore_U_sub_fifo_n219));
   CLKBUF_X1 FE_PHC4770_U_dfifo_U_dcore_U_sub_fifo_n344 (.Z(FE_PHN4770_U_dfifo_U_dcore_U_sub_fifo_n344), 
	.A(FE_PHN3767_U_dfifo_U_dcore_U_sub_fifo_n344));
   CLKBUF_X1 FE_PHC4769_U_dfifo_U_dcore_U_sub_fifo_n333 (.Z(FE_PHN4769_U_dfifo_U_dcore_U_sub_fifo_n333), 
	.A(FE_PHN3783_U_dfifo_U_dcore_U_sub_fifo_n333));
   CLKBUF_X1 FE_PHC4768_U_dfifo_U_dcore_U_sub_fifo_n403 (.Z(FE_PHN4768_U_dfifo_U_dcore_U_sub_fifo_n403), 
	.A(FE_PHN3747_U_dfifo_U_dcore_U_sub_fifo_n403));
   CLKBUF_X1 FE_PHC4766_U_dfifo_U_dcore_U_sub_fifo_n397 (.Z(FE_PHN4766_U_dfifo_U_dcore_U_sub_fifo_n397), 
	.A(FE_PHN3746_U_dfifo_U_dcore_U_sub_fifo_n397));
   CLKBUF_X1 FE_PHC4765_U_dfifo_U_dcore_U_sub_fifo_n398 (.Z(FE_PHN4765_U_dfifo_U_dcore_U_sub_fifo_n398), 
	.A(FE_PHN3740_U_dfifo_U_dcore_U_sub_fifo_n398));
   CLKBUF_X1 FE_PHC4764_U_dfifo_U_dcore_U_sub_fifo_n208 (.Z(FE_PHN4764_U_dfifo_U_dcore_U_sub_fifo_n208), 
	.A(FE_PHN3734_U_dfifo_U_dcore_U_sub_fifo_n208));
   CLKBUF_X1 FE_PHC4762_U_dfifo_U_dcore_U_sub_fifo_n220 (.Z(FE_PHN4762_U_dfifo_U_dcore_U_sub_fifo_n220), 
	.A(FE_PHN3820_U_dfifo_U_dcore_U_sub_fifo_n220));
   CLKBUF_X1 FE_PHC4758_U_afifo_U_acore_U_sub_fifo_n269 (.Z(FE_PHN4758_U_afifo_U_acore_U_sub_fifo_n269), 
	.A(FE_PHN3285_U_afifo_U_acore_U_sub_fifo_n269));
   CLKBUF_X1 FE_PHC4757_U_dfifo_U_dcore_U_sub_fifo_n206 (.Z(FE_PHN4757_U_dfifo_U_dcore_U_sub_fifo_n206), 
	.A(FE_PHN3834_U_dfifo_U_dcore_U_sub_fifo_n206));
   CLKBUF_X1 FE_PHC4755_U_dfifo_U_dcore_U_sub_fifo_n442 (.Z(FE_PHN4755_U_dfifo_U_dcore_U_sub_fifo_n442), 
	.A(FE_PHN3731_U_dfifo_U_dcore_U_sub_fifo_n442));
   CLKBUF_X1 FE_PHC4754_U_dfifo_U_dcore_U_sub_fifo_n356 (.Z(FE_PHN4754_U_dfifo_U_dcore_U_sub_fifo_n356), 
	.A(FE_PHN3729_U_dfifo_U_dcore_U_sub_fifo_n356));
   CLKBUF_X1 FE_PHC4753_U_dfifo_U_dcore_U_sub_fifo_n167 (.Z(FE_PHN4753_U_dfifo_U_dcore_U_sub_fifo_n167), 
	.A(FE_PHN3749_U_dfifo_U_dcore_U_sub_fifo_n167));
   CLKBUF_X1 FE_PHC4752_U_dfifo_U_dcore_U_sub_fifo_n440 (.Z(FE_PHN4752_U_dfifo_U_dcore_U_sub_fifo_n440), 
	.A(FE_PHN3719_U_dfifo_U_dcore_U_sub_fifo_n440));
   CLKBUF_X1 FE_PHC4751_U_dfifo_U_dcore_U_sub_fifo_n327 (.Z(FE_PHN4751_U_dfifo_U_dcore_U_sub_fifo_n327), 
	.A(FE_PHN3708_U_dfifo_U_dcore_U_sub_fifo_n327));
   CLKBUF_X1 FE_PHC4747_U_dfifo_U_dcore_U_sub_fifo_n412 (.Z(FE_PHN4747_U_dfifo_U_dcore_U_sub_fifo_n412), 
	.A(FE_PHN3709_U_dfifo_U_dcore_U_sub_fifo_n412));
   CLKBUF_X1 FE_PHC4746_U_dfifo_U_dcore_U_sub_fifo_n320 (.Z(FE_PHN4746_U_dfifo_U_dcore_U_sub_fifo_n320), 
	.A(FE_PHN3700_U_dfifo_U_dcore_U_sub_fifo_n320));
   CLKBUF_X1 FE_PHC4745_U_dfifo_U_dcore_U_sub_fifo_n452 (.Z(FE_PHN4745_U_dfifo_U_dcore_U_sub_fifo_n452), 
	.A(FE_PHN3218_U_dfifo_U_dcore_U_sub_fifo_n452));
   CLKBUF_X1 FE_PHC4744_U_dfifo_U_dcore_U_sub_fifo_n402 (.Z(FE_PHN4744_U_dfifo_U_dcore_U_sub_fifo_n402), 
	.A(FE_PHN3720_U_dfifo_U_dcore_U_sub_fifo_n402));
   CLKBUF_X1 FE_PHC4742_U_dfifo_U_dcore_U_sub_fifo_n316 (.Z(FE_PHN4742_U_dfifo_U_dcore_U_sub_fifo_n316), 
	.A(FE_PHN3644_U_dfifo_U_dcore_U_sub_fifo_n316));
   CLKBUF_X1 FE_PHC4741_U_dfifo_U_dcore_U_sub_fifo_n204 (.Z(FE_PHN4741_U_dfifo_U_dcore_U_sub_fifo_n204), 
	.A(FE_PHN3805_U_dfifo_U_dcore_U_sub_fifo_n204));
   CLKBUF_X1 FE_PHC4740_U_dfifo_U_dcore_U_sub_fifo_n340 (.Z(FE_PHN4740_U_dfifo_U_dcore_U_sub_fifo_n340), 
	.A(FE_PHN3723_U_dfifo_U_dcore_U_sub_fifo_n340));
   CLKBUF_X1 FE_PHC4738_U_dfifo_U_dcore_U_sub_fifo_n446 (.Z(FE_PHN4738_U_dfifo_U_dcore_U_sub_fifo_n446), 
	.A(FE_PHN3673_U_dfifo_U_dcore_U_sub_fifo_n446));
   CLKBUF_X1 FE_PHC4719_U_afifo_U_acore_n97 (.Z(FE_PHN4719_U_afifo_U_acore_n97), 
	.A(FE_PHN3310_U_afifo_U_acore_n97));
   BUF_X32 FE_PHC4705_U_ctl_N89 (.Z(FE_PHN4705_U_ctl_N89), 
	.A(FE_PHN5218_U_ctl_N89));
   CLKBUF_X1 FE_PHC4677_U_afifo_U_acore_U_sub_fifo_n297 (.Z(FE_PHN4677_U_afifo_U_acore_U_sub_fifo_n297), 
	.A(FE_PHN3175_U_afifo_U_acore_U_sub_fifo_n297));
   BUF_X32 FE_PHC4665_U_rbuf_n69 (.Z(FE_PHN4665_U_rbuf_n69), 
	.A(FE_PHN5240_U_rbuf_n69));
   BUF_X32 FE_PHC4664_miu_data_27_ (.Z(FE_PHN4664_miu_data_27_), 
	.A(FE_PHN5191_miu_data_27_));
   BUF_X32 FE_PHC4663_U_rbuf_n175 (.Z(FE_PHN4663_U_rbuf_n175), 
	.A(FE_PHN5241_U_rbuf_n175));
   BUF_X8 FE_PHC4650_U_rbuf_n63 (.Z(FE_PHN4650_U_rbuf_n63), 
	.A(U_rbuf_n63));
   BUF_X16 FE_PHC4649_U_rbuf_n59 (.Z(FE_PHN4649_U_rbuf_n59), 
	.A(U_rbuf_n59));
   BUF_X16 FE_PHC4647_U_rbuf_n174 (.Z(FE_PHN4647_U_rbuf_n174), 
	.A(U_rbuf_n174));
   BUF_X32 FE_PHC4646_U_rbuf_n179 (.Z(FE_PHN4646_U_rbuf_n179), 
	.A(U_rbuf_n179));
   CLKBUF_X1 FE_PHC4644_U_rbuf_n182 (.Z(FE_PHN4644_U_rbuf_n182), 
	.A(U_rbuf_n182));
   BUF_X16 FE_PHC4643_U_rbuf_n56 (.Z(FE_PHN4643_U_rbuf_n56), 
	.A(U_rbuf_n56));
   CLKBUF_X1 FE_PHC4642_U_rbuf_n75 (.Z(FE_PHN4642_U_rbuf_n75), 
	.A(U_rbuf_n75));
   BUF_X32 FE_PHC4640_U_ctl_n_bh_state_0_ (.Z(FE_PHN4640_U_ctl_n_bh_state_0_), 
	.A(U_ctl_n_bh_state[0]));
   BUF_X8 FE_PHC4636_hsel_reg (.Z(FE_PHN4636_hsel_reg), 
	.A(FE_PHN2917_hsel_reg));
   CLKBUF_X1 FE_PHC4635_U_rbuf_n188 (.Z(FE_PHN4635_U_rbuf_n188), 
	.A(FE_PHN5175_U_rbuf_n188));
   BUF_X32 FE_PHC4633_U_ctl_n212 (.Z(FE_PHN4633_U_ctl_n212), 
	.A(U_ctl_n212));
   BUF_X32 FE_PHC4632_U_ctl_n_sel_buf (.Z(FE_PHN4632_U_ctl_n_sel_buf), 
	.A(U_ctl_n_sel_buf));
   BUF_X32 FE_PHC4628_U_ctl_n382 (.Z(FE_PHN4628_U_ctl_n382), 
	.A(U_ctl_n382));
   BUF_X32 FE_PHC4626_m_af_push1_n (.Z(FE_PHN4626_m_af_push1_n), 
	.A(m_af_push1_n));
   BUF_X32 FE_PHC4619_U_ctl_f_burst_done (.Z(FE_PHN4619_U_ctl_f_burst_done), 
	.A(U_ctl_f_burst_done));
   CLKBUF_X1 FE_PHC4384_U_dfifo_U_dcore_n_empty (.Z(FE_PHN4384_U_dfifo_U_dcore_n_empty), 
	.A(FE_PHN1660_U_dfifo_U_dcore_n_empty));
   CLKBUF_X1 FE_PHC4370_U_dfifo_U_dcore_U_sub_fifo_n272 (.Z(FE_PHN4370_U_dfifo_U_dcore_U_sub_fifo_n272), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n272));
   CLKBUF_X1 FE_PHC4347_U_dfifo_U_dcore_U_sub_fifo_n303 (.Z(FE_PHN4347_U_dfifo_U_dcore_U_sub_fifo_n303), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n303));
   CLKBUF_X1 FE_PHC4341_U_dfifo_U_dcore_U_sub_fifo_n262 (.Z(FE_PHN4341_U_dfifo_U_dcore_U_sub_fifo_n262), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n262));
   CLKBUF_X1 FE_PHC4321_U_dfifo_U_dcore_U_sub_fifo_n55 (.Z(FE_PHN4321_U_dfifo_U_dcore_U_sub_fifo_n55), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n55));
   CLKBUF_X1 FE_PHC4310_U_dfifo_U_dcore_U_sub_fifo_n258 (.Z(FE_PHN4310_U_dfifo_U_dcore_U_sub_fifo_n258), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n258));
   CLKBUF_X1 FE_PHC4309_U_dfifo_U_dcore_U_sub_fifo_n278 (.Z(FE_PHN4309_U_dfifo_U_dcore_U_sub_fifo_n278), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n278));
   CLKBUF_X1 FE_PHC4300_U_dfifo_U_dcore_U_sub_fifo_n306 (.Z(FE_PHN4300_U_dfifo_U_dcore_U_sub_fifo_n306), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n306));
   CLKBUF_X1 FE_PHC4299_U_dfifo_U_dcore_U_sub_fifo_n451 (.Z(FE_PHN4299_U_dfifo_U_dcore_U_sub_fifo_n451), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n451));
   CLKBUF_X1 FE_PHC4296_U_dfifo_U_dcore_U_sub_fifo_n276 (.Z(FE_PHN4296_U_dfifo_U_dcore_U_sub_fifo_n276), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n276));
   CLKBUF_X1 FE_PHC4294_U_dfifo_U_dcore_U_sub_fifo_n448 (.Z(FE_PHN4294_U_dfifo_U_dcore_U_sub_fifo_n448), 
	.A(FE_PHN2421_U_dfifo_U_dcore_U_sub_fifo_n448));
   CLKBUF_X1 FE_PHC4292_U_dfifo_U_dcore_U_sub_fifo_n271 (.Z(FE_PHN4292_U_dfifo_U_dcore_U_sub_fifo_n271), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n271));
   CLKBUF_X1 FE_PHC4290_U_dfifo_U_dcore_U_sub_fifo_n270 (.Z(FE_PHN4290_U_dfifo_U_dcore_U_sub_fifo_n270), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n270));
   CLKBUF_X1 FE_PHC4285_U_dfifo_U_dcore_U_sub_fifo_n294 (.Z(FE_PHN4285_U_dfifo_U_dcore_U_sub_fifo_n294), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n294));
   CLKBUF_X1 FE_PHC4284_U_dfifo_U_dcore_U_sub_fifo_n260 (.Z(FE_PHN4284_U_dfifo_U_dcore_U_sub_fifo_n260), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n260));
   CLKBUF_X1 FE_PHC4281_U_dfifo_U_dcore_U_sub_fifo_n264 (.Z(FE_PHN4281_U_dfifo_U_dcore_U_sub_fifo_n264), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n264));
   CLKBUF_X1 FE_PHC4278_U_dfifo_U_dcore_U_sub_fifo_n265 (.Z(FE_PHN4278_U_dfifo_U_dcore_U_sub_fifo_n265), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n265));
   CLKBUF_X1 FE_PHC4276_U_dfifo_U_dcore_U_sub_fifo_n283 (.Z(FE_PHN4276_U_dfifo_U_dcore_U_sub_fifo_n283), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n283));
   CLKBUF_X1 FE_PHC4275_U_dfifo_U_dcore_U_sub_fifo_n295 (.Z(FE_PHN4275_U_dfifo_U_dcore_U_sub_fifo_n295), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n295));
   CLKBUF_X1 FE_PHC4268_U_dfifo_U_dcore_U_sub_fifo_n277 (.Z(FE_PHN4268_U_dfifo_U_dcore_U_sub_fifo_n277), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n277));
   CLKBUF_X1 FE_PHC4256_U_dfifo_U_dcore_U_sub_fifo_n243 (.Z(FE_PHN4256_U_dfifo_U_dcore_U_sub_fifo_n243), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n243));
   CLKBUF_X1 FE_PHC4255_U_dfifo_U_dcore_U_sub_fifo_n259 (.Z(FE_PHN4255_U_dfifo_U_dcore_U_sub_fifo_n259), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n259));
   CLKBUF_X1 FE_PHC4254_U_dfifo_U_dcore_U_sub_fifo_n282 (.Z(FE_PHN4254_U_dfifo_U_dcore_U_sub_fifo_n282), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n282));
   CLKBUF_X1 FE_PHC4253_U_dfifo_U_dcore_U_sub_fifo_n268 (.Z(FE_PHN4253_U_dfifo_U_dcore_U_sub_fifo_n268), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n268));
   CLKBUF_X1 FE_PHC4252_U_dfifo_U_dcore_U_sub_fifo_n309 (.Z(FE_PHN4252_U_dfifo_U_dcore_U_sub_fifo_n309), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n309));
   CLKBUF_X1 FE_PHC4251_U_dfifo_U_dcore_U_sub_fifo_n250 (.Z(FE_PHN4251_U_dfifo_U_dcore_U_sub_fifo_n250), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n250));
   CLKBUF_X1 FE_PHC4250_U_dfifo_U_dcore_U_sub_fifo_n248 (.Z(FE_PHN4250_U_dfifo_U_dcore_U_sub_fifo_n248), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n248));
   CLKBUF_X1 FE_PHC4245_U_dfifo_U_dcore_U_sub_fifo_n269 (.Z(FE_PHN4245_U_dfifo_U_dcore_U_sub_fifo_n269), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n269));
   CLKBUF_X1 FE_PHC4244_U_dfifo_U_dcore_U_sub_fifo_n299 (.Z(FE_PHN4244_U_dfifo_U_dcore_U_sub_fifo_n299), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n299));
   CLKBUF_X1 FE_PHC4243_U_dfifo_U_dcore_U_sub_fifo_n305 (.Z(FE_PHN4243_U_dfifo_U_dcore_U_sub_fifo_n305), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n305));
   CLKBUF_X1 FE_PHC4242_U_dfifo_U_dcore_U_sub_fifo_n300 (.Z(FE_PHN4242_U_dfifo_U_dcore_U_sub_fifo_n300), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n300));
   CLKBUF_X1 FE_PHC4241_U_dfifo_U_dcore_U_sub_fifo_n286 (.Z(FE_PHN4241_U_dfifo_U_dcore_U_sub_fifo_n286), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n286));
   CLKBUF_X1 FE_PHC4239_U_dfifo_U_dcore_U_sub_fifo_n273 (.Z(FE_PHN4239_U_dfifo_U_dcore_U_sub_fifo_n273), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n273));
   CLKBUF_X1 FE_PHC4238_U_dfifo_U_dcore_U_sub_fifo_n284 (.Z(FE_PHN4238_U_dfifo_U_dcore_U_sub_fifo_n284), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n284));
   CLKBUF_X1 FE_PHC4236_U_dfifo_U_dcore_U_sub_fifo_n257 (.Z(FE_PHN4236_U_dfifo_U_dcore_U_sub_fifo_n257), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n257));
   CLKBUF_X1 FE_PHC4228_U_dfifo_U_dcore_U_sub_fifo_n254 (.Z(FE_PHN4228_U_dfifo_U_dcore_U_sub_fifo_n254), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n254));
   CLKBUF_X1 FE_PHC4226_U_afifo_U_acore_U_sub_fifo_n279 (.Z(FE_PHN4226_U_afifo_U_acore_U_sub_fifo_n279), 
	.A(U_afifo_U_acore_U_sub_fifo_n279));
   CLKBUF_X1 FE_PHC4225_U_dfifo_U_dcore_U_sub_fifo_n310 (.Z(FE_PHN4225_U_dfifo_U_dcore_U_sub_fifo_n310), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n310));
   CLKBUF_X1 FE_PHC4224_U_dfifo_U_dcore_U_sub_fifo_n293 (.Z(FE_PHN4224_U_dfifo_U_dcore_U_sub_fifo_n293), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n293));
   CLKBUF_X1 FE_PHC4223_U_afifo_U_acore_U_sub_fifo_n309 (.Z(FE_PHN4223_U_afifo_U_acore_U_sub_fifo_n309), 
	.A(U_afifo_U_acore_U_sub_fifo_n309));
   CLKBUF_X1 FE_PHC4222_U_dfifo_U_dcore_U_sub_fifo_n274 (.Z(FE_PHN4222_U_dfifo_U_dcore_U_sub_fifo_n274), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n274));
   CLKBUF_X1 FE_PHC4211_U_dfifo_U_dcore_U_sub_fifo_n292 (.Z(FE_PHN4211_U_dfifo_U_dcore_U_sub_fifo_n292), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n292));
   CLKBUF_X1 FE_PHC4210_U_dfifo_U_dcore_U_sub_fifo_n255 (.Z(FE_PHN4210_U_dfifo_U_dcore_U_sub_fifo_n255), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n255));
   CLKBUF_X1 FE_PHC4209_U_dfifo_U_dcore_U_sub_fifo_n288 (.Z(FE_PHN4209_U_dfifo_U_dcore_U_sub_fifo_n288), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n288));
   CLKBUF_X1 FE_PHC4208_U_dfifo_U_dcore_U_sub_fifo_n245 (.Z(FE_PHN4208_U_dfifo_U_dcore_U_sub_fifo_n245), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n245));
   CLKBUF_X1 FE_PHC4207_U_dfifo_U_dcore_n156 (.Z(FE_PHN4207_U_dfifo_U_dcore_n156), 
	.A(U_dfifo_U_dcore_n156));
   CLKBUF_X1 FE_PHC4206_U_dfifo_U_dcore_U_sub_fifo_n290 (.Z(FE_PHN4206_U_dfifo_U_dcore_U_sub_fifo_n290), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n290));
   CLKBUF_X1 FE_PHC4203_U_afifo_U_acore_U_sub_fifo_n196 (.Z(FE_PHN4203_U_afifo_U_acore_U_sub_fifo_n196), 
	.A(U_afifo_U_acore_U_sub_fifo_n196));
   BUF_X8 FE_PHC4197_U_afifo_U_acore_U_sub_fifo_n208 (.Z(FE_PHN4197_U_afifo_U_acore_U_sub_fifo_n208), 
	.A(U_afifo_U_acore_U_sub_fifo_n208));
   CLKBUF_X1 FE_PHC4195_U_dfifo_U_dcore_U_sub_fifo_n308 (.Z(FE_PHN4195_U_dfifo_U_dcore_U_sub_fifo_n308), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n308));
   CLKBUF_X1 FE_PHC4194_U_dfifo_U_dcore_U_sub_fifo_n307 (.Z(FE_PHN4194_U_dfifo_U_dcore_U_sub_fifo_n307), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n307));
   CLKBUF_X1 FE_PHC4190_U_dfifo_U_dcore_U_sub_fifo_n285 (.Z(FE_PHN4190_U_dfifo_U_dcore_U_sub_fifo_n285), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n285));
   CLKBUF_X1 FE_PHC4189_U_dfifo_U_dcore_U_sub_fifo_n249 (.Z(FE_PHN4189_U_dfifo_U_dcore_U_sub_fifo_n249), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n249));
   CLKBUF_X1 FE_PHC4188_U_dfifo_U_dcore_U_sub_fifo_n280 (.Z(FE_PHN4188_U_dfifo_U_dcore_U_sub_fifo_n280), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n280));
   CLKBUF_X1 FE_PHC4186_U_afifo_n159 (.Z(FE_PHN4186_U_afifo_n159), 
	.A(U_afifo_n159));
   CLKBUF_X1 FE_PHC4184_U_dfifo_U_dcore_U_sub_fifo_n247 (.Z(FE_PHN4184_U_dfifo_U_dcore_U_sub_fifo_n247), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n247));
   CLKBUF_X1 FE_PHC4183_U_dfifo_U_dcore_U_sub_fifo_n246 (.Z(FE_PHN4183_U_dfifo_U_dcore_U_sub_fifo_n246), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n246));
   CLKBUF_X1 FE_PHC4179_U_afifo_U_acore_U_sub_fifo_n192 (.Z(FE_PHN4179_U_afifo_U_acore_U_sub_fifo_n192), 
	.A(U_afifo_U_acore_U_sub_fifo_n192));
   CLKBUF_X1 FE_PHC4173_U_dfifo_U_dcore_U_sub_fifo_n251 (.Z(FE_PHN4173_U_dfifo_U_dcore_U_sub_fifo_n251), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n251));
   CLKBUF_X1 FE_PHC4164_U_afifo_U_acore_U_sub_fifo_n275 (.Z(FE_PHN4164_U_afifo_U_acore_U_sub_fifo_n275), 
	.A(U_afifo_U_acore_U_sub_fifo_n275));
   CLKBUF_X1 FE_PHC4163_U_afifo_U_acore_U_sub_fifo_n205 (.Z(FE_PHN4163_U_afifo_U_acore_U_sub_fifo_n205), 
	.A(U_afifo_U_acore_U_sub_fifo_n205));
   CLKBUF_X1 FE_PHC4162_U_dfifo_U_dcore_n154 (.Z(FE_PHN4162_U_dfifo_U_dcore_n154), 
	.A(U_dfifo_U_dcore_n154));
   CLKBUF_X1 FE_PHC4159_U_afifo_U_acore_U_sub_fifo_n187 (.Z(FE_PHN4159_U_afifo_U_acore_U_sub_fifo_n187), 
	.A(U_afifo_U_acore_U_sub_fifo_n187));
   CLKBUF_X1 FE_PHC4158_U_afifo_U_acore_U_sub_fifo_n191 (.Z(FE_PHN4158_U_afifo_U_acore_U_sub_fifo_n191), 
	.A(U_afifo_U_acore_U_sub_fifo_n191));
   CLKBUF_X1 FE_PHC4157_U_dfifo_U_dcore_U_sub_fifo_n275 (.Z(FE_PHN4157_U_dfifo_U_dcore_U_sub_fifo_n275), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n275));
   CLKBUF_X1 FE_PHC4156_U_dfifo_U_dcore_U_sub_fifo_n291 (.Z(FE_PHN4156_U_dfifo_U_dcore_U_sub_fifo_n291), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n291));
   CLKBUF_X1 FE_PHC4155_U_dfifo_U_dcore_n153 (.Z(FE_PHN4155_U_dfifo_U_dcore_n153), 
	.A(U_dfifo_U_dcore_n153));
   CLKBUF_X1 FE_PHC4153_U_afifo_U_acore_U_sub_fifo_n184 (.Z(FE_PHN4153_U_afifo_U_acore_U_sub_fifo_n184), 
	.A(U_afifo_U_acore_U_sub_fifo_n184));
   CLKBUF_X1 FE_PHC4151_U_dfifo_U_dcore_U_sub_fifo_n304 (.Z(FE_PHN4151_U_dfifo_U_dcore_U_sub_fifo_n304), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n304));
   CLKBUF_X1 FE_PHC4144_U_dfifo_U_dcore_U_sub_fifo_n267 (.Z(FE_PHN4144_U_dfifo_U_dcore_U_sub_fifo_n267), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n267));
   CLKBUF_X1 FE_PHC4143_U_dfifo_U_dcore_U_sub_fifo_n279 (.Z(FE_PHN4143_U_dfifo_U_dcore_U_sub_fifo_n279), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n279));
   CLKBUF_X1 FE_PHC4137_U_dfifo_U_dcore_U_sub_fifo_n253 (.Z(FE_PHN4137_U_dfifo_U_dcore_U_sub_fifo_n253), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n253));
   CLKBUF_X1 FE_PHC4134_U_afifo_U_acore_U_sub_fifo_n210 (.Z(FE_PHN4134_U_afifo_U_acore_U_sub_fifo_n210), 
	.A(U_afifo_U_acore_U_sub_fifo_n210));
   CLKBUF_X1 FE_PHC4131_U_dfifo_U_dcore_U_sub_fifo_n296 (.Z(FE_PHN4131_U_dfifo_U_dcore_U_sub_fifo_n296), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n296));
   CLKBUF_X1 FE_PHC4130_U_dfifo_U_dcore_U_sub_fifo_n281 (.Z(FE_PHN4130_U_dfifo_U_dcore_U_sub_fifo_n281), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n281));
   CLKBUF_X1 FE_PHC4128_U_afifo_U_acore_U_sub_fifo_n188 (.Z(FE_PHN4128_U_afifo_U_acore_U_sub_fifo_n188), 
	.A(U_afifo_U_acore_U_sub_fifo_n188));
   CLKBUF_X1 FE_PHC4127_U_afifo_U_acore_U_sub_fifo_n291 (.Z(FE_PHN4127_U_afifo_U_acore_U_sub_fifo_n291), 
	.A(U_afifo_U_acore_U_sub_fifo_n291));
   CLKBUF_X1 FE_PHC4125_U_dfifo_U_dcore_U_sub_fifo_n263 (.Z(FE_PHN4125_U_dfifo_U_dcore_U_sub_fifo_n263), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n263));
   CLKBUF_X1 FE_PHC4121_U_afifo_U_acore_U_sub_fifo_n265 (.Z(FE_PHN4121_U_afifo_U_acore_U_sub_fifo_n265), 
	.A(U_afifo_U_acore_U_sub_fifo_n265));
   CLKBUF_X1 FE_PHC4116_U_dfifo_U_dcore_U_sub_fifo_n261 (.Z(FE_PHN4116_U_dfifo_U_dcore_U_sub_fifo_n261), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n261));
   CLKBUF_X1 FE_PHC4114_U_afifo_U_acore_U_sub_fifo_n218 (.Z(FE_PHN4114_U_afifo_U_acore_U_sub_fifo_n218), 
	.A(U_afifo_U_acore_U_sub_fifo_n218));
   CLKBUF_X1 FE_PHC4113_U_afifo_U_acore_U_sub_fifo_n314 (.Z(FE_PHN4113_U_afifo_U_acore_U_sub_fifo_n314), 
	.A(U_afifo_U_acore_U_sub_fifo_n314));
   BUF_X8 FE_PHC4112_U_afifo_U_acore_U_sub_fifo_n317 (.Z(FE_PHN4112_U_afifo_U_acore_U_sub_fifo_n317), 
	.A(U_afifo_U_acore_U_sub_fifo_n317));
   CLKBUF_X1 FE_PHC4111_U_afifo_U_acore_U_sub_fifo_n180 (.Z(FE_PHN4111_U_afifo_U_acore_U_sub_fifo_n180), 
	.A(U_afifo_U_acore_U_sub_fifo_n180));
   BUF_X8 FE_PHC4107_U_afifo_U_acore_U_sub_fifo_n190 (.Z(FE_PHN4107_U_afifo_U_acore_U_sub_fifo_n190), 
	.A(U_afifo_U_acore_U_sub_fifo_n190));
   CLKBUF_X1 FE_PHC4106_U_afifo_U_acore_U_sub_fifo_n285 (.Z(FE_PHN4106_U_afifo_U_acore_U_sub_fifo_n285), 
	.A(U_afifo_U_acore_U_sub_fifo_n285));
   CLKBUF_X1 FE_PHC4105_U_afifo_n17 (.Z(FE_PHN4105_U_afifo_n17), 
	.A(U_afifo_n17));
   CLKBUF_X1 FE_PHC4103_U_dfifo_U_dcore_U_sub_fifo_n266 (.Z(FE_PHN4103_U_dfifo_U_dcore_U_sub_fifo_n266), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n266));
   BUF_X8 FE_PHC4100_U_afifo_U_acore_U_sub_fifo_n263 (.Z(FE_PHN4100_U_afifo_U_acore_U_sub_fifo_n263), 
	.A(U_afifo_U_acore_U_sub_fifo_n263));
   CLKBUF_X1 FE_PHC4099_U_afifo_U_acore_U_sub_fifo_n264 (.Z(FE_PHN4099_U_afifo_U_acore_U_sub_fifo_n264), 
	.A(U_afifo_U_acore_U_sub_fifo_n264));
   CLKBUF_X1 FE_PHC4098_U_afifo_U_acore_U_sub_fifo_n283 (.Z(FE_PHN4098_U_afifo_U_acore_U_sub_fifo_n283), 
	.A(U_afifo_U_acore_U_sub_fifo_n283));
   BUF_X8 FE_PHC4097_U_afifo_U_acore_U_sub_fifo_n284 (.Z(FE_PHN4097_U_afifo_U_acore_U_sub_fifo_n284), 
	.A(U_afifo_U_acore_U_sub_fifo_n284));
   CLKBUF_X1 FE_PHC4095_U_dfifo_U_dcore_U_sub_fifo_n287 (.Z(FE_PHN4095_U_dfifo_U_dcore_U_sub_fifo_n287), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n287));
   BUF_X8 FE_PHC4092_U_afifo_U_acore_U_sub_fifo_n288 (.Z(FE_PHN4092_U_afifo_U_acore_U_sub_fifo_n288), 
	.A(U_afifo_U_acore_U_sub_fifo_n288));
   BUF_X8 FE_PHC4091_U_dfifo_U_dcore_U_sub_fifo_n289 (.Z(FE_PHN4091_U_dfifo_U_dcore_U_sub_fifo_n289), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n289));
   CLKBUF_X1 FE_PHC4087_U_afifo_U_acore_U_sub_fifo_n214 (.Z(FE_PHN4087_U_afifo_U_acore_U_sub_fifo_n214), 
	.A(U_afifo_U_acore_U_sub_fifo_n214));
   CLKBUF_X1 FE_PHC4086_U_afifo_n191 (.Z(FE_PHN4086_U_afifo_n191), 
	.A(U_afifo_n191));
   CLKBUF_X1 FE_PHC4081_U_afifo_U_acore_U_sub_fifo_n213 (.Z(FE_PHN4081_U_afifo_U_acore_U_sub_fifo_n213), 
	.A(U_afifo_U_acore_U_sub_fifo_n213));
   BUF_X8 FE_PHC4080_U_afifo_U_acore_U_sub_fifo_n230 (.Z(FE_PHN4080_U_afifo_U_acore_U_sub_fifo_n230), 
	.A(U_afifo_U_acore_U_sub_fifo_n230));
   BUF_X1 FE_PHC4079_U_afifo_n166 (.Z(FE_PHN4079_U_afifo_n166), 
	.A(U_afifo_n166));
   BUF_X8 FE_PHC4074_U_afifo_U_acore_U_sub_fifo_n232 (.Z(FE_PHN4074_U_afifo_U_acore_U_sub_fifo_n232), 
	.A(U_afifo_U_acore_U_sub_fifo_n232));
   CLKBUF_X1 FE_PHC4073_U_dfifo_U_dcore_U_sub_fifo_n297 (.Z(FE_PHN4073_U_dfifo_U_dcore_U_sub_fifo_n297), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n297));
   BUF_X8 FE_PHC4071_U_afifo_U_acore_U_sub_fifo_n224 (.Z(FE_PHN4071_U_afifo_U_acore_U_sub_fifo_n224), 
	.A(U_afifo_U_acore_U_sub_fifo_n224));
   BUF_X8 FE_PHC4070_U_afifo_U_acore_U_sub_fifo_n181 (.Z(FE_PHN4070_U_afifo_U_acore_U_sub_fifo_n181), 
	.A(U_afifo_U_acore_U_sub_fifo_n181));
   CLKBUF_X1 FE_PHC4069_U_afifo_U_acore_U_sub_fifo_n315 (.Z(FE_PHN4069_U_afifo_U_acore_U_sub_fifo_n315), 
	.A(U_afifo_U_acore_U_sub_fifo_n315));
   BUF_X8 FE_PHC4068_U_dfifo_U_dcore_U_sub_fifo_n301 (.Z(FE_PHN4068_U_dfifo_U_dcore_U_sub_fifo_n301), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n301));
   BUF_X8 FE_PHC4066_U_afifo_U_acore_U_sub_fifo_n178 (.Z(FE_PHN4066_U_afifo_U_acore_U_sub_fifo_n178), 
	.A(U_afifo_U_acore_U_sub_fifo_n178));
   BUF_X8 FE_PHC4065_U_afifo_U_acore_U_sub_fifo_n175 (.Z(FE_PHN4065_U_afifo_U_acore_U_sub_fifo_n175), 
	.A(U_afifo_U_acore_U_sub_fifo_n175));
   CLKBUF_X1 FE_PHC4064_U_dfifo_U_dcore_U_sub_fifo_n179 (.Z(FE_PHN4064_U_dfifo_U_dcore_U_sub_fifo_n179), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n179));
   BUF_X8 FE_PHC4063_U_dfifo_U_dcore_U_sub_fifo_n244 (.Z(FE_PHN4063_U_dfifo_U_dcore_U_sub_fifo_n244), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n244));
   CLKBUF_X1 FE_PHC4062_U_dfifo_U_dcore_U_sub_fifo_n256 (.Z(FE_PHN4062_U_dfifo_U_dcore_U_sub_fifo_n256), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n256));
   BUF_X8 FE_PHC4056_U_afifo_U_acore_U_sub_fifo_n215 (.Z(FE_PHN4056_U_afifo_U_acore_U_sub_fifo_n215), 
	.A(U_afifo_U_acore_U_sub_fifo_n215));
   BUF_X8 FE_PHC4055_U_afifo_U_acore_U_sub_fifo_n290 (.Z(FE_PHN4055_U_afifo_U_acore_U_sub_fifo_n290), 
	.A(U_afifo_U_acore_U_sub_fifo_n290));
   CLKBUF_X1 FE_PHC4049_U_afifo_U_acore_U_sub_fifo_n247 (.Z(FE_PHN4049_U_afifo_U_acore_U_sub_fifo_n247), 
	.A(U_afifo_U_acore_U_sub_fifo_n247));
   BUF_X8 FE_PHC4046_U_dfifo_U_dcore_n150 (.Z(FE_PHN4046_U_dfifo_U_dcore_n150), 
	.A(U_dfifo_U_dcore_n150));
   BUF_X8 FE_PHC4038_U_afifo_U_acore_U_sub_fifo_n259 (.Z(FE_PHN4038_U_afifo_U_acore_U_sub_fifo_n259), 
	.A(U_afifo_U_acore_U_sub_fifo_n259));
   CLKBUF_X1 FE_PHC4037_U_afifo_U_acore_U_sub_fifo_n320 (.Z(FE_PHN4037_U_afifo_U_acore_U_sub_fifo_n320), 
	.A(U_afifo_U_acore_U_sub_fifo_n320));
   BUF_X8 FE_PHC4036_U_afifo_U_acore_U_sub_fifo_n197 (.Z(FE_PHN4036_U_afifo_U_acore_U_sub_fifo_n197), 
	.A(U_afifo_U_acore_U_sub_fifo_n197));
   CLKBUF_X1 FE_PHC4033_U_dfifo_U_dcore_U_sub_fifo_n302 (.Z(FE_PHN4033_U_dfifo_U_dcore_U_sub_fifo_n302), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n302));
   BUF_X8 FE_PHC4030_U_afifo_U_acore_U_sub_fifo_n257 (.Z(FE_PHN4030_U_afifo_U_acore_U_sub_fifo_n257), 
	.A(U_afifo_U_acore_U_sub_fifo_n257));
   CLKBUF_X1 FE_PHC4028_U_afifo_n192 (.Z(FE_PHN4028_U_afifo_n192), 
	.A(FE_PHN4957_U_afifo_n192));
   CLKBUF_X1 FE_PHC4025_U_afifo_n165 (.Z(FE_PHN4025_U_afifo_n165), 
	.A(U_afifo_n165));
   BUF_X8 FE_PHC4019_U_afifo_U_acore_U_sub_fifo_n304 (.Z(FE_PHN4019_U_afifo_U_acore_U_sub_fifo_n304), 
	.A(U_afifo_U_acore_U_sub_fifo_n304));
   BUF_X8 FE_PHC4016_U_afifo_U_acore_U_sub_fifo_n211 (.Z(FE_PHN4016_U_afifo_U_acore_U_sub_fifo_n211), 
	.A(U_afifo_U_acore_U_sub_fifo_n211));
   BUF_X8 FE_PHC4015_U_afifo_U_acore_U_sub_fifo_n183 (.Z(FE_PHN4015_U_afifo_U_acore_U_sub_fifo_n183), 
	.A(U_afifo_U_acore_U_sub_fifo_n183));
   BUF_X8 FE_PHC4014_U_afifo_U_acore_U_sub_fifo_n207 (.Z(FE_PHN4014_U_afifo_U_acore_U_sub_fifo_n207), 
	.A(U_afifo_U_acore_U_sub_fifo_n207));
   BUF_X8 FE_PHC4011_U_afifo_U_acore_U_sub_fifo_n195 (.Z(FE_PHN4011_U_afifo_U_acore_U_sub_fifo_n195), 
	.A(U_afifo_U_acore_U_sub_fifo_n195));
   BUF_X8 FE_PHC4010_U_afifo_U_acore_U_sub_fifo_n182 (.Z(FE_PHN4010_U_afifo_U_acore_U_sub_fifo_n182), 
	.A(U_afifo_U_acore_U_sub_fifo_n182));
   BUF_X8 FE_PHC4009_U_afifo_U_acore_U_sub_fifo_n242 (.Z(FE_PHN4009_U_afifo_U_acore_U_sub_fifo_n242), 
	.A(U_afifo_U_acore_U_sub_fifo_n242));
   CLKBUF_X1 FE_PHC4008_U_dfifo_U_dcore_U_sub_fifo_n298 (.Z(FE_PHN4008_U_dfifo_U_dcore_U_sub_fifo_n298), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n298));
   BUF_X8 FE_PHC4007_U_dfifo_U_dcore_U_sub_fifo_n252 (.Z(FE_PHN4007_U_dfifo_U_dcore_U_sub_fifo_n252), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n252));
   BUF_X8 FE_PHC3999_U_afifo_U_acore_U_sub_fifo_n261 (.Z(FE_PHN3999_U_afifo_U_acore_U_sub_fifo_n261), 
	.A(U_afifo_U_acore_U_sub_fifo_n261));
   BUF_X8 FE_PHC3998_U_afifo_U_acore_U_sub_fifo_n174 (.Z(FE_PHN3998_U_afifo_U_acore_U_sub_fifo_n174), 
	.A(U_afifo_U_acore_U_sub_fifo_n174));
   BUF_X8 FE_PHC3997_U_afifo_U_acore_U_sub_fifo_n179 (.Z(FE_PHN3997_U_afifo_U_acore_U_sub_fifo_n179), 
	.A(U_afifo_U_acore_U_sub_fifo_n179));
   BUF_X8 FE_PHC3996_U_afifo_U_acore_U_sub_fifo_n204 (.Z(FE_PHN3996_U_afifo_U_acore_U_sub_fifo_n204), 
	.A(U_afifo_U_acore_U_sub_fifo_n204));
   BUF_X8 FE_PHC3995_U_afifo_U_acore_U_sub_fifo_n238 (.Z(FE_PHN3995_U_afifo_U_acore_U_sub_fifo_n238), 
	.A(U_afifo_U_acore_U_sub_fifo_n238));
   CLKBUF_X1 FE_PHC3994_U_afifo_U_acore_U_sub_fifo_n229 (.Z(FE_PHN3994_U_afifo_U_acore_U_sub_fifo_n229), 
	.A(U_afifo_U_acore_U_sub_fifo_n229));
   BUF_X8 FE_PHC3993_U_afifo_U_acore_U_sub_fifo_n254 (.Z(FE_PHN3993_U_afifo_U_acore_U_sub_fifo_n254), 
	.A(U_afifo_U_acore_U_sub_fifo_n254));
   CLKBUF_X1 FE_PHC3992_U_afifo_U_acore_U_sub_fifo_n240 (.Z(FE_PHN3992_U_afifo_U_acore_U_sub_fifo_n240), 
	.A(U_afifo_U_acore_U_sub_fifo_n240));
   BUF_X8 FE_PHC3991_U_afifo_U_acore_U_sub_fifo_n189 (.Z(FE_PHN3991_U_afifo_U_acore_U_sub_fifo_n189), 
	.A(U_afifo_U_acore_U_sub_fifo_n189));
   CLKBUF_X1 FE_PHC3990_U_afifo_U_acore_U_sub_fifo_n222 (.Z(FE_PHN3990_U_afifo_U_acore_U_sub_fifo_n222), 
	.A(U_afifo_U_acore_U_sub_fifo_n222));
   BUF_X8 FE_PHC3984_U_afifo_U_acore_U_sub_fifo_n216 (.Z(FE_PHN3984_U_afifo_U_acore_U_sub_fifo_n216), 
	.A(U_afifo_U_acore_U_sub_fifo_n216));
   BUF_X8 FE_PHC3980_U_afifo_U_acore_U_sub_fifo_n289 (.Z(FE_PHN3980_U_afifo_U_acore_U_sub_fifo_n289), 
	.A(U_afifo_U_acore_U_sub_fifo_n289));
   CLKBUF_X1 FE_PHC3979_U_afifo_U_acore_U_sub_fifo_n258 (.Z(FE_PHN3979_U_afifo_U_acore_U_sub_fifo_n258), 
	.A(U_afifo_U_acore_U_sub_fifo_n258));
   BUF_X8 FE_PHC3978_U_afifo_U_acore_U_sub_fifo_n244 (.Z(FE_PHN3978_U_afifo_U_acore_U_sub_fifo_n244), 
	.A(U_afifo_U_acore_U_sub_fifo_n244));
   BUF_X8 FE_PHC3967_U_afifo_U_acore_U_sub_fifo_n245 (.Z(FE_PHN3967_U_afifo_U_acore_U_sub_fifo_n245), 
	.A(U_afifo_U_acore_U_sub_fifo_n245));
   BUF_X8 FE_PHC3966_U_afifo_U_acore_U_sub_fifo_n228 (.Z(FE_PHN3966_U_afifo_U_acore_U_sub_fifo_n228), 
	.A(U_afifo_U_acore_U_sub_fifo_n228));
   BUF_X8 FE_PHC3965_U_dfifo_U_dcore_n152 (.Z(FE_PHN3965_U_dfifo_U_dcore_n152), 
	.A(U_dfifo_U_dcore_n152));
   CLKBUF_X1 FE_PHC3964_U_dfifo_U_dcore_U_sub_fifo_n205 (.Z(FE_PHN3964_U_dfifo_U_dcore_U_sub_fifo_n205), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n205));
   BUF_X8 FE_PHC3957_U_afifo_U_acore_U_sub_fifo_n186 (.Z(FE_PHN3957_U_afifo_U_acore_U_sub_fifo_n186), 
	.A(U_afifo_U_acore_U_sub_fifo_n186));
   BUF_X8 FE_PHC3956_U_afifo_U_acore_U_sub_fifo_n233 (.Z(FE_PHN3956_U_afifo_U_acore_U_sub_fifo_n233), 
	.A(U_afifo_U_acore_U_sub_fifo_n233));
   BUF_X8 FE_PHC3955_U_afifo_U_acore_U_sub_fifo_n281 (.Z(FE_PHN3955_U_afifo_U_acore_U_sub_fifo_n281), 
	.A(U_afifo_U_acore_U_sub_fifo_n281));
   BUF_X8 FE_PHC3953_U_afifo_U_acore_U_sub_fifo_n234 (.Z(FE_PHN3953_U_afifo_U_acore_U_sub_fifo_n234), 
	.A(U_afifo_U_acore_U_sub_fifo_n234));
   BUF_X8 FE_PHC3952_U_afifo_U_acore_U_sub_fifo_n286 (.Z(FE_PHN3952_U_afifo_U_acore_U_sub_fifo_n286), 
	.A(U_afifo_U_acore_U_sub_fifo_n286));
   BUF_X8 FE_PHC3947_U_afifo_U_acore_U_sub_fifo_n194 (.Z(FE_PHN3947_U_afifo_U_acore_U_sub_fifo_n194), 
	.A(U_afifo_U_acore_U_sub_fifo_n194));
   BUF_X8 FE_PHC3946_U_afifo_U_acore_U_sub_fifo_n282 (.Z(FE_PHN3946_U_afifo_U_acore_U_sub_fifo_n282), 
	.A(U_afifo_U_acore_U_sub_fifo_n282));
   BUF_X8 FE_PHC3945_U_afifo_U_acore_U_sub_fifo_n225 (.Z(FE_PHN3945_U_afifo_U_acore_U_sub_fifo_n225), 
	.A(U_afifo_U_acore_U_sub_fifo_n225));
   BUF_X8 FE_PHC3944_U_dfifo_U_dcore_U_sub_fifo_n171 (.Z(FE_PHN3944_U_dfifo_U_dcore_U_sub_fifo_n171), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n171));
   BUF_X8 FE_PHC3940_U_afifo_U_acore_U_sub_fifo_n239 (.Z(FE_PHN3940_U_afifo_U_acore_U_sub_fifo_n239), 
	.A(U_afifo_U_acore_U_sub_fifo_n239));
   BUF_X8 FE_PHC3939_U_afifo_U_acore_U_sub_fifo_n209 (.Z(FE_PHN3939_U_afifo_U_acore_U_sub_fifo_n209), 
	.A(U_afifo_U_acore_U_sub_fifo_n209));
   BUF_X8 FE_PHC3936_U_afifo_U_acore_U_sub_fifo_n231 (.Z(FE_PHN3936_U_afifo_U_acore_U_sub_fifo_n231), 
	.A(U_afifo_U_acore_U_sub_fifo_n231));
   BUF_X8 FE_PHC3935_U_afifo_U_acore_U_sub_fifo_n220 (.Z(FE_PHN3935_U_afifo_U_acore_U_sub_fifo_n220), 
	.A(U_afifo_U_acore_U_sub_fifo_n220));
   CLKBUF_X1 FE_PHC3933_U_dfifo_U_dcore_U_sub_fifo_n210 (.Z(FE_PHN3933_U_dfifo_U_dcore_U_sub_fifo_n210), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n210));
   CLKBUF_X1 FE_PHC3932_U_dfifo_U_dcore_U_sub_fifo_n170 (.Z(FE_PHN3932_U_dfifo_U_dcore_U_sub_fifo_n170), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n170));
   BUF_X8 FE_PHC3929_U_afifo_U_acore_U_sub_fifo_n241 (.Z(FE_PHN3929_U_afifo_U_acore_U_sub_fifo_n241), 
	.A(U_afifo_U_acore_U_sub_fifo_n241));
   BUF_X8 FE_PHC3920_U_afifo_U_acore_U_sub_fifo_n260 (.Z(FE_PHN3920_U_afifo_U_acore_U_sub_fifo_n260), 
	.A(U_afifo_U_acore_U_sub_fifo_n260));
   BUF_X8 FE_PHC3914_U_afifo_U_acore_U_sub_fifo_n217 (.Z(FE_PHN3914_U_afifo_U_acore_U_sub_fifo_n217), 
	.A(U_afifo_U_acore_U_sub_fifo_n217));
   CLKBUF_X1 FE_PHC3913_U_dfifo_U_dcore_U_sub_fifo_n164 (.Z(FE_PHN3913_U_dfifo_U_dcore_U_sub_fifo_n164), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n164));
   BUF_X8 FE_PHC3905_U_afifo_U_acore_U_sub_fifo_n237 (.Z(FE_PHN3905_U_afifo_U_acore_U_sub_fifo_n237), 
	.A(U_afifo_U_acore_U_sub_fifo_n237));
   BUF_X8 FE_PHC3901_U_afifo_U_acore_U_sub_fifo_n236 (.Z(FE_PHN3901_U_afifo_U_acore_U_sub_fifo_n236), 
	.A(U_afifo_U_acore_U_sub_fifo_n236));
   BUF_X8 FE_PHC3899_U_dfifo_U_dcore_U_sub_fifo_n213 (.Z(FE_PHN3899_U_dfifo_U_dcore_U_sub_fifo_n213), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n213));
   BUF_X8 FE_PHC3897_U_afifo_n158 (.Z(FE_PHN3897_U_afifo_n158), 
	.A(U_afifo_n158));
   BUF_X8 FE_PHC3895_U_afifo_U_acore_U_sub_fifo_n235 (.Z(FE_PHN3895_U_afifo_U_acore_U_sub_fifo_n235), 
	.A(U_afifo_U_acore_U_sub_fifo_n235));
   BUF_X8 FE_PHC3894_U_dfifo_U_dcore_U_sub_fifo_n216 (.Z(FE_PHN3894_U_dfifo_U_dcore_U_sub_fifo_n216), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n216));
   BUF_X8 FE_PHC3891_U_afifo_U_acore_U_sub_fifo_n185 (.Z(FE_PHN3891_U_afifo_U_acore_U_sub_fifo_n185), 
	.A(U_afifo_U_acore_U_sub_fifo_n185));
   BUF_X8 FE_PHC3890_U_afifo_U_acore_U_sub_fifo_n255 (.Z(FE_PHN3890_U_afifo_U_acore_U_sub_fifo_n255), 
	.A(U_afifo_U_acore_U_sub_fifo_n255));
   BUF_X8 FE_PHC3881_U_afifo_U_acore_U_sub_fifo_n246 (.Z(FE_PHN3881_U_afifo_U_acore_U_sub_fifo_n246), 
	.A(U_afifo_U_acore_U_sub_fifo_n246));
   BUF_X8 FE_PHC3873_U_dfifo_U_dcore_n151 (.Z(FE_PHN3873_U_dfifo_U_dcore_n151), 
	.A(U_dfifo_U_dcore_n151));
   BUF_X8 FE_PHC3861_U_dfifo_U_dcore_U_sub_fifo_n214 (.Z(FE_PHN3861_U_dfifo_U_dcore_U_sub_fifo_n214), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n214));
   BUF_X8 FE_PHC3860_U_dfifo_U_dcore_U_sub_fifo_n218 (.Z(FE_PHN3860_U_dfifo_U_dcore_U_sub_fifo_n218), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n218));
   BUF_X8 FE_PHC3859_U_dfifo_U_dcore_U_sub_fifo_n163 (.Z(FE_PHN3859_U_dfifo_U_dcore_U_sub_fifo_n163), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n163));
   BUF_X8 FE_PHC3858_U_dfifo_U_dcore_U_sub_fifo_n209 (.Z(FE_PHN3858_U_dfifo_U_dcore_U_sub_fifo_n209), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n209));
   BUF_X8 FE_PHC3855_U_dfifo_U_dcore_U_sub_fifo_n215 (.Z(FE_PHN3855_U_dfifo_U_dcore_U_sub_fifo_n215), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n215));
   BUF_X8 FE_PHC3854_U_dfifo_U_dcore_U_sub_fifo_n219 (.Z(FE_PHN3854_U_dfifo_U_dcore_U_sub_fifo_n219), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n219));
   BUF_X8 FE_PHC3852_U_dfifo_U_dcore_U_sub_fifo_n202 (.Z(FE_PHN3852_U_dfifo_U_dcore_U_sub_fifo_n202), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n202));
   BUF_X8 FE_PHC3850_U_dfifo_U_dcore_U_sub_fifo_n178 (.Z(FE_PHN3850_U_dfifo_U_dcore_U_sub_fifo_n178), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n178));
   BUF_X8 FE_PHC3849_U_dfifo_U_dcore_U_sub_fifo_n175 (.Z(FE_PHN3849_U_dfifo_U_dcore_U_sub_fifo_n175), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n175));
   BUF_X8 FE_PHC3848_U_dfifo_U_dcore_U_sub_fifo_n166 (.Z(FE_PHN3848_U_dfifo_U_dcore_U_sub_fifo_n166), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n166));
   BUF_X8 FE_PHC3846_U_dfifo_U_dcore_U_sub_fifo_n211 (.Z(FE_PHN3846_U_dfifo_U_dcore_U_sub_fifo_n211), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n211));
   BUF_X8 FE_PHC3841_U_dfifo_U_dcore_U_sub_fifo_n207 (.Z(FE_PHN3841_U_dfifo_U_dcore_U_sub_fifo_n207), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n207));
   BUF_X8 FE_PHC3840_U_dfifo_U_dcore_U_sub_fifo_n314 (.Z(FE_PHN3840_U_dfifo_U_dcore_U_sub_fifo_n314), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n314));
   BUF_X16 FE_PHC3838_U_dfifo_U_dcore_U_sub_fifo_n177 (.Z(FE_PHN3838_U_dfifo_U_dcore_U_sub_fifo_n177), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n177));
   BUF_X16 FE_PHC3837_U_afifo_U_acore_U_sub_fifo_n268 (.Z(FE_PHN3837_U_afifo_U_acore_U_sub_fifo_n268), 
	.A(U_afifo_U_acore_U_sub_fifo_n268));
   BUF_X8 FE_PHC3835_U_dfifo_U_dcore_U_sub_fifo_n169 (.Z(FE_PHN3835_U_dfifo_U_dcore_U_sub_fifo_n169), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n169));
   CLKBUF_X1 FE_PHC3834_U_dfifo_U_dcore_U_sub_fifo_n206 (.Z(FE_PHN3834_U_dfifo_U_dcore_U_sub_fifo_n206), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n206));
   BUF_X8 FE_PHC3832_U_dfifo_U_dcore_U_sub_fifo_n174 (.Z(FE_PHN3832_U_dfifo_U_dcore_U_sub_fifo_n174), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n174));
   BUF_X16 FE_PHC3829_U_dfifo_U_dcore_U_sub_fifo_n337 (.Z(FE_PHN3829_U_dfifo_U_dcore_U_sub_fifo_n337), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n337));
   BUF_X16 FE_PHC3827_U_dfifo_U_dcore_U_sub_fifo_n162 (.Z(FE_PHN3827_U_dfifo_U_dcore_U_sub_fifo_n162), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n162));
   BUF_X8 FE_PHC3825_U_dfifo_U_dcore_U_sub_fifo_n445 (.Z(FE_PHN3825_U_dfifo_U_dcore_U_sub_fifo_n445), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n445));
   BUF_X8 FE_PHC3824_U_dfifo_U_dcore_U_sub_fifo_n168 (.Z(FE_PHN3824_U_dfifo_U_dcore_U_sub_fifo_n168), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n168));
   BUF_X8 FE_PHC3822_U_dfifo_U_dcore_U_sub_fifo_n413 (.Z(FE_PHN3822_U_dfifo_U_dcore_U_sub_fifo_n413), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n413));
   BUF_X8 FE_PHC3820_U_dfifo_U_dcore_U_sub_fifo_n220 (.Z(FE_PHN3820_U_dfifo_U_dcore_U_sub_fifo_n220), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n220));
   BUF_X8 FE_PHC3819_U_dfifo_U_dcore_U_sub_fifo_n165 (.Z(FE_PHN3819_U_dfifo_U_dcore_U_sub_fifo_n165), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n165));
   BUF_X8 FE_PHC3818_U_dfifo_U_dcore_U_sub_fifo_n173 (.Z(FE_PHN3818_U_dfifo_U_dcore_U_sub_fifo_n173), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n173));
   BUF_X8 FE_PHC3817_U_afifo_U_acore_U_sub_fifo_n267 (.Z(FE_PHN3817_U_afifo_U_acore_U_sub_fifo_n267), 
	.A(U_afifo_U_acore_U_sub_fifo_n267));
   BUF_X8 FE_PHC3815_U_dfifo_U_dcore_U_sub_fifo_n212 (.Z(FE_PHN3815_U_dfifo_U_dcore_U_sub_fifo_n212), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n212));
   BUF_X16 FE_PHC3813_U_afifo_U_acore_U_sub_fifo_n272 (.Z(FE_PHN3813_U_afifo_U_acore_U_sub_fifo_n272), 
	.A(U_afifo_U_acore_U_sub_fifo_n272));
   BUF_X8 FE_PHC3812_U_dfifo_U_dcore_U_sub_fifo_n176 (.Z(FE_PHN3812_U_dfifo_U_dcore_U_sub_fifo_n176), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n176));
   BUF_X16 FE_PHC3809_U_dfifo_U_dcore_U_sub_fifo_n329 (.Z(FE_PHN3809_U_dfifo_U_dcore_U_sub_fifo_n329), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n329));
   BUF_X8 FE_PHC3807_U_dfifo_U_dcore_U_sub_fifo_n172 (.Z(FE_PHN3807_U_dfifo_U_dcore_U_sub_fifo_n172), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n172));
   BUF_X8 FE_PHC3805_U_dfifo_U_dcore_U_sub_fifo_n204 (.Z(FE_PHN3805_U_dfifo_U_dcore_U_sub_fifo_n204), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n204));
   BUF_X16 FE_PHC3804_U_dfifo_U_dcore_U_sub_fifo_n330 (.Z(FE_PHN3804_U_dfifo_U_dcore_U_sub_fifo_n330), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n330));
   BUF_X16 FE_PHC3801_U_dfifo_U_dcore_U_sub_fifo_n415 (.Z(FE_PHN3801_U_dfifo_U_dcore_U_sub_fifo_n415), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n415));
   BUF_X8 FE_PHC3795_U_afifo_U_acore_U_sub_fifo_n266 (.Z(FE_PHN3795_U_afifo_U_acore_U_sub_fifo_n266), 
	.A(U_afifo_U_acore_U_sub_fifo_n266));
   BUF_X16 FE_PHC3794_U_dfifo_U_dcore_U_sub_fifo_n321 (.Z(FE_PHN3794_U_dfifo_U_dcore_U_sub_fifo_n321), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n321));
   BUF_X16 FE_PHC3792_U_dfifo_U_dcore_U_sub_fifo_n217 (.Z(FE_PHN3792_U_dfifo_U_dcore_U_sub_fifo_n217), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n217));
   BUF_X8 FE_PHC3791_U_dfifo_U_dcore_U_sub_fifo_n401 (.Z(FE_PHN3791_U_dfifo_U_dcore_U_sub_fifo_n401), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n401));
   BUF_X8 FE_PHC3790_U_dfifo_U_dcore_U_sub_fifo_n338 (.Z(FE_PHN3790_U_dfifo_U_dcore_U_sub_fifo_n338), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n338));
   BUF_X16 FE_PHC3789_U_dfifo_U_dcore_n144 (.Z(FE_PHN3789_U_dfifo_U_dcore_n144), 
	.A(U_dfifo_U_dcore_n144));
   BUF_X16 FE_PHC3788_U_dfifo_U_dcore_U_sub_fifo_n317 (.Z(FE_PHN3788_U_dfifo_U_dcore_U_sub_fifo_n317), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n317));
   BUF_X8 FE_PHC3783_U_dfifo_U_dcore_U_sub_fifo_n333 (.Z(FE_PHN3783_U_dfifo_U_dcore_U_sub_fifo_n333), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n333));
   BUF_X16 FE_PHC3772_U_afifo_U_acore_U_sub_fifo_n270 (.Z(FE_PHN3772_U_afifo_U_acore_U_sub_fifo_n270), 
	.A(U_afifo_U_acore_U_sub_fifo_n270));
   BUF_X16 FE_PHC3770_U_afifo_n20 (.Z(FE_PHN3770_U_afifo_n20), 
	.A(U_afifo_n20));
   BUF_X8 FE_PHC3767_U_dfifo_U_dcore_U_sub_fifo_n344 (.Z(FE_PHN3767_U_dfifo_U_dcore_U_sub_fifo_n344), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n344));
   BUF_X16 FE_PHC3761_U_dfifo_U_dcore_U_sub_fifo_n203 (.Z(FE_PHN3761_U_dfifo_U_dcore_U_sub_fifo_n203), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n203));
   BUF_X16 FE_PHC3756_U_dfifo_U_dcore_n143 (.Z(FE_PHN3756_U_dfifo_U_dcore_n143), 
	.A(U_dfifo_U_dcore_n143));
   BUF_X16 FE_PHC3754_U_dfifo_U_dcore_U_sub_fifo_n315 (.Z(FE_PHN3754_U_dfifo_U_dcore_U_sub_fifo_n315), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n315));
   BUF_X16 FE_PHC3752_U_dfifo_U_dcore_U_sub_fifo_n416 (.Z(FE_PHN3752_U_dfifo_U_dcore_U_sub_fifo_n416), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n416));
   BUF_X16 FE_PHC3750_U_dfifo_U_dcore_U_sub_fifo_n407 (.Z(FE_PHN3750_U_dfifo_U_dcore_U_sub_fifo_n407), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n407));
   BUF_X8 FE_PHC3749_U_dfifo_U_dcore_U_sub_fifo_n167 (.Z(FE_PHN3749_U_dfifo_U_dcore_U_sub_fifo_n167), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n167));
   BUF_X16 FE_PHC3748_U_dfifo_U_dcore_U_sub_fifo_n313 (.Z(FE_PHN3748_U_dfifo_U_dcore_U_sub_fifo_n313), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n313));
   BUF_X8 FE_PHC3747_U_dfifo_U_dcore_U_sub_fifo_n403 (.Z(FE_PHN3747_U_dfifo_U_dcore_U_sub_fifo_n403), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n403));
   BUF_X8 FE_PHC3746_U_dfifo_U_dcore_U_sub_fifo_n397 (.Z(FE_PHN3746_U_dfifo_U_dcore_U_sub_fifo_n397), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n397));
   BUF_X16 FE_PHC3743_U_dfifo_U_dcore_U_sub_fifo_n417 (.Z(FE_PHN3743_U_dfifo_U_dcore_U_sub_fifo_n417), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n417));
   BUF_X16 FE_PHC3742_U_dfifo_U_dcore_U_sub_fifo_n324 (.Z(FE_PHN3742_U_dfifo_U_dcore_U_sub_fifo_n324), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n324));
   BUF_X16 FE_PHC3741_U_dfifo_U_dcore_U_sub_fifo_n325 (.Z(FE_PHN3741_U_dfifo_U_dcore_U_sub_fifo_n325), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n325));
   BUF_X8 FE_PHC3740_U_dfifo_U_dcore_U_sub_fifo_n398 (.Z(FE_PHN3740_U_dfifo_U_dcore_U_sub_fifo_n398), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n398));
   BUF_X8 FE_PHC3734_U_dfifo_U_dcore_U_sub_fifo_n208 (.Z(FE_PHN3734_U_dfifo_U_dcore_U_sub_fifo_n208), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n208));
   BUF_X16 FE_PHC3732_U_dfifo_U_dcore_U_sub_fifo_n326 (.Z(FE_PHN3732_U_dfifo_U_dcore_U_sub_fifo_n326), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n326));
   BUF_X8 FE_PHC3731_U_dfifo_U_dcore_U_sub_fifo_n442 (.Z(FE_PHN3731_U_dfifo_U_dcore_U_sub_fifo_n442), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n442));
   BUF_X8 FE_PHC3729_U_dfifo_U_dcore_U_sub_fifo_n356 (.Z(FE_PHN3729_U_dfifo_U_dcore_U_sub_fifo_n356), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n356));
   BUF_X16 FE_PHC3728_U_dfifo_U_dcore_U_sub_fifo_n318 (.Z(FE_PHN3728_U_dfifo_U_dcore_U_sub_fifo_n318), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n318));
   BUF_X16 FE_PHC3727_U_dfifo_U_dcore_U_sub_fifo_n443 (.Z(FE_PHN3727_U_dfifo_U_dcore_U_sub_fifo_n443), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n443));
   BUF_X8 FE_PHC3723_U_dfifo_U_dcore_U_sub_fifo_n340 (.Z(FE_PHN3723_U_dfifo_U_dcore_U_sub_fifo_n340), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n340));
   BUF_X16 FE_PHC3721_U_dfifo_U_dcore_U_sub_fifo_n411 (.Z(FE_PHN3721_U_dfifo_U_dcore_U_sub_fifo_n411), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n411));
   BUF_X8 FE_PHC3720_U_dfifo_U_dcore_U_sub_fifo_n402 (.Z(FE_PHN3720_U_dfifo_U_dcore_U_sub_fifo_n402), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n402));
   BUF_X8 FE_PHC3719_U_dfifo_U_dcore_U_sub_fifo_n440 (.Z(FE_PHN3719_U_dfifo_U_dcore_U_sub_fifo_n440), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n440));
   BUF_X16 FE_PHC3716_U_dfifo_U_dcore_n147 (.Z(FE_PHN3716_U_dfifo_U_dcore_n147), 
	.A(U_dfifo_U_dcore_n147));
   BUF_X16 FE_PHC3715_U_dfifo_U_dcore_U_sub_fifo_n127 (.Z(FE_PHN3715_U_dfifo_U_dcore_U_sub_fifo_n127), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n127));
   BUF_X16 FE_PHC3711_U_dfifo_U_dcore_U_sub_fifo_n405 (.Z(FE_PHN3711_U_dfifo_U_dcore_U_sub_fifo_n405), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n405));
   BUF_X16 FE_PHC3710_U_dfifo_U_dcore_U_sub_fifo_n406 (.Z(FE_PHN3710_U_dfifo_U_dcore_U_sub_fifo_n406), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n406));
   BUF_X8 FE_PHC3709_U_dfifo_U_dcore_U_sub_fifo_n412 (.Z(FE_PHN3709_U_dfifo_U_dcore_U_sub_fifo_n412), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n412));
   BUF_X8 FE_PHC3708_U_dfifo_U_dcore_U_sub_fifo_n327 (.Z(FE_PHN3708_U_dfifo_U_dcore_U_sub_fifo_n327), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n327));
   BUF_X16 FE_PHC3706_U_dfifo_U_dcore_U_sub_fifo_n399 (.Z(FE_PHN3706_U_dfifo_U_dcore_U_sub_fifo_n399), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n399));
   BUF_X16 FE_PHC3705_U_dfifo_U_dcore_U_sub_fifo_n339 (.Z(FE_PHN3705_U_dfifo_U_dcore_U_sub_fifo_n339), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n339));
   BUF_X16 FE_PHC3703_U_dfifo_U_dcore_U_sub_fifo_n414 (.Z(FE_PHN3703_U_dfifo_U_dcore_U_sub_fifo_n414), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n414));
   BUF_X16 FE_PHC3701_U_dfifo_U_dcore_U_sub_fifo_n400 (.Z(FE_PHN3701_U_dfifo_U_dcore_U_sub_fifo_n400), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n400));
   BUF_X8 FE_PHC3700_U_dfifo_U_dcore_U_sub_fifo_n320 (.Z(FE_PHN3700_U_dfifo_U_dcore_U_sub_fifo_n320), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n320));
   BUF_X16 FE_PHC3696_U_dfifo_U_dcore_U_sub_fifo_n323 (.Z(FE_PHN3696_U_dfifo_U_dcore_U_sub_fifo_n323), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n323));
   BUF_X16 FE_PHC3695_U_dfifo_U_dcore_U_sub_fifo_n311 (.Z(FE_PHN3695_U_dfifo_U_dcore_U_sub_fifo_n311), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n311));
   BUF_X16 FE_PHC3694_U_dfifo_U_dcore_U_sub_fifo_n404 (.Z(FE_PHN3694_U_dfifo_U_dcore_U_sub_fifo_n404), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n404));
   BUF_X16 FE_PHC3693_U_dfifo_U_dcore_U_sub_fifo_n331 (.Z(FE_PHN3693_U_dfifo_U_dcore_U_sub_fifo_n331), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n331));
   BUF_X16 FE_PHC3691_U_dfifo_U_dcore_U_sub_fifo_n334 (.Z(FE_PHN3691_U_dfifo_U_dcore_U_sub_fifo_n334), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n334));
   BUF_X16 FE_PHC3689_U_dfifo_U_dcore_U_sub_fifo_n441 (.Z(FE_PHN3689_U_dfifo_U_dcore_U_sub_fifo_n441), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n441));
   BUF_X16 FE_PHC3688_U_dfifo_U_dcore_U_sub_fifo_n439 (.Z(FE_PHN3688_U_dfifo_U_dcore_U_sub_fifo_n439), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n439));
   BUF_X16 FE_PHC3685_U_dfifo_U_dcore_U_sub_fifo_n418 (.Z(FE_PHN3685_U_dfifo_U_dcore_U_sub_fifo_n418), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n418));
   BUF_X16 FE_PHC3679_U_dfifo_U_dcore_U_sub_fifo_n343 (.Z(FE_PHN3679_U_dfifo_U_dcore_U_sub_fifo_n343), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n343));
   BUF_X16 FE_PHC3678_U_dfifo_U_dcore_U_sub_fifo_n319 (.Z(FE_PHN3678_U_dfifo_U_dcore_U_sub_fifo_n319), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n319));
   BUF_X16 FE_PHC3677_U_dfifo_U_dcore_U_sub_fifo_n332 (.Z(FE_PHN3677_U_dfifo_U_dcore_U_sub_fifo_n332), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n332));
   BUF_X16 FE_PHC3676_U_dfifo_U_dcore_U_sub_fifo_n444 (.Z(FE_PHN3676_U_dfifo_U_dcore_U_sub_fifo_n444), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n444));
   BUF_X16 FE_PHC3675_U_dfifo_U_dcore_U_sub_fifo_n438 (.Z(FE_PHN3675_U_dfifo_U_dcore_U_sub_fifo_n438), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n438));
   BUF_X16 FE_PHC3674_U_dfifo_U_dcore_U_sub_fifo_n322 (.Z(FE_PHN3674_U_dfifo_U_dcore_U_sub_fifo_n322), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n322));
   BUF_X8 FE_PHC3673_U_dfifo_U_dcore_U_sub_fifo_n446 (.Z(FE_PHN3673_U_dfifo_U_dcore_U_sub_fifo_n446), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n446));
   BUF_X16 FE_PHC3671_U_afifo_n18 (.Z(FE_PHN3671_U_afifo_n18), 
	.A(U_afifo_n18));
   BUF_X16 FE_PHC3670_U_dfifo_U_dcore_U_sub_fifo_n328 (.Z(FE_PHN3670_U_dfifo_U_dcore_U_sub_fifo_n328), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n328));
   BUF_X16 FE_PHC3668_U_dfifo_U_dcore_U_sub_fifo_n341 (.Z(FE_PHN3668_U_dfifo_U_dcore_U_sub_fifo_n341), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n341));
   BUF_X16 FE_PHC3667_U_dfifo_U_dcore_U_sub_fifo_n408 (.Z(FE_PHN3667_U_dfifo_U_dcore_U_sub_fifo_n408), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n408));
   BUF_X16 FE_PHC3664_U_dfifo_U_dcore_U_sub_fifo_n410 (.Z(FE_PHN3664_U_dfifo_U_dcore_U_sub_fifo_n410), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n410));
   BUF_X16 FE_PHC3658_U_dfifo_U_dcore_U_sub_fifo_n409 (.Z(FE_PHN3658_U_dfifo_U_dcore_U_sub_fifo_n409), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n409));
   BUF_X16 FE_PHC3656_U_dfifo_U_dcore_U_sub_fifo_n335 (.Z(FE_PHN3656_U_dfifo_U_dcore_U_sub_fifo_n335), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n335));
   BUF_X16 FE_PHC3655_U_dfifo_U_dcore_n146 (.Z(FE_PHN3655_U_dfifo_U_dcore_n146), 
	.A(U_dfifo_U_dcore_n146));
   BUF_X16 FE_PHC3652_U_dfifo_U_dcore_U_sub_fifo_n312 (.Z(FE_PHN3652_U_dfifo_U_dcore_U_sub_fifo_n312), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n312));
   BUF_X16 FE_PHC3650_U_dfifo_U_dcore_U_sub_fifo_n342 (.Z(FE_PHN3650_U_dfifo_U_dcore_U_sub_fifo_n342), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n342));
   BUF_X16 FE_PHC3649_U_dfifo_U_dcore_U_sub_fifo_n336 (.Z(FE_PHN3649_U_dfifo_U_dcore_U_sub_fifo_n336), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n336));
   BUF_X16 FE_PHC3646_U_afifo_n19 (.Z(FE_PHN3646_U_afifo_n19), 
	.A(U_afifo_n19));
   BUF_X8 FE_PHC3644_U_dfifo_U_dcore_U_sub_fifo_n316 (.Z(FE_PHN3644_U_dfifo_U_dcore_U_sub_fifo_n316), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n316));
   BUF_X16 FE_PHC3632_U_dfifo_U_dcore_n13 (.Z(FE_PHN3632_U_dfifo_U_dcore_n13), 
	.A(U_dfifo_U_dcore_n13));
   BUF_X16 FE_PHC3618_U_dfifo_U_dcore_n14 (.Z(FE_PHN3618_U_dfifo_U_dcore_n14), 
	.A(U_dfifo_U_dcore_n14));
   BUF_X32 FE_PHC3543_U_afifo_n164 (.Z(FE_PHN3543_U_afifo_n164), 
	.A(U_afifo_n164));
   CLKBUF_X1 FE_PHC3504_U_afifo_U_acore_U_sub_fifo_n223 (.Z(FE_PHN3504_U_afifo_U_acore_U_sub_fifo_n223), 
	.A(U_afifo_U_acore_U_sub_fifo_n223));
   CLKBUF_X1 FE_PHC3499_U_afifo_U_acore_U_sub_fifo_n248 (.Z(FE_PHN3499_U_afifo_U_acore_U_sub_fifo_n248), 
	.A(U_afifo_U_acore_U_sub_fifo_n248));
   CLKBUF_X1 FE_PHC3498_U_afifo_U_acore_U_sub_fifo_n250 (.Z(FE_PHN3498_U_afifo_U_acore_U_sub_fifo_n250), 
	.A(U_afifo_U_acore_U_sub_fifo_n250));
   CLKBUF_X1 FE_PHC3495_U_afifo_U_acore_U_sub_fifo_n173 (.Z(FE_PHN3495_U_afifo_U_acore_U_sub_fifo_n173), 
	.A(U_afifo_U_acore_U_sub_fifo_n173));
   BUF_X8 FE_PHC3494_U_afifo_U_acore_U_sub_fifo_n219 (.Z(FE_PHN3494_U_afifo_U_acore_U_sub_fifo_n219), 
	.A(U_afifo_U_acore_U_sub_fifo_n219));
   BUF_X8 FE_PHC3493_U_afifo_U_acore_U_sub_fifo_n253 (.Z(FE_PHN3493_U_afifo_U_acore_U_sub_fifo_n253), 
	.A(U_afifo_U_acore_U_sub_fifo_n253));
   BUF_X8 FE_PHC3492_U_afifo_U_acore_U_sub_fifo_n226 (.Z(FE_PHN3492_U_afifo_U_acore_U_sub_fifo_n226), 
	.A(U_afifo_U_acore_U_sub_fifo_n226));
   CLKBUF_X1 FE_PHC3491_U_afifo_U_acore_U_sub_fifo_n177 (.Z(FE_PHN3491_U_afifo_U_acore_U_sub_fifo_n177), 
	.A(U_afifo_U_acore_U_sub_fifo_n177));
   BUF_X1 FE_PHC3490_U_afifo_U_acore_U_sub_fifo_n227 (.Z(FE_PHN3490_U_afifo_U_acore_U_sub_fifo_n227), 
	.A(U_afifo_U_acore_U_sub_fifo_n227));
   CLKBUF_X1 FE_PHC3489_U_afifo_U_acore_U_sub_fifo_n256 (.Z(FE_PHN3489_U_afifo_U_acore_U_sub_fifo_n256), 
	.A(U_afifo_U_acore_U_sub_fifo_n256));
   BUF_X8 FE_PHC3488_U_afifo_U_acore_U_sub_fifo_n252 (.Z(FE_PHN3488_U_afifo_U_acore_U_sub_fifo_n252), 
	.A(U_afifo_U_acore_U_sub_fifo_n252));
   BUF_X8 FE_PHC3487_U_afifo_U_acore_U_sub_fifo_n199 (.Z(FE_PHN3487_U_afifo_U_acore_U_sub_fifo_n199), 
	.A(U_afifo_U_acore_U_sub_fifo_n199));
   BUF_X8 FE_PHC3486_U_afifo_U_acore_U_sub_fifo_n193 (.Z(FE_PHN3486_U_afifo_U_acore_U_sub_fifo_n193), 
	.A(U_afifo_U_acore_U_sub_fifo_n193));
   BUF_X8 FE_PHC3484_U_afifo_U_acore_U_sub_fifo_n251 (.Z(FE_PHN3484_U_afifo_U_acore_U_sub_fifo_n251), 
	.A(U_afifo_U_acore_U_sub_fifo_n251));
   BUF_X8 FE_PHC3483_U_afifo_U_acore_U_sub_fifo_n243 (.Z(FE_PHN3483_U_afifo_U_acore_U_sub_fifo_n243), 
	.A(U_afifo_U_acore_U_sub_fifo_n243));
   BUF_X16 FE_PHC3481_U_afifo_n157 (.Z(FE_PHN3481_U_afifo_n157), 
	.A(U_afifo_n157));
   BUF_X32 FE_PHC3471_U_afifo_m_data_in_49_ (.Z(FE_PHN3471_U_afifo_m_data_in_49_), 
	.A(U_afifo_m_data_in[49]));
   BUF_X32 FE_PHC3469_U_ctl_n136 (.Z(FE_PHN3469_U_ctl_n136), 
	.A(U_ctl_n136));
   CLKBUF_X1 FE_PHC3468_U_ctl_n103 (.Z(FE_PHN3468_U_ctl_n103), 
	.A(FE_PHN1102_U_ctl_n103));
   CLKBUF_X2 FE_PHC3465_U_afifo_U_acore_f_obuf_34_ (.Z(FE_PHN3465_U_afifo_U_acore_f_obuf_34_), 
	.A(U_afifo_U_acore_f_obuf_34_));
   BUF_X1 FE_PHC3462_U_ctl_n101 (.Z(FE_PHN3462_U_ctl_n101), 
	.A(FE_PHN1342_U_ctl_n101));
   CLKBUF_X1 FE_PHC3460_U_afifo_U_acore_n157 (.Z(FE_PHN3460_U_afifo_U_acore_n157), 
	.A(U_afifo_U_acore_n157));
   CLKBUF_X1 FE_PHC3459_U_afifo_U_acore_n91 (.Z(FE_PHN3459_U_afifo_U_acore_n91), 
	.A(U_afifo_U_acore_n91));
   BUF_X1 FE_PHC3458_U_afifo_n186 (.Z(FE_PHN3458_U_afifo_n186), 
	.A(U_afifo_n186));
   CLKBUF_X1 FE_PHC3457_U_afifo_U_acore_n69 (.Z(FE_PHN3457_U_afifo_U_acore_n69), 
	.A(U_afifo_U_acore_n69));
   CLKBUF_X1 FE_PHC3455_U_afifo_U_acore_n164 (.Z(FE_PHN3455_U_afifo_U_acore_n164), 
	.A(U_afifo_U_acore_n164));
   CLKBUF_X1 FE_PHC3453_U_afifo_U_acore_n75 (.Z(FE_PHN3453_U_afifo_U_acore_n75), 
	.A(U_afifo_U_acore_n75));
   CLKBUF_X1 FE_PHC3451_U_ctl_n102 (.Z(FE_PHN3451_U_ctl_n102), 
	.A(FE_PHN1226_U_ctl_n102));
   CLKBUF_X1 FE_PHC3448_U_afifo_U_acore_n89 (.Z(FE_PHN3448_U_afifo_U_acore_n89), 
	.A(U_afifo_U_acore_n89));
   CLKBUF_X1 FE_PHC3447_U_afifo_U_acore_n101 (.Z(FE_PHN3447_U_afifo_U_acore_n101), 
	.A(U_afifo_U_acore_n101));
   CLKBUF_X1 FE_PHC3444_U_afifo_U_acore_n87 (.Z(FE_PHN3444_U_afifo_U_acore_n87), 
	.A(U_afifo_U_acore_n87));
   CLKBUF_X1 FE_PHC3441_U_afifo_n202 (.Z(FE_PHN3441_U_afifo_n202), 
	.A(U_afifo_n202));
   CLKBUF_X1 FE_PHC3439_U_afifo_n212 (.Z(FE_PHN3439_U_afifo_n212), 
	.A(U_afifo_n212));
   CLKBUF_X1 FE_PHC3438_U_dfifo_U_dcore_n200 (.Z(FE_PHN3438_U_dfifo_U_dcore_n200), 
	.A(U_dfifo_U_dcore_n200));
   CLKBUF_X1 FE_PHC3436_U_afifo_n208 (.Z(FE_PHN3436_U_afifo_n208), 
	.A(U_afifo_n208));
   CLKBUF_X1 FE_PHC3435_U_afifo_n198 (.Z(FE_PHN3435_U_afifo_n198), 
	.A(U_afifo_n198));
   CLKBUF_X1 FE_PHC3434_U_afifo_n210 (.Z(FE_PHN3434_U_afifo_n210), 
	.A(U_afifo_n210));
   CLKBUF_X1 FE_PHC3433_U_afifo_U_acore_n155 (.Z(FE_PHN3433_U_afifo_U_acore_n155), 
	.A(U_afifo_U_acore_n155));
   CLKBUF_X1 FE_PHC3430_U_afifo_U_acore_n143 (.Z(FE_PHN3430_U_afifo_U_acore_n143), 
	.A(U_afifo_U_acore_n143));
   CLKBUF_X1 FE_PHC3429_U_afifo_n220 (.Z(FE_PHN3429_U_afifo_n220), 
	.A(U_afifo_n220));
   CLKBUF_X1 FE_PHC3428_U_dfifo_U_dcore_n140 (.Z(FE_PHN3428_U_dfifo_U_dcore_n140), 
	.A(U_dfifo_U_dcore_n140));
   CLKBUF_X1 FE_PHC3426_U_afifo_U_acore_n_obuf_empty (.Z(FE_PHN3426_U_afifo_U_acore_n_obuf_empty), 
	.A(FE_PHN750_U_afifo_U_acore_n_obuf_empty));
   CLKBUF_X1 FE_PHC3425_U_afifo_n188 (.Z(FE_PHN3425_U_afifo_n188), 
	.A(U_afifo_n188));
   CLKBUF_X1 FE_PHC3424_U_afifo_n232 (.Z(FE_PHN3424_U_afifo_n232), 
	.A(U_afifo_n232));
   CLKBUF_X1 FE_PHC3423_U_afifo_U_acore_n29 (.Z(FE_PHN3423_U_afifo_U_acore_n29), 
	.A(U_afifo_U_acore_n29));
   CLKBUF_X1 FE_PHC3422_U_afifo_n226 (.Z(FE_PHN3422_U_afifo_n226), 
	.A(U_afifo_n226));
   CLKBUF_X1 FE_PHC3420_U_afifo_n206 (.Z(FE_PHN3420_U_afifo_n206), 
	.A(U_afifo_n206));
   CLKBUF_X1 FE_PHC3419_U_afifo_n248 (.Z(FE_PHN3419_U_afifo_n248), 
	.A(U_afifo_n248));
   CLKBUF_X1 FE_PHC3418_U_afifo_n236 (.Z(FE_PHN3418_U_afifo_n236), 
	.A(U_afifo_n236));
   CLKBUF_X1 FE_PHC3417_U_dfifo_U_dcore_n194 (.Z(FE_PHN3417_U_dfifo_U_dcore_n194), 
	.A(U_dfifo_U_dcore_n194));
   CLKBUF_X1 FE_PHC3416_U_afifo_U_acore_n67 (.Z(FE_PHN3416_U_afifo_U_acore_n67), 
	.A(U_afifo_U_acore_n67));
   CLKBUF_X1 FE_PHC3413_U_afifo_n204 (.Z(FE_PHN3413_U_afifo_n204), 
	.A(U_afifo_n204));
   CLKBUF_X1 FE_PHC3412_U_afifo_U_acore_n158 (.Z(FE_PHN3412_U_afifo_U_acore_n158), 
	.A(U_afifo_U_acore_n158));
   CLKBUF_X1 FE_PHC3410_U_afifo_n230 (.Z(FE_PHN3410_U_afifo_n230), 
	.A(U_afifo_n230));
   CLKBUF_X1 FE_PHC3409_U_afifo_U_acore_n153 (.Z(FE_PHN3409_U_afifo_U_acore_n153), 
	.A(U_afifo_U_acore_n153));
   CLKBUF_X1 FE_PHC3408_U_afifo_n234 (.Z(FE_PHN3408_U_afifo_n234), 
	.A(U_afifo_n234));
   CLKBUF_X1 FE_PHC3406_U_afifo_U_acore_n99 (.Z(FE_PHN3406_U_afifo_U_acore_n99), 
	.A(U_afifo_U_acore_n99));
   CLKBUF_X1 FE_PHC3404_U_afifo_n218 (.Z(FE_PHN3404_U_afifo_n218), 
	.A(U_afifo_n218));
   CLKBUF_X1 FE_PHC3403_U_afifo_n224 (.Z(FE_PHN3403_U_afifo_n224), 
	.A(U_afifo_n224));
   CLKBUF_X1 FE_PHC3402_U_afifo_n238 (.Z(FE_PHN3402_U_afifo_n238), 
	.A(U_afifo_n238));
   CLKBUF_X1 FE_PHC3401_U_afifo_U_acore_n77 (.Z(FE_PHN3401_U_afifo_U_acore_n77), 
	.A(U_afifo_U_acore_n77));
   CLKBUF_X1 FE_PHC3400_U_afifo_n250 (.Z(FE_PHN3400_U_afifo_n250), 
	.A(U_afifo_n250));
   CLKBUF_X1 FE_PHC3398_U_dfifo_U_dcore_n195 (.Z(FE_PHN3398_U_dfifo_U_dcore_n195), 
	.A(U_dfifo_U_dcore_n195));
   CLKBUF_X1 FE_PHC3397_U_afifo_n200 (.Z(FE_PHN3397_U_afifo_n200), 
	.A(U_afifo_n200));
   CLKBUF_X1 FE_PHC3396_U_afifo_n240 (.Z(FE_PHN3396_U_afifo_n240), 
	.A(U_afifo_n240));
   CLKBUF_X1 FE_PHC3395_U_afifo_n244 (.Z(FE_PHN3395_U_afifo_n244), 
	.A(U_afifo_n244));
   CLKBUF_X1 FE_PHC3394_U_afifo_n246 (.Z(FE_PHN3394_U_afifo_n246), 
	.A(U_afifo_n246));
   CLKBUF_X1 FE_PHC3393_U_afifo_n216 (.Z(FE_PHN3393_U_afifo_n216), 
	.A(U_afifo_n216));
   CLKBUF_X1 FE_PHC3392_U_afifo_n222 (.Z(FE_PHN3392_U_afifo_n222), 
	.A(U_afifo_n222));
   CLKBUF_X1 FE_PHC3390_U_afifo_n173 (.Z(FE_PHN3390_U_afifo_n173), 
	.A(U_afifo_n173));
   CLKBUF_X1 FE_PHC3388_U_afifo_n214 (.Z(FE_PHN3388_U_afifo_n214), 
	.A(U_afifo_n214));
   CLKBUF_X1 FE_PHC3386_U_afifo_U_acore_n71 (.Z(FE_PHN3386_U_afifo_U_acore_n71), 
	.A(U_afifo_U_acore_n71));
   CLKBUF_X1 FE_PHC3385_U_afifo_n228 (.Z(FE_PHN3385_U_afifo_n228), 
	.A(U_afifo_n228));
   CLKBUF_X1 FE_PHC3384_U_afifo_U_acore_n156 (.Z(FE_PHN3384_U_afifo_U_acore_n156), 
	.A(U_afifo_U_acore_n156));
   CLKBUF_X1 FE_PHC3383_U_afifo_n242 (.Z(FE_PHN3383_U_afifo_n242), 
	.A(U_afifo_n242));
   CLKBUF_X1 FE_PHC3382_U_ctl_n105 (.Z(FE_PHN3382_U_ctl_n105), 
	.A(U_ctl_n105));
   CLKBUF_X1 FE_PHC3381_U_afifo_n171 (.Z(FE_PHN3381_U_afifo_n171), 
	.A(U_afifo_n171));
   CLKBUF_X1 FE_PHC3380_U_afifo_U_acore_n73 (.Z(FE_PHN3380_U_afifo_U_acore_n73), 
	.A(U_afifo_U_acore_n73));
   CLKBUF_X1 FE_PHC3376_U_afifo_U_acore_n200 (.Z(FE_PHN3376_U_afifo_U_acore_n200), 
	.A(U_afifo_U_acore_n200));
   CLKBUF_X1 FE_PHC3374_U_afifo_f_clr_pers (.Z(FE_PHN3374_U_afifo_f_clr_pers), 
	.A(U_afifo_f_clr_pers));
   CLKBUF_X1 FE_PHC3372_U_dfifo_U_dcore_n178 (.Z(FE_PHN3372_U_dfifo_U_dcore_n178), 
	.A(U_dfifo_U_dcore_n178));
   CLKBUF_X1 FE_PHC3369_U_afifo_U_acore_n183 (.Z(FE_PHN3369_U_afifo_U_acore_n183), 
	.A(U_afifo_U_acore_n183));
   CLKBUF_X1 FE_PHC3368_U_dfifo_U_dcore_n192 (.Z(FE_PHN3368_U_dfifo_U_dcore_n192), 
	.A(U_dfifo_U_dcore_n192));
   CLKBUF_X1 FE_PHC3367_U_afifo_U_acore_n189 (.Z(FE_PHN3367_U_afifo_U_acore_n189), 
	.A(U_afifo_U_acore_n189));
   CLKBUF_X1 FE_PHC3366_U_afifo_U_acore_n180 (.Z(FE_PHN3366_U_afifo_U_acore_n180), 
	.A(U_afifo_U_acore_n180));
   CLKBUF_X1 FE_PHC3365_U_afifo_U_acore_n171 (.Z(FE_PHN3365_U_afifo_U_acore_n171), 
	.A(U_afifo_U_acore_n171));
   CLKBUF_X1 FE_PHC3364_U_dfifo_U_dcore_n180 (.Z(FE_PHN3364_U_dfifo_U_dcore_n180), 
	.A(U_dfifo_U_dcore_n180));
   CLKBUF_X1 FE_PHC3363_U_dfifo_U_dcore_n184 (.Z(FE_PHN3363_U_dfifo_U_dcore_n184), 
	.A(U_dfifo_U_dcore_n184));
   CLKBUF_X1 FE_PHC3362_U_afifo_U_acore_n193 (.Z(FE_PHN3362_U_afifo_U_acore_n193), 
	.A(U_afifo_U_acore_n193));
   CLKBUF_X1 FE_PHC3361_U_afifo_U_acore_n209 (.Z(FE_PHN3361_U_afifo_U_acore_n209), 
	.A(U_afifo_U_acore_n209));
   CLKBUF_X1 FE_PHC3360_U_afifo_U_acore_n182 (.Z(FE_PHN3360_U_afifo_U_acore_n182), 
	.A(U_afifo_U_acore_n182));
   CLKBUF_X1 FE_PHC3359_U_afifo_U_acore_n174 (.Z(FE_PHN3359_U_afifo_U_acore_n174), 
	.A(U_afifo_U_acore_n174));
   CLKBUF_X1 FE_PHC3358_U_dfifo_U_dcore_n176 (.Z(FE_PHN3358_U_dfifo_U_dcore_n176), 
	.A(U_dfifo_U_dcore_n176));
   CLKBUF_X1 FE_PHC3357_U_afifo_U_acore_f_afull (.Z(FE_PHN3357_U_afifo_U_acore_f_afull), 
	.A(U_afifo_U_acore_f_afull));
   CLKBUF_X1 FE_PHC3356_U_afifo_U_acore_n187 (.Z(FE_PHN3356_U_afifo_U_acore_n187), 
	.A(U_afifo_U_acore_n187));
   CLKBUF_X1 FE_PHC3354_U_dfifo_U_dcore_n181 (.Z(FE_PHN3354_U_dfifo_U_dcore_n181), 
	.A(U_dfifo_U_dcore_n181));
   CLKBUF_X1 FE_PHC3351_U_dfifo_U_dcore_n193 (.Z(FE_PHN3351_U_dfifo_U_dcore_n193), 
	.A(U_dfifo_U_dcore_n193));
   CLKBUF_X1 FE_PHC3350_U_afifo_U_acore_n206 (.Z(FE_PHN3350_U_afifo_U_acore_n206), 
	.A(U_afifo_U_acore_n206));
   CLKBUF_X1 FE_PHC3348_U_afifo_U_acore_n202 (.Z(FE_PHN3348_U_afifo_U_acore_n202), 
	.A(U_afifo_U_acore_n202));
   CLKBUF_X1 FE_PHC3347_U_afifo_U_acore_n172 (.Z(FE_PHN3347_U_afifo_U_acore_n172), 
	.A(U_afifo_U_acore_n172));
   CLKBUF_X1 FE_PHC3344_U_afifo_U_acore_n191 (.Z(FE_PHN3344_U_afifo_U_acore_n191), 
	.A(U_afifo_U_acore_n191));
   CLKBUF_X1 FE_PHC3342_U_afifo_U_acore_n196 (.Z(FE_PHN3342_U_afifo_U_acore_n196), 
	.A(U_afifo_U_acore_n196));
   CLKBUF_X1 FE_PHC3341_U_dfifo_U_dcore_n189 (.Z(FE_PHN3341_U_dfifo_U_dcore_n189), 
	.A(U_dfifo_U_dcore_n189));
   CLKBUF_X1 FE_PHC3340_U_afifo_U_acore_n185 (.Z(FE_PHN3340_U_afifo_U_acore_n185), 
	.A(U_afifo_U_acore_n185));
   CLKBUF_X1 FE_PHC3339_U_dfifo_U_dcore_n182 (.Z(FE_PHN3339_U_dfifo_U_dcore_n182), 
	.A(U_dfifo_U_dcore_n182));
   CLKBUF_X1 FE_PHC3338_U_dfifo_U_dcore_n186 (.Z(FE_PHN3338_U_dfifo_U_dcore_n186), 
	.A(U_dfifo_U_dcore_n186));
   CLKBUF_X1 FE_PHC3336_U_afifo_U_acore_n208 (.Z(FE_PHN3336_U_afifo_U_acore_n208), 
	.A(U_afifo_U_acore_n208));
   CLKBUF_X1 FE_PHC3335_U_afifo_U_acore_n178 (.Z(FE_PHN3335_U_afifo_U_acore_n178), 
	.A(U_afifo_U_acore_n178));
   CLKBUF_X1 FE_PHC3334_U_dfifo_U_dcore_n188 (.Z(FE_PHN3334_U_dfifo_U_dcore_n188), 
	.A(U_dfifo_U_dcore_n188));
   CLKBUF_X1 FE_PHC3333_U_afifo_U_acore_n176 (.Z(FE_PHN3333_U_afifo_U_acore_n176), 
	.A(U_afifo_U_acore_n176));
   CLKBUF_X1 FE_PHC3332_U_dfifo_U_dcore_n197 (.Z(FE_PHN3332_U_dfifo_U_dcore_n197), 
	.A(U_dfifo_U_dcore_n197));
   CLKBUF_X1 FE_PHC3331_U_afifo_U_acore_n204 (.Z(FE_PHN3331_U_afifo_U_acore_n204), 
	.A(U_afifo_U_acore_n204));
   CLKBUF_X1 FE_PHC3330_U_dfifo_U_dcore_n179 (.Z(FE_PHN3330_U_dfifo_U_dcore_n179), 
	.A(U_dfifo_U_dcore_n179));
   CLKBUF_X1 FE_PHC3329_U_dfifo_U_dcore_n191 (.Z(FE_PHN3329_U_dfifo_U_dcore_n191), 
	.A(U_dfifo_U_dcore_n191));
   CLKBUF_X1 FE_PHC3323_U_afifo_U_acore_n95 (.Z(FE_PHN3323_U_afifo_U_acore_n95), 
	.A(U_afifo_U_acore_n95));
   CLKBUF_X1 FE_PHC3310_U_afifo_U_acore_n97 (.Z(FE_PHN3310_U_afifo_U_acore_n97), 
	.A(U_afifo_U_acore_n97));
   CLKBUF_X1 FE_PHC3308_U_afifo_U_acore_U_sub_fifo_n273 (.Z(FE_PHN3308_U_afifo_U_acore_U_sub_fifo_n273), 
	.A(U_afifo_U_acore_U_sub_fifo_n273));
   CLKBUF_X1 FE_PHC3307_U_afifo_U_acore_U_sub_fifo_n202 (.Z(FE_PHN3307_U_afifo_U_acore_U_sub_fifo_n202), 
	.A(U_afifo_U_acore_U_sub_fifo_n202));
   BUF_X8 FE_PHC3306_U_afifo_U_acore_U_sub_fifo_n176 (.Z(FE_PHN3306_U_afifo_U_acore_U_sub_fifo_n176), 
	.A(U_afifo_U_acore_U_sub_fifo_n176));
   CLKBUF_X1 FE_PHC3304_U_afifo_U_acore_U_sub_fifo_n277 (.Z(FE_PHN3304_U_afifo_U_acore_U_sub_fifo_n277), 
	.A(U_afifo_U_acore_U_sub_fifo_n277));
   CLKBUF_X1 FE_PHC3303_U_afifo_U_acore_U_sub_fifo_n203 (.Z(FE_PHN3303_U_afifo_U_acore_U_sub_fifo_n203), 
	.A(U_afifo_U_acore_U_sub_fifo_n203));
   BUF_X8 FE_PHC3302_U_afifo_U_acore_U_sub_fifo_n206 (.Z(FE_PHN3302_U_afifo_U_acore_U_sub_fifo_n206), 
	.A(U_afifo_U_acore_U_sub_fifo_n206));
   BUF_X8 FE_PHC3301_U_afifo_U_acore_U_sub_fifo_n201 (.Z(FE_PHN3301_U_afifo_U_acore_U_sub_fifo_n201), 
	.A(U_afifo_U_acore_U_sub_fifo_n201));
   BUF_X8 FE_PHC3300_U_afifo_U_acore_U_sub_fifo_n200 (.Z(FE_PHN3300_U_afifo_U_acore_U_sub_fifo_n200), 
	.A(U_afifo_U_acore_U_sub_fifo_n200));
   BUF_X8 FE_PHC3296_U_afifo_U_acore_U_sub_fifo_n198 (.Z(FE_PHN3296_U_afifo_U_acore_U_sub_fifo_n198), 
	.A(U_afifo_U_acore_U_sub_fifo_n198));
   CLKBUF_X1 FE_PHC3295_U_dfifo_U_dcore_U_sub_fifo_n450 (.Z(FE_PHN3295_U_dfifo_U_dcore_U_sub_fifo_n450), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n450));
   BUF_X8 FE_PHC3294_U_afifo_U_acore_U_sub_fifo_n249 (.Z(FE_PHN3294_U_afifo_U_acore_U_sub_fifo_n249), 
	.A(U_afifo_U_acore_U_sub_fifo_n249));
   BUF_X8 FE_PHC3285_U_afifo_U_acore_U_sub_fifo_n269 (.Z(FE_PHN3285_U_afifo_U_acore_U_sub_fifo_n269), 
	.A(U_afifo_U_acore_U_sub_fifo_n269));
   BUF_X16 FE_PHC3284_U_dfifo_n3 (.Z(FE_PHN3284_U_dfifo_n3), 
	.A(U_dfifo_n3));
   BUF_X32 FE_PHC3281_U_rbuf_n82 (.Z(FE_PHN3281_U_rbuf_n82), 
	.A(U_rbuf_n82));
   BUF_X32 FE_PHC3280_U_rbuf_n84 (.Z(FE_PHN3280_U_rbuf_n84), 
	.A(U_rbuf_n84));
   BUF_X32 FE_PHC3279_U_rbuf_n85 (.Z(FE_PHN3279_U_rbuf_n85), 
	.A(U_rbuf_n85));
   BUF_X32 FE_PHC3272_U_rbuf_n71 (.Z(FE_PHN3272_U_rbuf_n71), 
	.A(U_rbuf_n71));
   BUF_X32 FE_PHC3271_U_ctl_n141 (.Z(FE_PHN3271_U_ctl_n141), 
	.A(U_ctl_n141));
   BUF_X32 FE_PHC3270_U_ctl_n123 (.Z(FE_PHN3270_U_ctl_n123), 
	.A(U_ctl_n123));
   BUF_X32 FE_PHC3269_U_ctl_n139 (.Z(FE_PHN3269_U_ctl_n139), 
	.A(U_ctl_n139));
   CLKBUF_X1 FE_PHC3267_U_afifo_U_acore_n142 (.Z(FE_PHN3267_U_afifo_U_acore_n142), 
	.A(U_afifo_U_acore_n142));
   CLKBUF_X1 FE_PHC3266_U_dfifo_U_dcore_n167 (.Z(FE_PHN3266_U_dfifo_U_dcore_n167), 
	.A(U_dfifo_U_dcore_n167));
   CLKBUF_X1 FE_PHC3265_U_afifo_U_acore_n144 (.Z(FE_PHN3265_U_afifo_U_acore_n144), 
	.A(U_afifo_U_acore_n144));
   CLKBUF_X1 FE_PHC3264_U_afifo_U_acore_n138 (.Z(FE_PHN3264_U_afifo_U_acore_n138), 
	.A(U_afifo_U_acore_n138));
   CLKBUF_X1 FE_PHC3263_U_afifo_U_acore_n162 (.Z(FE_PHN3263_U_afifo_U_acore_n162), 
	.A(U_afifo_U_acore_n162));
   BUF_X1 FE_PHC3262_U_afifo_U_acore_n160 (.Z(FE_PHN3262_U_afifo_U_acore_n160), 
	.A(U_afifo_U_acore_n160));
   CLKBUF_X1 FE_PHC3261_U_afifo_U_acore_n33 (.Z(FE_PHN3261_U_afifo_U_acore_n33), 
	.A(U_afifo_U_acore_n33));
   BUF_X1 FE_PHC3257_U_afifo_U_acore_n104 (.Z(FE_PHN3257_U_afifo_U_acore_n104), 
	.A(U_afifo_U_acore_n104));
   CLKBUF_X1 FE_PHC3254_U_afifo_U_acore_n121 (.Z(FE_PHN3254_U_afifo_U_acore_n121), 
	.A(U_afifo_U_acore_n121));
   CLKBUF_X1 FE_PHC3253_U_afifo_U_acore_n115 (.Z(FE_PHN3253_U_afifo_U_acore_n115), 
	.A(U_afifo_U_acore_n115));
   CLKBUF_X1 FE_PHC3251_U_afifo_U_acore_n147 (.Z(FE_PHN3251_U_afifo_U_acore_n147), 
	.A(U_afifo_U_acore_n147));
   CLKBUF_X1 FE_PHC3248_U_afifo_U_acore_n94 (.Z(FE_PHN3248_U_afifo_U_acore_n94), 
	.A(U_afifo_U_acore_n94));
   CLKBUF_X1 FE_PHC3246_U_dfifo_U_dcore_f_buf_data_0_ (.Z(FE_PHN3246_U_dfifo_U_dcore_f_buf_data_0_), 
	.A(U_dfifo_U_dcore_f_buf_data_0_));
   CLKBUF_X1 FE_PHC3243_U_afifo_U_acore_n199 (.Z(FE_PHN3243_U_afifo_U_acore_n199), 
	.A(U_afifo_U_acore_n199));
   CLKBUF_X1 FE_PHC3236_U_dfifo_U_dcore_n157 (.Z(FE_PHN3236_U_dfifo_U_dcore_n157), 
	.A(U_dfifo_U_dcore_n157));
   BUF_X8 FE_PHC3226_U_dfifo_U_dcore_n155 (.Z(FE_PHN3226_U_dfifo_U_dcore_n155), 
	.A(U_dfifo_U_dcore_n155));
   CLKBUF_X1 FE_PHC3225_U_afifo_m_data_in_14_ (.Z(FE_PHN3225_U_afifo_m_data_in_14_), 
	.A(U_afifo_m_data_in[14]));
   BUF_X8 FE_PHC3219_U_dfifo_U_dcore_n145 (.Z(FE_PHN3219_U_dfifo_U_dcore_n145), 
	.A(U_dfifo_U_dcore_n145));
   BUF_X8 FE_PHC3218_U_dfifo_U_dcore_U_sub_fifo_n452 (.Z(FE_PHN3218_U_dfifo_U_dcore_U_sub_fifo_n452), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n452));
   BUF_X16 FE_PHC3214_U_dfifo_U_dcore_n148 (.Z(FE_PHN3214_U_dfifo_U_dcore_n148), 
	.A(U_dfifo_U_dcore_n148));
   BUF_X16 FE_PHC3213_U_afifo_m_data_in_12_ (.Z(FE_PHN3213_U_afifo_m_data_in_12_), 
	.A(U_afifo_m_data_in[12]));
   BUF_X32 FE_PHC3210_U_afifo_m_data_in_4_ (.Z(FE_PHN3210_U_afifo_m_data_in_4_), 
	.A(U_afifo_m_data_in[4]));
   BUF_X32 FE_PHC3207_U_ctl_n117 (.Z(FE_PHN3207_U_ctl_n117), 
	.A(U_ctl_n117));
   BUF_X32 FE_PHC3203_U_ctl_n120 (.Z(FE_PHN3203_U_ctl_n120), 
	.A(U_ctl_n120));
   CLKBUF_X1 FE_PHC3184_U_afifo_U_acore_U_sub_fifo_n287 (.Z(FE_PHN3184_U_afifo_U_acore_U_sub_fifo_n287), 
	.A(U_afifo_U_acore_U_sub_fifo_n287));
   CLKBUF_X1 FE_PHC3181_U_afifo_U_acore_U_sub_fifo_n322 (.Z(FE_PHN3181_U_afifo_U_acore_U_sub_fifo_n322), 
	.A(U_afifo_U_acore_U_sub_fifo_n322));
   CLKBUF_X1 FE_PHC3180_U_afifo_U_acore_n133 (.Z(FE_PHN3180_U_afifo_U_acore_n133), 
	.A(FE_PHN1314_U_afifo_U_acore_n133));
   CLKBUF_X1 FE_PHC3179_U_afifo_U_acore_U_sub_fifo_n305 (.Z(FE_PHN3179_U_afifo_U_acore_U_sub_fifo_n305), 
	.A(U_afifo_U_acore_U_sub_fifo_n305));
   CLKBUF_X1 FE_PHC3178_U_afifo_U_acore_U_sub_fifo_n292 (.Z(FE_PHN3178_U_afifo_U_acore_U_sub_fifo_n292), 
	.A(U_afifo_U_acore_U_sub_fifo_n292));
   CLKBUF_X1 FE_PHC3177_U_afifo_U_acore_U_sub_fifo_n310 (.Z(FE_PHN3177_U_afifo_U_acore_U_sub_fifo_n310), 
	.A(U_afifo_U_acore_U_sub_fifo_n310));
   CLKBUF_X1 FE_PHC3176_U_afifo_U_acore_U_sub_fifo_n316 (.Z(FE_PHN3176_U_afifo_U_acore_U_sub_fifo_n316), 
	.A(U_afifo_U_acore_U_sub_fifo_n316));
   CLKBUF_X1 FE_PHC3175_U_afifo_U_acore_U_sub_fifo_n297 (.Z(FE_PHN3175_U_afifo_U_acore_U_sub_fifo_n297), 
	.A(U_afifo_U_acore_U_sub_fifo_n297));
   CLKBUF_X1 FE_PHC3174_U_afifo_U_acore_U_sub_fifo_n294 (.Z(FE_PHN3174_U_afifo_U_acore_U_sub_fifo_n294), 
	.A(U_afifo_U_acore_U_sub_fifo_n294));
   CLKBUF_X1 FE_PHC3173_U_afifo_U_acore_U_sub_fifo_n278 (.Z(FE_PHN3173_U_afifo_U_acore_U_sub_fifo_n278), 
	.A(U_afifo_U_acore_U_sub_fifo_n278));
   CLKBUF_X1 FE_PHC3172_U_afifo_U_acore_U_sub_fifo_n274 (.Z(FE_PHN3172_U_afifo_U_acore_U_sub_fifo_n274), 
	.A(U_afifo_U_acore_U_sub_fifo_n274));
   CLKBUF_X1 FE_PHC3171_U_afifo_U_acore_U_sub_fifo_n308 (.Z(FE_PHN3171_U_afifo_U_acore_U_sub_fifo_n308), 
	.A(U_afifo_U_acore_U_sub_fifo_n308));
   BUF_X8 FE_PHC3163_U_afifo_U_acore_U_sub_fifo_n296 (.Z(FE_PHN3163_U_afifo_U_acore_U_sub_fifo_n296), 
	.A(U_afifo_U_acore_U_sub_fifo_n296));
   BUF_X16 FE_PHC3161_U_afifo_U_acore_U_sub_fifo_n295 (.Z(FE_PHN3161_U_afifo_U_acore_U_sub_fifo_n295), 
	.A(U_afifo_U_acore_U_sub_fifo_n295));
   BUF_X16 FE_PHC3159_U_afifo_U_acore_U_sub_fifo_n280 (.Z(FE_PHN3159_U_afifo_U_acore_U_sub_fifo_n280), 
	.A(U_afifo_U_acore_U_sub_fifo_n280));
   BUF_X16 FE_PHC3158_U_afifo_U_acore_U_sub_fifo_n318 (.Z(FE_PHN3158_U_afifo_U_acore_U_sub_fifo_n318), 
	.A(U_afifo_U_acore_U_sub_fifo_n318));
   BUF_X16 FE_PHC3157_U_afifo_U_acore_U_sub_fifo_n307 (.Z(FE_PHN3157_U_afifo_U_acore_U_sub_fifo_n307), 
	.A(U_afifo_U_acore_U_sub_fifo_n307));
   BUF_X32 FE_PHC3155_U_ctl_n133 (.Z(FE_PHN3155_U_ctl_n133), 
	.A(U_ctl_n133));
   BUF_X32 FE_PHC3154_U_ctl_n134 (.Z(FE_PHN3154_U_ctl_n134), 
	.A(U_ctl_n134));
   BUF_X32 FE_PHC3152_U_ctl_n118 (.Z(FE_PHN3152_U_ctl_n118), 
	.A(FE_PHN1605_U_ctl_n118));
   BUF_X32 FE_PHC3151_U_ctl_n130 (.Z(FE_PHN3151_U_ctl_n130), 
	.A(U_ctl_n130));
   BUF_X32 FE_PHC3150_U_ctl_n137 (.Z(FE_PHN3150_U_ctl_n137), 
	.A(U_ctl_n137));
   BUF_X32 FE_PHC3149_U_ctl_n140 (.Z(FE_PHN3149_U_ctl_n140), 
	.A(U_ctl_n140));
   BUF_X32 FE_PHC3148_U_ctl_n129 (.Z(FE_PHN3148_U_ctl_n129), 
	.A(U_ctl_n129));
   BUF_X32 FE_PHC3147_U_ctl_n131 (.Z(FE_PHN3147_U_ctl_n131), 
	.A(U_ctl_n131));
   BUF_X32 FE_PHC3146_U_ctl_n128 (.Z(FE_PHN3146_U_ctl_n128), 
	.A(U_ctl_n128));
   BUF_X32 FE_PHC3145_U_ctl_n125 (.Z(FE_PHN3145_U_ctl_n125), 
	.A(U_ctl_n125));
   BUF_X32 FE_PHC3144_U_ctl_n106 (.Z(FE_PHN3144_U_ctl_n106), 
	.A(U_ctl_n106));
   BUF_X32 FE_PHC3141_U_ctl_n421 (.Z(FE_PHN3141_U_ctl_n421), 
	.A(FE_PHN1675_U_ctl_n421));
   CLKBUF_X1 FE_PHC3132_U_dfifo_U_dcore_n139 (.Z(FE_PHN3132_U_dfifo_U_dcore_n139), 
	.A(U_dfifo_U_dcore_n139));
   CLKBUF_X1 FE_PHC3131_U_dfifo_U_dcore_n141 (.Z(FE_PHN3131_U_dfifo_U_dcore_n141), 
	.A(U_dfifo_U_dcore_n141));
   CLKBUF_X1 FE_PHC3130_U_dfifo_U_dcore_n137 (.Z(FE_PHN3130_U_dfifo_U_dcore_n137), 
	.A(U_dfifo_U_dcore_n137));
   CLKBUF_X1 FE_PHC3129_U_dfifo_U_dcore_n138 (.Z(FE_PHN3129_U_dfifo_U_dcore_n138), 
	.A(U_dfifo_U_dcore_n138));
   CLKBUF_X1 FE_PHC3128_U_dfifo_U_dcore_n135 (.Z(FE_PHN3128_U_dfifo_U_dcore_n135), 
	.A(U_dfifo_U_dcore_n135));
   CLKBUF_X1 FE_PHC3125_U_dfifo_U_dcore_n203 (.Z(FE_PHN3125_U_dfifo_U_dcore_n203), 
	.A(FE_PHN1498_U_dfifo_U_dcore_n203));
   CLKBUF_X1 FE_PHC3124_U_dfifo_U_dcore_f_buf_data_6_ (.Z(FE_PHN3124_U_dfifo_U_dcore_f_buf_data_6_), 
	.A(U_dfifo_U_dcore_f_buf_data_6_));
   CLKBUF_X1 FE_PHC3122_U_dfifo_U_dcore_f_buf_data_19_ (.Z(FE_PHN3122_U_dfifo_U_dcore_f_buf_data_19_), 
	.A(U_dfifo_U_dcore_f_buf_data_19_));
   CLKBUF_X1 FE_PHC3121_U_dfifo_U_dcore_f_buf_data_7_ (.Z(FE_PHN3121_U_dfifo_U_dcore_f_buf_data_7_), 
	.A(U_dfifo_U_dcore_f_buf_data_7_));
   CLKBUF_X1 FE_PHC3120_U_dfifo_U_dcore_f_buf_data_3_ (.Z(FE_PHN3120_U_dfifo_U_dcore_f_buf_data_3_), 
	.A(U_dfifo_U_dcore_f_buf_data_3_));
   CLKBUF_X1 FE_PHC3118_U_dfifo_U_dcore_f_buf_data_15_ (.Z(FE_PHN3118_U_dfifo_U_dcore_f_buf_data_15_), 
	.A(U_dfifo_U_dcore_f_buf_data_15_));
   CLKBUF_X1 FE_PHC3117_U_dfifo_U_dcore_f_buf_data_17_ (.Z(FE_PHN3117_U_dfifo_U_dcore_f_buf_data_17_), 
	.A(U_dfifo_U_dcore_f_buf_data_17_));
   CLKBUF_X1 FE_PHC3116_U_dfifo_U_dcore_f_buf_data_22_ (.Z(FE_PHN3116_U_dfifo_U_dcore_f_buf_data_22_), 
	.A(U_dfifo_U_dcore_f_buf_data_22_));
   CLKBUF_X1 FE_PHC3114_U_dfifo_U_dcore_f_buf_data_9_ (.Z(FE_PHN3114_U_dfifo_U_dcore_f_buf_data_9_), 
	.A(U_dfifo_U_dcore_f_buf_data_9_));
   BUF_X32 FE_PHC3096_U_ctl_n135 (.Z(FE_PHN3096_U_ctl_n135), 
	.A(U_ctl_n135));
   BUF_X32 FE_PHC3095_U_ctl_n119 (.Z(FE_PHN3095_U_ctl_n119), 
	.A(U_ctl_n119));
   BUF_X32 FE_PHC3062_U_ctl_n122 (.Z(FE_PHN3062_U_ctl_n122), 
	.A(U_ctl_n122));
   BUF_X32 FE_PHC3042_U_ctl_n138 (.Z(FE_PHN3042_U_ctl_n138), 
	.A(U_ctl_n138));
   CLKBUF_X1 FE_PHC3040_U_dfifo_U_dcore_f_buf_data_30_ (.Z(FE_PHN3040_U_dfifo_U_dcore_f_buf_data_30_), 
	.A(U_dfifo_U_dcore_f_buf_data_30_));
   CLKBUF_X1 FE_PHC3039_U_dfifo_U_dcore_f_buf_data_2_ (.Z(FE_PHN3039_U_dfifo_U_dcore_f_buf_data_2_), 
	.A(U_dfifo_U_dcore_f_buf_data_2_));
   CLKBUF_X1 FE_PHC3038_U_dfifo_U_dcore_f_buf_data_5_ (.Z(FE_PHN3038_U_dfifo_U_dcore_f_buf_data_5_), 
	.A(U_dfifo_U_dcore_f_buf_data_5_));
   CLKBUF_X1 FE_PHC3037_U_dfifo_U_dcore_f_buf_data_31_ (.Z(FE_PHN3037_U_dfifo_U_dcore_f_buf_data_31_), 
	.A(U_dfifo_U_dcore_f_buf_data_31_));
   CLKBUF_X1 FE_PHC3036_U_dfifo_U_dcore_f_buf_data_4_ (.Z(FE_PHN3036_U_dfifo_U_dcore_f_buf_data_4_), 
	.A(U_dfifo_U_dcore_f_buf_data_4_));
   CLKBUF_X1 FE_PHC3035_U_dfifo_U_dcore_f_buf_data_28_ (.Z(FE_PHN3035_U_dfifo_U_dcore_f_buf_data_28_), 
	.A(U_dfifo_U_dcore_f_buf_data_28_));
   BUF_X8 FE_PHC3032_U_afifo_n_new_req (.Z(FE_PHN3032_U_afifo_n_new_req), 
	.A(U_afifo_n_new_req));
   BUF_X32 FE_PHC3027_U_rbuf_n63 (.Z(FE_PHN3027_U_rbuf_n63), 
	.A(FE_PHN5180_U_rbuf_n63));
   BUF_X32 FE_PHC3026_U_rbuf_n64 (.Z(FE_PHN3026_U_rbuf_n64), 
	.A(U_rbuf_n64));
   BUF_X32 FE_PHC3025_U_rbuf_n83 (.Z(FE_PHN3025_U_rbuf_n83), 
	.A(U_rbuf_n83));
   BUF_X32 FE_PHC3024_U_rbuf_n65 (.Z(FE_PHN3024_U_rbuf_n65), 
	.A(U_rbuf_n65));
   BUF_X32 FE_PHC3023_U_rbuf_n72 (.Z(FE_PHN3023_U_rbuf_n72), 
	.A(FE_PHN5179_U_rbuf_n72));
   BUF_X32 FE_PHC3022_U_rbuf_n59 (.Z(FE_PHN3022_U_rbuf_n59), 
	.A(FE_PHN4649_U_rbuf_n59));
   BUF_X32 FE_PHC3021_U_rbuf_n77 (.Z(FE_PHN3021_U_rbuf_n77), 
	.A(U_rbuf_n77));
   BUF_X32 FE_PHC3020_U_rbuf_n60 (.Z(FE_PHN3020_U_rbuf_n60), 
	.A(U_rbuf_n60));
   BUF_X32 FE_PHC3019_U_rbuf_n80 (.Z(FE_PHN3019_U_rbuf_n80), 
	.A(U_rbuf_n80));
   BUF_X32 FE_PHC3017_U_rbuf_n76 (.Z(FE_PHN3017_U_rbuf_n76), 
	.A(U_rbuf_n76));
   BUF_X32 FE_PHC3016_U_rbuf_n81 (.Z(FE_PHN3016_U_rbuf_n81), 
	.A(U_rbuf_n81));
   BUF_X32 FE_PHC3015_U_rbuf_n74 (.Z(FE_PHN3015_U_rbuf_n74), 
	.A(U_rbuf_n74));
   BUF_X32 FE_PHC3014_U_ctl_n124 (.Z(FE_PHN3014_U_ctl_n124), 
	.A(U_ctl_n124));
   BUF_X32 FE_PHC3008_U_rbuf_n56 (.Z(FE_PHN3008_U_rbuf_n56), 
	.A(FE_PHN4643_U_rbuf_n56));
   BUF_X32 FE_PHC3007_U_rbuf_n67 (.Z(FE_PHN3007_U_rbuf_n67), 
	.A(U_rbuf_n67));
   BUF_X32 FE_PHC3006_U_rbuf_n61 (.Z(FE_PHN3006_U_rbuf_n61), 
	.A(U_rbuf_n61));
   BUF_X32 FE_PHC3005_U_rbuf_n70 (.Z(FE_PHN3005_U_rbuf_n70), 
	.A(U_rbuf_n70));
   BUF_X32 FE_PHC3004_U_rbuf_n57 (.Z(FE_PHN3004_U_rbuf_n57), 
	.A(U_rbuf_n57));
   BUF_X32 FE_PHC3003_U_rbuf_n58 (.Z(FE_PHN3003_U_rbuf_n58), 
	.A(U_rbuf_n58));
   BUF_X32 FE_PHC3002_hiu_terminate (.Z(FE_PHN3002_hiu_terminate), 
	.A(FE_PHN676_hiu_terminate));
   BUF_X32 FE_PHC2999_U_rbuf_n73 (.Z(FE_PHN2999_U_rbuf_n73), 
	.A(U_rbuf_n73));
   BUF_X32 FE_PHC2998_U_rbuf_n86 (.Z(FE_PHN2998_U_rbuf_n86), 
	.A(U_rbuf_n86));
   BUF_X32 FE_PHC2997_U_rbuf_n79 (.Z(FE_PHN2997_U_rbuf_n79), 
	.A(U_rbuf_n79));
   BUF_X32 FE_PHC2996_U_rbuf_n75 (.Z(FE_PHN2996_U_rbuf_n75), 
	.A(FE_PHN4642_U_rbuf_n75));
   CLKBUF_X1 FE_PHC2979_U_afifo_U_acore_U_sub_fifo_count_0_ (.Z(FE_PHN2979_U_afifo_U_acore_U_sub_fifo_count_0_), 
	.A(U_afifo_U_acore_U_sub_fifo_count_0_));
   BUF_X32 FE_PHC2963_U_ctl_n132 (.Z(FE_PHN2963_U_ctl_n132), 
	.A(U_ctl_n132));
   BUF_X32 FE_PHC2957_U_rbuf_n62 (.Z(FE_PHN2957_U_rbuf_n62), 
	.A(U_rbuf_n62));
   BUF_X32 FE_PHC2949_U_rbuf_n78 (.Z(FE_PHN2949_U_rbuf_n78), 
	.A(U_rbuf_n78));
   BUF_X32 FE_PHC2940_U_rbuf_n55 (.Z(FE_PHN2940_U_rbuf_n55), 
	.A(U_rbuf_n55));
   BUF_X32 FE_PHC2938_U_rbuf_n69 (.Z(FE_PHN2938_U_rbuf_n69), 
	.A(FE_PHN4665_U_rbuf_n69));
   BUF_X32 FE_PHC2937_U_rbuf_n66 (.Z(FE_PHN2937_U_rbuf_n66), 
	.A(U_rbuf_n66));
   BUF_X32 FE_PHC2934_U_rbuf_n68 (.Z(FE_PHN2934_U_rbuf_n68), 
	.A(U_rbuf_n68));
   BUF_X32 FE_PHC2933_U_ctl_n127 (.Z(FE_PHN2933_U_ctl_n127), 
	.A(U_ctl_n127));
   BUF_X32 FE_PHC2930_U_rbuf_n89 (.Z(FE_PHN2930_U_rbuf_n89), 
	.A(FE_PHN782_U_rbuf_n89));
   BUF_X32 FE_PHC2924_m_rb_overflow (.Z(FE_PHN2924_m_rb_overflow), 
	.A(m_rb_overflow));
   BUF_X32 FE_PHC2923_U_ctl_n212 (.Z(FE_PHN2923_U_ctl_n212), 
	.A(FE_PHN4633_U_ctl_n212));
   BUF_X32 FE_PHC2917_hsel_reg (.Z(FE_PHN2917_hsel_reg), 
	.A(FE_PHN695_hsel_reg));
   BUF_X32 FE_PHC2914_U_ctl_n382 (.Z(FE_PHN2914_U_ctl_n382), 
	.A(FE_PHN4628_U_ctl_n382));
   BUF_X2 FE_PHC2913_U_ctl_n422 (.Z(FE_PHN2913_U_ctl_n422), 
	.A(FE_PHN687_U_ctl_n422));
   BUF_X32 FE_PHC2908_m_af_push1_n (.Z(FE_PHN2908_m_af_push1_n), 
	.A(FE_PHN4626_m_af_push1_n));
   BUF_X32 FE_PHC2904_U_ctl_f_burst_done (.Z(FE_PHN2904_U_ctl_f_burst_done), 
	.A(FE_PHN4619_U_ctl_f_burst_done));
   BUF_X32 FE_PHC2704_U_afifo_n20 (.Z(FE_PHN2704_U_afifo_n20), 
	.A(FE_PHN3770_U_afifo_n20));
   BUF_X32 FE_PHC2677_U_afifo_n19 (.Z(FE_PHN2677_U_afifo_n19), 
	.A(FE_PHN3646_U_afifo_n19));
   BUF_X32 FE_PHC2656_U_afifo_n18 (.Z(FE_PHN2656_U_afifo_n18), 
	.A(FE_PHN3671_U_afifo_n18));
   BUF_X32 FE_PHC2638_U_afifo_n159 (.Z(FE_PHN2638_U_afifo_n159), 
	.A(FE_PHN5100_U_afifo_n159));
   BUF_X32 FE_PHC2575_U_afifo_n166 (.Z(FE_PHN2575_U_afifo_n166), 
	.A(FE_PHN5021_U_afifo_n166));
   BUF_X32 FE_PHC2567_U_afifo_n165 (.Z(FE_PHN2567_U_afifo_n165), 
	.A(FE_PHN5004_U_afifo_n165));
   BUF_X32 FE_PHC2565_U_afifo_n191 (.Z(FE_PHN2565_U_afifo_n191), 
	.A(FE_PHN4917_U_afifo_n191));
   BUF_X32 FE_PHC2558_U_afifo_n160 (.Z(FE_PHN2558_U_afifo_n160), 
	.A(U_afifo_n160));
   BUF_X32 FE_PHC2434_U_afifo_n158 (.Z(FE_PHN2434_U_afifo_n158), 
	.A(FE_PHN5132_U_afifo_n158));
   BUF_X32 FE_PHC2433_U_afifo_n164 (.Z(FE_PHN2433_U_afifo_n164), 
	.A(FE_PHN3543_U_afifo_n164));
   BUF_X16 FE_PHC2421_U_dfifo_U_dcore_U_sub_fifo_n448 (.Z(FE_PHN2421_U_dfifo_U_dcore_U_sub_fifo_n448), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n448));
   BUF_X32 FE_PHC2375_U_dfifo_U_dcore_U_sub_fifo_n272 (.Z(FE_PHN2375_U_dfifo_U_dcore_U_sub_fifo_n272), 
	.A(FE_PHN4370_U_dfifo_U_dcore_U_sub_fifo_n272));
   BUF_X32 FE_PHC2374_U_dfifo_U_dcore_U_sub_fifo_n271 (.Z(FE_PHN2374_U_dfifo_U_dcore_U_sub_fifo_n271), 
	.A(FE_PHN4292_U_dfifo_U_dcore_U_sub_fifo_n271));
   BUF_X32 FE_PHC2372_U_dfifo_U_dcore_U_sub_fifo_n303 (.Z(FE_PHN2372_U_dfifo_U_dcore_U_sub_fifo_n303), 
	.A(FE_PHN4347_U_dfifo_U_dcore_U_sub_fifo_n303));
   BUF_X32 FE_PHC2371_U_dfifo_U_dcore_U_sub_fifo_n306 (.Z(FE_PHN2371_U_dfifo_U_dcore_U_sub_fifo_n306), 
	.A(FE_PHN4300_U_dfifo_U_dcore_U_sub_fifo_n306));
   BUF_X32 FE_PHC2370_U_dfifo_U_dcore_U_sub_fifo_n294 (.Z(FE_PHN2370_U_dfifo_U_dcore_U_sub_fifo_n294), 
	.A(FE_PHN4285_U_dfifo_U_dcore_U_sub_fifo_n294));
   BUF_X32 FE_PHC2369_U_dfifo_U_dcore_U_sub_fifo_n260 (.Z(FE_PHN2369_U_dfifo_U_dcore_U_sub_fifo_n260), 
	.A(FE_PHN4284_U_dfifo_U_dcore_U_sub_fifo_n260));
   BUF_X32 FE_PHC2368_U_dfifo_U_dcore_U_sub_fifo_n295 (.Z(FE_PHN2368_U_dfifo_U_dcore_U_sub_fifo_n295), 
	.A(FE_PHN4275_U_dfifo_U_dcore_U_sub_fifo_n295));
   BUF_X32 FE_PHC2367_U_dfifo_U_dcore_U_sub_fifo_n309 (.Z(FE_PHN2367_U_dfifo_U_dcore_U_sub_fifo_n309), 
	.A(FE_PHN4252_U_dfifo_U_dcore_U_sub_fifo_n309));
   BUF_X32 FE_PHC2366_U_dfifo_U_dcore_U_sub_fifo_n278 (.Z(FE_PHN2366_U_dfifo_U_dcore_U_sub_fifo_n278), 
	.A(FE_PHN4309_U_dfifo_U_dcore_U_sub_fifo_n278));
   BUF_X32 FE_PHC2365_U_dfifo_U_dcore_U_sub_fifo_n305 (.Z(FE_PHN2365_U_dfifo_U_dcore_U_sub_fifo_n305), 
	.A(FE_PHN4243_U_dfifo_U_dcore_U_sub_fifo_n305));
   BUF_X32 FE_PHC2363_U_dfifo_U_dcore_U_sub_fifo_n275 (.Z(FE_PHN2363_U_dfifo_U_dcore_U_sub_fifo_n275), 
	.A(FE_PHN5159_U_dfifo_U_dcore_U_sub_fifo_n275));
   BUF_X32 FE_PHC2362_U_afifo_U_acore_U_sub_fifo_n248 (.Z(FE_PHN2362_U_afifo_U_acore_U_sub_fifo_n248), 
	.A(FE_PHN3499_U_afifo_U_acore_U_sub_fifo_n248));
   BUF_X32 FE_PHC2361_U_dfifo_U_dcore_U_sub_fifo_n269 (.Z(FE_PHN2361_U_dfifo_U_dcore_U_sub_fifo_n269), 
	.A(FE_PHN4245_U_dfifo_U_dcore_U_sub_fifo_n269));
   BUF_X32 FE_PHC2360_U_dfifo_U_dcore_U_sub_fifo_n270 (.Z(FE_PHN2360_U_dfifo_U_dcore_U_sub_fifo_n270), 
	.A(FE_PHN4290_U_dfifo_U_dcore_U_sub_fifo_n270));
   BUF_X32 FE_PHC2359_U_afifo_U_acore_U_sub_fifo_n197 (.Z(FE_PHN2359_U_afifo_U_acore_U_sub_fifo_n197), 
	.A(FE_PHN4036_U_afifo_U_acore_U_sub_fifo_n197));
   BUF_X32 FE_PHC2358_U_dfifo_U_dcore_U_sub_fifo_n283 (.Z(FE_PHN2358_U_dfifo_U_dcore_U_sub_fifo_n283), 
	.A(FE_PHN4276_U_dfifo_U_dcore_U_sub_fifo_n283));
   BUF_X32 FE_PHC2357_U_dfifo_U_dcore_U_sub_fifo_n268 (.Z(FE_PHN2357_U_dfifo_U_dcore_U_sub_fifo_n268), 
	.A(FE_PHN4253_U_dfifo_U_dcore_U_sub_fifo_n268));
   BUF_X32 FE_PHC2356_U_dfifo_U_dcore_U_sub_fifo_n307 (.Z(FE_PHN2356_U_dfifo_U_dcore_U_sub_fifo_n307), 
	.A(FE_PHN5138_U_dfifo_U_dcore_U_sub_fifo_n307));
   BUF_X32 FE_PHC2354_U_dfifo_U_dcore_U_sub_fifo_n292 (.Z(FE_PHN2354_U_dfifo_U_dcore_U_sub_fifo_n292), 
	.A(FE_PHN5115_U_dfifo_U_dcore_U_sub_fifo_n292));
   BUF_X32 FE_PHC2353_U_dfifo_U_dcore_U_sub_fifo_n257 (.Z(FE_PHN2353_U_dfifo_U_dcore_U_sub_fifo_n257), 
	.A(FE_PHN5148_U_dfifo_U_dcore_U_sub_fifo_n257));
   BUF_X32 FE_PHC2352_U_dfifo_U_dcore_U_sub_fifo_n253 (.Z(FE_PHN2352_U_dfifo_U_dcore_U_sub_fifo_n253), 
	.A(FE_PHN4939_U_dfifo_U_dcore_U_sub_fifo_n253));
   BUF_X32 FE_PHC2351_U_afifo_U_acore_U_sub_fifo_n208 (.Z(FE_PHN2351_U_afifo_U_acore_U_sub_fifo_n208), 
	.A(FE_PHN4197_U_afifo_U_acore_U_sub_fifo_n208));
   BUF_X32 FE_PHC2350_U_dfifo_U_dcore_U_sub_fifo_n279 (.Z(FE_PHN2350_U_dfifo_U_dcore_U_sub_fifo_n279), 
	.A(FE_PHN4993_U_dfifo_U_dcore_U_sub_fifo_n279));
   BUF_X32 FE_PHC2349_U_dfifo_U_dcore_U_sub_fifo_n265 (.Z(FE_PHN2349_U_dfifo_U_dcore_U_sub_fifo_n265), 
	.A(FE_PHN4278_U_dfifo_U_dcore_U_sub_fifo_n265));
   BUF_X32 FE_PHC2345_U_dfifo_U_dcore_U_sub_fifo_n290 (.Z(FE_PHN2345_U_dfifo_U_dcore_U_sub_fifo_n290), 
	.A(FE_PHN4206_U_dfifo_U_dcore_U_sub_fifo_n290));
   BUF_X32 FE_PHC2344_U_dfifo_U_dcore_U_sub_fifo_n258 (.Z(FE_PHN2344_U_dfifo_U_dcore_U_sub_fifo_n258), 
	.A(FE_PHN4310_U_dfifo_U_dcore_U_sub_fifo_n258));
   BUF_X32 FE_PHC2343_U_afifo_U_acore_U_sub_fifo_n205 (.Z(FE_PHN2343_U_afifo_U_acore_U_sub_fifo_n205), 
	.A(FE_PHN5058_U_afifo_U_acore_U_sub_fifo_n205));
   BUF_X32 FE_PHC2342_U_dfifo_U_dcore_U_sub_fifo_n255 (.Z(FE_PHN2342_U_dfifo_U_dcore_U_sub_fifo_n255), 
	.A(FE_PHN5036_U_dfifo_U_dcore_U_sub_fifo_n255));
   BUF_X32 FE_PHC2341_U_dfifo_U_dcore_U_sub_fifo_n254 (.Z(FE_PHN2341_U_dfifo_U_dcore_U_sub_fifo_n254), 
	.A(FE_PHN5051_U_dfifo_U_dcore_U_sub_fifo_n254));
   BUF_X32 FE_PHC2340_U_dfifo_U_dcore_U_sub_fifo_n274 (.Z(FE_PHN2340_U_dfifo_U_dcore_U_sub_fifo_n274), 
	.A(FE_PHN5083_U_dfifo_U_dcore_U_sub_fifo_n274));
   BUF_X32 FE_PHC2339_U_dfifo_U_dcore_U_sub_fifo_n267 (.Z(FE_PHN2339_U_dfifo_U_dcore_U_sub_fifo_n267), 
	.A(FE_PHN4925_U_dfifo_U_dcore_U_sub_fifo_n267));
   BUF_X32 FE_PHC2338_U_dfifo_U_dcore_U_sub_fifo_n277 (.Z(FE_PHN2338_U_dfifo_U_dcore_U_sub_fifo_n277), 
	.A(FE_PHN4268_U_dfifo_U_dcore_U_sub_fifo_n277));
   BUF_X32 FE_PHC2337_U_dfifo_U_dcore_U_sub_fifo_n286 (.Z(FE_PHN2337_U_dfifo_U_dcore_U_sub_fifo_n286), 
	.A(FE_PHN4241_U_dfifo_U_dcore_U_sub_fifo_n286));
   BUF_X32 FE_PHC2336_U_dfifo_U_dcore_U_sub_fifo_n276 (.Z(FE_PHN2336_U_dfifo_U_dcore_U_sub_fifo_n276), 
	.A(FE_PHN4296_U_dfifo_U_dcore_U_sub_fifo_n276));
   BUF_X32 FE_PHC2335_U_dfifo_U_dcore_U_sub_fifo_n262 (.Z(FE_PHN2335_U_dfifo_U_dcore_U_sub_fifo_n262), 
	.A(FE_PHN4341_U_dfifo_U_dcore_U_sub_fifo_n262));
   BUF_X32 FE_PHC2334_U_dfifo_U_dcore_U_sub_fifo_n246 (.Z(FE_PHN2334_U_dfifo_U_dcore_U_sub_fifo_n246), 
	.A(FE_PHN4183_U_dfifo_U_dcore_U_sub_fifo_n246));
   BUF_X32 FE_PHC2332_U_dfifo_U_dcore_U_sub_fifo_n249 (.Z(FE_PHN2332_U_dfifo_U_dcore_U_sub_fifo_n249), 
	.A(FE_PHN4189_U_dfifo_U_dcore_U_sub_fifo_n249));
   BUF_X32 FE_PHC2331_U_dfifo_U_dcore_U_sub_fifo_n248 (.Z(FE_PHN2331_U_dfifo_U_dcore_U_sub_fifo_n248), 
	.A(FE_PHN4250_U_dfifo_U_dcore_U_sub_fifo_n248));
   BUF_X32 FE_PHC2329_U_dfifo_U_dcore_U_sub_fifo_n282 (.Z(FE_PHN2329_U_dfifo_U_dcore_U_sub_fifo_n282), 
	.A(FE_PHN4254_U_dfifo_U_dcore_U_sub_fifo_n282));
   BUF_X32 FE_PHC2328_U_afifo_U_acore_U_sub_fifo_n301 (.Z(FE_PHN2328_U_afifo_U_acore_U_sub_fifo_n301), 
	.A(U_afifo_U_acore_U_sub_fifo_n301));
   BUF_X32 FE_PHC2327_U_dfifo_U_dcore_U_sub_fifo_n299 (.Z(FE_PHN2327_U_dfifo_U_dcore_U_sub_fifo_n299), 
	.A(FE_PHN5157_U_dfifo_U_dcore_U_sub_fifo_n299));
   BUF_X32 FE_PHC2326_U_dfifo_U_dcore_U_sub_fifo_n256 (.Z(FE_PHN2326_U_dfifo_U_dcore_U_sub_fifo_n256), 
	.A(FE_PHN4881_U_dfifo_U_dcore_U_sub_fifo_n256));
   BUF_X32 FE_PHC2325_U_dfifo_U_dcore_U_sub_fifo_n263 (.Z(FE_PHN2325_U_dfifo_U_dcore_U_sub_fifo_n263), 
	.A(FE_PHN5072_U_dfifo_U_dcore_U_sub_fifo_n263));
   BUF_X32 FE_PHC2324_U_afifo_U_acore_U_sub_fifo_n265 (.Z(FE_PHN2324_U_afifo_U_acore_U_sub_fifo_n265), 
	.A(FE_PHN5087_U_afifo_U_acore_U_sub_fifo_n265));
   BUF_X32 FE_PHC2323_U_dfifo_U_dcore_U_sub_fifo_n250 (.Z(FE_PHN2323_U_dfifo_U_dcore_U_sub_fifo_n250), 
	.A(FE_PHN4251_U_dfifo_U_dcore_U_sub_fifo_n250));
   BUF_X32 FE_PHC2322_U_dfifo_U_dcore_U_sub_fifo_n302 (.Z(FE_PHN2322_U_dfifo_U_dcore_U_sub_fifo_n302), 
	.A(FE_PHN4998_U_dfifo_U_dcore_U_sub_fifo_n302));
   BUF_X32 FE_PHC2321_U_afifo_U_acore_U_sub_fifo_n257 (.Z(FE_PHN2321_U_afifo_U_acore_U_sub_fifo_n257), 
	.A(FE_PHN4030_U_afifo_U_acore_U_sub_fifo_n257));
   BUF_X32 FE_PHC2320_U_dfifo_U_dcore_U_sub_fifo_n243 (.Z(FE_PHN2320_U_dfifo_U_dcore_U_sub_fifo_n243), 
	.A(FE_PHN4256_U_dfifo_U_dcore_U_sub_fifo_n243));
   BUF_X32 FE_PHC2319_U_dfifo_U_dcore_U_sub_fifo_n261 (.Z(FE_PHN2319_U_dfifo_U_dcore_U_sub_fifo_n261), 
	.A(FE_PHN4948_U_dfifo_U_dcore_U_sub_fifo_n261));
   BUF_X32 FE_PHC2318_U_dfifo_U_dcore_U_sub_fifo_n259 (.Z(FE_PHN2318_U_dfifo_U_dcore_U_sub_fifo_n259), 
	.A(FE_PHN5147_U_dfifo_U_dcore_U_sub_fifo_n259));
   BUF_X32 FE_PHC2317_U_dfifo_U_dcore_U_sub_fifo_n284 (.Z(FE_PHN2317_U_dfifo_U_dcore_U_sub_fifo_n284), 
	.A(FE_PHN4238_U_dfifo_U_dcore_U_sub_fifo_n284));
   BUF_X32 FE_PHC2316_U_afifo_U_acore_U_sub_fifo_n302 (.Z(FE_PHN2316_U_afifo_U_acore_U_sub_fifo_n302), 
	.A(U_afifo_U_acore_U_sub_fifo_n302));
   BUF_X32 FE_PHC2315_U_afifo_U_acore_U_sub_fifo_n279 (.Z(FE_PHN2315_U_afifo_U_acore_U_sub_fifo_n279), 
	.A(FE_PHN4226_U_afifo_U_acore_U_sub_fifo_n279));
   BUF_X32 FE_PHC2314_U_dfifo_U_dcore_U_sub_fifo_n289 (.Z(FE_PHN2314_U_dfifo_U_dcore_U_sub_fifo_n289), 
	.A(FE_PHN4091_U_dfifo_U_dcore_U_sub_fifo_n289));
   BUF_X32 FE_PHC2313_U_dfifo_U_dcore_U_sub_fifo_n287 (.Z(FE_PHN2313_U_dfifo_U_dcore_U_sub_fifo_n287), 
	.A(FE_PHN5092_U_dfifo_U_dcore_U_sub_fifo_n287));
   BUF_X32 FE_PHC2312_U_afifo_U_acore_U_sub_fifo_n306 (.Z(FE_PHN2312_U_afifo_U_acore_U_sub_fifo_n306), 
	.A(U_afifo_U_acore_U_sub_fifo_n306));
   BUF_X32 FE_PHC2311_U_dfifo_U_dcore_U_sub_fifo_n298 (.Z(FE_PHN2311_U_dfifo_U_dcore_U_sub_fifo_n298), 
	.A(FE_PHN4843_U_dfifo_U_dcore_U_sub_fifo_n298));
   BUF_X32 FE_PHC2310_U_dfifo_U_dcore_U_sub_fifo_n266 (.Z(FE_PHN2310_U_dfifo_U_dcore_U_sub_fifo_n266), 
	.A(FE_PHN4968_U_dfifo_U_dcore_U_sub_fifo_n266));
   BUF_X32 FE_PHC2309_U_dfifo_U_dcore_U_sub_fifo_n245 (.Z(FE_PHN2309_U_dfifo_U_dcore_U_sub_fifo_n245), 
	.A(FE_PHN4208_U_dfifo_U_dcore_U_sub_fifo_n245));
   BUF_X32 FE_PHC2308_U_afifo_U_acore_U_sub_fifo_n259 (.Z(FE_PHN2308_U_afifo_U_acore_U_sub_fifo_n259), 
	.A(FE_PHN4038_U_afifo_U_acore_U_sub_fifo_n259));
   BUF_X32 FE_PHC2307_U_dfifo_U_dcore_U_sub_fifo_n310 (.Z(FE_PHN2307_U_dfifo_U_dcore_U_sub_fifo_n310), 
	.A(FE_PHN5109_U_dfifo_U_dcore_U_sub_fifo_n310));
   BUF_X32 FE_PHC2306_U_dfifo_U_dcore_U_sub_fifo_n300 (.Z(FE_PHN2306_U_dfifo_U_dcore_U_sub_fifo_n300), 
	.A(FE_PHN4242_U_dfifo_U_dcore_U_sub_fifo_n300));
   BUF_X32 FE_PHC2305_U_dfifo_U_dcore_U_sub_fifo_n244 (.Z(FE_PHN2305_U_dfifo_U_dcore_U_sub_fifo_n244), 
	.A(FE_PHN4063_U_dfifo_U_dcore_U_sub_fifo_n244));
   BUF_X32 FE_PHC2304_U_dfifo_U_dcore_U_sub_fifo_n273 (.Z(FE_PHN2304_U_dfifo_U_dcore_U_sub_fifo_n273), 
	.A(FE_PHN4239_U_dfifo_U_dcore_U_sub_fifo_n273));
   BUF_X32 FE_PHC2303_U_dfifo_U_dcore_U_sub_fifo_n301 (.Z(FE_PHN2303_U_dfifo_U_dcore_U_sub_fifo_n301), 
	.A(FE_PHN4068_U_dfifo_U_dcore_U_sub_fifo_n301));
   BUF_X32 FE_PHC2301_U_dfifo_U_dcore_U_sub_fifo_n296 (.Z(FE_PHN2301_U_dfifo_U_dcore_U_sub_fifo_n296), 
	.A(FE_PHN4918_U_dfifo_U_dcore_U_sub_fifo_n296));
   BUF_X32 FE_PHC2299_U_dfifo_U_dcore_U_sub_fifo_n304 (.Z(FE_PHN2299_U_dfifo_U_dcore_U_sub_fifo_n304), 
	.A(FE_PHN5030_U_dfifo_U_dcore_U_sub_fifo_n304));
   BUF_X32 FE_PHC2298_U_dfifo_U_dcore_U_sub_fifo_n293 (.Z(FE_PHN2298_U_dfifo_U_dcore_U_sub_fifo_n293), 
	.A(FE_PHN4224_U_dfifo_U_dcore_U_sub_fifo_n293));
   BUF_X32 FE_PHC2297_U_dfifo_U_dcore_U_sub_fifo_n308 (.Z(FE_PHN2297_U_dfifo_U_dcore_U_sub_fifo_n308), 
	.A(FE_PHN5070_U_dfifo_U_dcore_U_sub_fifo_n308));
   BUF_X32 FE_PHC2296_U_dfifo_U_dcore_U_sub_fifo_n247 (.Z(FE_PHN2296_U_dfifo_U_dcore_U_sub_fifo_n247), 
	.A(FE_PHN5116_U_dfifo_U_dcore_U_sub_fifo_n247));
   BUF_X32 FE_PHC2295_U_afifo_U_acore_U_sub_fifo_n173 (.Z(FE_PHN2295_U_afifo_U_acore_U_sub_fifo_n173), 
	.A(FE_PHN4979_U_afifo_U_acore_U_sub_fifo_n173));
   BUF_X32 FE_PHC2293_U_dfifo_U_dcore_U_sub_fifo_n252 (.Z(FE_PHN2293_U_dfifo_U_dcore_U_sub_fifo_n252), 
	.A(FE_PHN4007_U_dfifo_U_dcore_U_sub_fifo_n252));
   BUF_X32 FE_PHC2292_U_afifo_U_acore_U_sub_fifo_n180 (.Z(FE_PHN2292_U_afifo_U_acore_U_sub_fifo_n180), 
	.A(FE_PHN5073_U_afifo_U_acore_U_sub_fifo_n180));
   BUF_X32 FE_PHC2291_U_dfifo_U_dcore_U_sub_fifo_n280 (.Z(FE_PHN2291_U_dfifo_U_dcore_U_sub_fifo_n280), 
	.A(FE_PHN5082_U_dfifo_U_dcore_U_sub_fifo_n280));
   BUF_X32 FE_PHC2290_U_afifo_U_acore_U_sub_fifo_n210 (.Z(FE_PHN2290_U_afifo_U_acore_U_sub_fifo_n210), 
	.A(FE_PHN4987_U_afifo_U_acore_U_sub_fifo_n210));
   BUF_X32 FE_PHC2289_U_dfifo_U_dcore_U_sub_fifo_n288 (.Z(FE_PHN2289_U_dfifo_U_dcore_U_sub_fifo_n288), 
	.A(FE_PHN4209_U_dfifo_U_dcore_U_sub_fifo_n288));
   BUF_X32 FE_PHC2288_U_dfifo_U_dcore_U_sub_fifo_n251 (.Z(FE_PHN2288_U_dfifo_U_dcore_U_sub_fifo_n251), 
	.A(FE_PHN5128_U_dfifo_U_dcore_U_sub_fifo_n251));
   BUF_X32 FE_PHC2287_U_afifo_U_acore_U_sub_fifo_n194 (.Z(FE_PHN2287_U_afifo_U_acore_U_sub_fifo_n194), 
	.A(FE_PHN5095_U_afifo_U_acore_U_sub_fifo_n194));
   BUF_X32 FE_PHC2285_U_dfifo_U_dcore_U_sub_fifo_n281 (.Z(FE_PHN2285_U_dfifo_U_dcore_U_sub_fifo_n281), 
	.A(FE_PHN5033_U_dfifo_U_dcore_U_sub_fifo_n281));
   BUF_X32 FE_PHC2284_U_dfifo_U_dcore_U_sub_fifo_n291 (.Z(FE_PHN2284_U_dfifo_U_dcore_U_sub_fifo_n291), 
	.A(FE_PHN4961_U_dfifo_U_dcore_U_sub_fifo_n291));
   BUF_X32 FE_PHC2283_U_dfifo_U_dcore_U_sub_fifo_n297 (.Z(FE_PHN2283_U_dfifo_U_dcore_U_sub_fifo_n297), 
	.A(FE_PHN5062_U_dfifo_U_dcore_U_sub_fifo_n297));
   BUF_X32 FE_PHC2282_U_afifo_U_acore_U_sub_fifo_n224 (.Z(FE_PHN2282_U_afifo_U_acore_U_sub_fifo_n224), 
	.A(FE_PHN4071_U_afifo_U_acore_U_sub_fifo_n224));
   BUF_X32 FE_PHC2281_U_afifo_U_acore_U_sub_fifo_n213 (.Z(FE_PHN2281_U_afifo_U_acore_U_sub_fifo_n213), 
	.A(FE_PHN5075_U_afifo_U_acore_U_sub_fifo_n213));
   BUF_X32 FE_PHC2280_U_dfifo_U_dcore_U_sub_fifo_n285 (.Z(FE_PHN2280_U_dfifo_U_dcore_U_sub_fifo_n285), 
	.A(FE_PHN5057_U_dfifo_U_dcore_U_sub_fifo_n285));
   BUF_X32 FE_PHC2279_U_afifo_U_acore_U_sub_fifo_n211 (.Z(FE_PHN2279_U_afifo_U_acore_U_sub_fifo_n211), 
	.A(FE_PHN4016_U_afifo_U_acore_U_sub_fifo_n211));
   BUF_X32 FE_PHC2278_U_afifo_U_acore_U_sub_fifo_n177 (.Z(FE_PHN2278_U_afifo_U_acore_U_sub_fifo_n177), 
	.A(FE_PHN5101_U_afifo_U_acore_U_sub_fifo_n177));
   BUF_X32 FE_PHC2277_U_afifo_U_acore_U_sub_fifo_n226 (.Z(FE_PHN2277_U_afifo_U_acore_U_sub_fifo_n226), 
	.A(FE_PHN3492_U_afifo_U_acore_U_sub_fifo_n226));
   BUF_X32 FE_PHC2276_U_afifo_U_acore_U_sub_fifo_n253 (.Z(FE_PHN2276_U_afifo_U_acore_U_sub_fifo_n253), 
	.A(FE_PHN3493_U_afifo_U_acore_U_sub_fifo_n253));
   BUF_X32 FE_PHC2275_U_afifo_U_acore_U_sub_fifo_n200 (.Z(FE_PHN2275_U_afifo_U_acore_U_sub_fifo_n200), 
	.A(FE_PHN3300_U_afifo_U_acore_U_sub_fifo_n200));
   BUF_X32 FE_PHC2274_U_afifo_U_acore_U_sub_fifo_n243 (.Z(FE_PHN2274_U_afifo_U_acore_U_sub_fifo_n243), 
	.A(FE_PHN5068_U_afifo_U_acore_U_sub_fifo_n243));
   BUF_X32 FE_PHC2273_U_afifo_U_acore_U_sub_fifo_n245 (.Z(FE_PHN2273_U_afifo_U_acore_U_sub_fifo_n245), 
	.A(FE_PHN5140_U_afifo_U_acore_U_sub_fifo_n245));
   BUF_X32 FE_PHC2272_U_afifo_U_acore_U_sub_fifo_n215 (.Z(FE_PHN2272_U_afifo_U_acore_U_sub_fifo_n215), 
	.A(FE_PHN4056_U_afifo_U_acore_U_sub_fifo_n215));
   BUF_X32 FE_PHC2271_U_afifo_U_acore_U_sub_fifo_n300 (.Z(FE_PHN2271_U_afifo_U_acore_U_sub_fifo_n300), 
	.A(U_afifo_U_acore_U_sub_fifo_n300));
   BUF_X32 FE_PHC2269_U_afifo_U_acore_U_sub_fifo_n252 (.Z(FE_PHN2269_U_afifo_U_acore_U_sub_fifo_n252), 
	.A(FE_PHN3488_U_afifo_U_acore_U_sub_fifo_n252));
   BUF_X32 FE_PHC2268_U_afifo_U_acore_U_sub_fifo_n256 (.Z(FE_PHN2268_U_afifo_U_acore_U_sub_fifo_n256), 
	.A(FE_PHN4899_U_afifo_U_acore_U_sub_fifo_n256));
   BUF_X32 FE_PHC2267_U_afifo_U_acore_U_sub_fifo_n249 (.Z(FE_PHN2267_U_afifo_U_acore_U_sub_fifo_n249), 
	.A(FE_PHN5154_U_afifo_U_acore_U_sub_fifo_n249));
   BUF_X32 FE_PHC2266_U_afifo_U_acore_U_sub_fifo_n203 (.Z(FE_PHN2266_U_afifo_U_acore_U_sub_fifo_n203), 
	.A(FE_PHN4965_U_afifo_U_acore_U_sub_fifo_n203));
   BUF_X32 FE_PHC2265_U_afifo_U_acore_U_sub_fifo_n319 (.Z(FE_PHN2265_U_afifo_U_acore_U_sub_fifo_n319), 
	.A(U_afifo_U_acore_U_sub_fifo_n319));
   BUF_X32 FE_PHC2264_U_afifo_U_acore_U_sub_fifo_n179 (.Z(FE_PHN2264_U_afifo_U_acore_U_sub_fifo_n179), 
	.A(FE_PHN3997_U_afifo_U_acore_U_sub_fifo_n179));
   BUF_X32 FE_PHC2263_U_afifo_U_acore_U_sub_fifo_n191 (.Z(FE_PHN2263_U_afifo_U_acore_U_sub_fifo_n191), 
	.A(FE_PHN5022_U_afifo_U_acore_U_sub_fifo_n191));
   BUF_X32 FE_PHC2262_U_afifo_U_acore_U_sub_fifo_n183 (.Z(FE_PHN2262_U_afifo_U_acore_U_sub_fifo_n183), 
	.A(FE_PHN4015_U_afifo_U_acore_U_sub_fifo_n183));
   BUF_X32 FE_PHC2261_U_afifo_U_acore_U_sub_fifo_n283 (.Z(FE_PHN2261_U_afifo_U_acore_U_sub_fifo_n283), 
	.A(FE_PHN5003_U_afifo_U_acore_U_sub_fifo_n283));
   BUF_X32 FE_PHC2260_U_afifo_U_acore_U_sub_fifo_n227 (.Z(FE_PHN2260_U_afifo_U_acore_U_sub_fifo_n227), 
	.A(FE_PHN5063_U_afifo_U_acore_U_sub_fifo_n227));
   BUF_X32 FE_PHC2259_U_afifo_U_acore_U_sub_fifo_n289 (.Z(FE_PHN2259_U_afifo_U_acore_U_sub_fifo_n289), 
	.A(FE_PHN3980_U_afifo_U_acore_U_sub_fifo_n289));
   BUF_X32 FE_PHC2258_U_afifo_U_acore_U_sub_fifo_n198 (.Z(FE_PHN2258_U_afifo_U_acore_U_sub_fifo_n198), 
	.A(FE_PHN3296_U_afifo_U_acore_U_sub_fifo_n198));
   BUF_X32 FE_PHC2257_U_afifo_U_acore_U_sub_fifo_n284 (.Z(FE_PHN2257_U_afifo_U_acore_U_sub_fifo_n284), 
	.A(FE_PHN4097_U_afifo_U_acore_U_sub_fifo_n284));
   BUF_X32 FE_PHC2256_U_afifo_U_acore_U_sub_fifo_n237 (.Z(FE_PHN2256_U_afifo_U_acore_U_sub_fifo_n237), 
	.A(FE_PHN5040_U_afifo_U_acore_U_sub_fifo_n237));
   BUF_X32 FE_PHC2255_U_afifo_U_acore_U_sub_fifo_n228 (.Z(FE_PHN2255_U_afifo_U_acore_U_sub_fifo_n228), 
	.A(FE_PHN3966_U_afifo_U_acore_U_sub_fifo_n228));
   BUF_X32 FE_PHC2253_U_afifo_U_acore_U_sub_fifo_n186 (.Z(FE_PHN2253_U_afifo_U_acore_U_sub_fifo_n186), 
	.A(FE_PHN3957_U_afifo_U_acore_U_sub_fifo_n186));
   BUF_X32 FE_PHC2252_U_afifo_U_acore_U_sub_fifo_n246 (.Z(FE_PHN2252_U_afifo_U_acore_U_sub_fifo_n246), 
	.A(FE_PHN5078_U_afifo_U_acore_U_sub_fifo_n246));
   BUF_X32 FE_PHC2251_U_afifo_U_acore_U_sub_fifo_n199 (.Z(FE_PHN2251_U_afifo_U_acore_U_sub_fifo_n199), 
	.A(FE_PHN3487_U_afifo_U_acore_U_sub_fifo_n199));
   BUF_X32 FE_PHC2250_U_afifo_U_acore_U_sub_fifo_n234 (.Z(FE_PHN2250_U_afifo_U_acore_U_sub_fifo_n234), 
	.A(FE_PHN3953_U_afifo_U_acore_U_sub_fifo_n234));
   BUF_X32 FE_PHC2249_U_afifo_U_acore_U_sub_fifo_n258 (.Z(FE_PHN2249_U_afifo_U_acore_U_sub_fifo_n258), 
	.A(FE_PHN4942_U_afifo_U_acore_U_sub_fifo_n258));
   BUF_X32 FE_PHC2248_U_afifo_U_acore_U_sub_fifo_n189 (.Z(FE_PHN2248_U_afifo_U_acore_U_sub_fifo_n189), 
	.A(FE_PHN3991_U_afifo_U_acore_U_sub_fifo_n189));
   BUF_X32 FE_PHC2247_U_afifo_U_acore_U_sub_fifo_n204 (.Z(FE_PHN2247_U_afifo_U_acore_U_sub_fifo_n204), 
	.A(FE_PHN3996_U_afifo_U_acore_U_sub_fifo_n204));
   BUF_X32 FE_PHC2246_U_afifo_U_acore_U_sub_fifo_n254 (.Z(FE_PHN2246_U_afifo_U_acore_U_sub_fifo_n254), 
	.A(FE_PHN3993_U_afifo_U_acore_U_sub_fifo_n254));
   BUF_X32 FE_PHC2244_U_afifo_U_acore_U_sub_fifo_n276 (.Z(FE_PHN2244_U_afifo_U_acore_U_sub_fifo_n276), 
	.A(U_afifo_U_acore_U_sub_fifo_n276));
   BUF_X32 FE_PHC2243_U_afifo_U_acore_U_sub_fifo_n241 (.Z(FE_PHN2243_U_afifo_U_acore_U_sub_fifo_n241), 
	.A(FE_PHN3929_U_afifo_U_acore_U_sub_fifo_n241));
   BUF_X32 FE_PHC2242_U_afifo_U_acore_U_sub_fifo_n185 (.Z(FE_PHN2242_U_afifo_U_acore_U_sub_fifo_n185), 
	.A(FE_PHN5069_U_afifo_U_acore_U_sub_fifo_n185));
   BUF_X32 FE_PHC2239_U_afifo_U_acore_U_sub_fifo_n235 (.Z(FE_PHN2239_U_afifo_U_acore_U_sub_fifo_n235), 
	.A(FE_PHN4992_U_afifo_U_acore_U_sub_fifo_n235));
   BUF_X32 FE_PHC2238_U_afifo_U_acore_U_sub_fifo_n286 (.Z(FE_PHN2238_U_afifo_U_acore_U_sub_fifo_n286), 
	.A(FE_PHN3952_U_afifo_U_acore_U_sub_fifo_n286));
   BUF_X32 FE_PHC2237_U_afifo_U_acore_U_sub_fifo_n231 (.Z(FE_PHN2237_U_afifo_U_acore_U_sub_fifo_n231), 
	.A(FE_PHN5079_U_afifo_U_acore_U_sub_fifo_n231));
   BUF_X32 FE_PHC2236_U_afifo_U_acore_U_sub_fifo_n192 (.Z(FE_PHN2236_U_afifo_U_acore_U_sub_fifo_n192), 
	.A(FE_PHN5032_U_afifo_U_acore_U_sub_fifo_n192));
   BUF_X32 FE_PHC2235_U_dfifo_U_dcore_U_sub_fifo_n396 (.Z(FE_PHN2235_U_dfifo_U_dcore_U_sub_fifo_n396), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n396));
   BUF_X32 FE_PHC2234_U_afifo_U_acore_U_sub_fifo_n181 (.Z(FE_PHN2234_U_afifo_U_acore_U_sub_fifo_n181), 
	.A(FE_PHN4070_U_afifo_U_acore_U_sub_fifo_n181));
   BUF_X32 FE_PHC2231_U_afifo_U_acore_U_sub_fifo_n182 (.Z(FE_PHN2231_U_afifo_U_acore_U_sub_fifo_n182), 
	.A(FE_PHN4010_U_afifo_U_acore_U_sub_fifo_n182));
   BUF_X32 FE_PHC2230_U_afifo_U_acore_U_sub_fifo_n232 (.Z(FE_PHN2230_U_afifo_U_acore_U_sub_fifo_n232), 
	.A(FE_PHN4074_U_afifo_U_acore_U_sub_fifo_n232));
   BUF_X32 FE_PHC2229_U_dfifo_U_dcore_U_sub_fifo_n374 (.Z(FE_PHN2229_U_dfifo_U_dcore_U_sub_fifo_n374), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n374));
   BUF_X32 FE_PHC2228_U_afifo_U_acore_U_sub_fifo_n290 (.Z(FE_PHN2228_U_afifo_U_acore_U_sub_fifo_n290), 
	.A(FE_PHN4055_U_afifo_U_acore_U_sub_fifo_n290));
   BUF_X32 FE_PHC2227_U_afifo_U_acore_U_sub_fifo_n190 (.Z(FE_PHN2227_U_afifo_U_acore_U_sub_fifo_n190), 
	.A(FE_PHN4107_U_afifo_U_acore_U_sub_fifo_n190));
   BUF_X32 FE_PHC2226_U_afifo_U_acore_U_sub_fifo_n288 (.Z(FE_PHN2226_U_afifo_U_acore_U_sub_fifo_n288), 
	.A(FE_PHN4092_U_afifo_U_acore_U_sub_fifo_n288));
   BUF_X32 FE_PHC2222_U_dfifo_U_dcore_U_sub_fifo_n376 (.Z(FE_PHN2222_U_dfifo_U_dcore_U_sub_fifo_n376), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n376));
   BUF_X32 FE_PHC2221_U_dfifo_U_dcore_U_sub_fifo_n350 (.Z(FE_PHN2221_U_dfifo_U_dcore_U_sub_fifo_n350), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n350));
   BUF_X32 FE_PHC2220_U_dfifo_U_dcore_U_sub_fifo_n430 (.Z(FE_PHN2220_U_dfifo_U_dcore_U_sub_fifo_n430), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n430));
   BUF_X32 FE_PHC2218_U_dfifo_U_dcore_U_sub_fifo_n422 (.Z(FE_PHN2218_U_dfifo_U_dcore_U_sub_fifo_n422), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n422));
   BUF_X32 FE_PHC2217_U_dfifo_U_dcore_U_sub_fifo_n381 (.Z(FE_PHN2217_U_dfifo_U_dcore_U_sub_fifo_n381), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n381));
   BUF_X32 FE_PHC2216_U_dfifo_U_dcore_U_sub_fifo_n337 (.Z(FE_PHN2216_U_dfifo_U_dcore_U_sub_fifo_n337), 
	.A(FE_PHN3829_U_dfifo_U_dcore_U_sub_fifo_n337));
   BUF_X32 FE_PHC2214_U_dfifo_U_dcore_U_sub_fifo_n388 (.Z(FE_PHN2214_U_dfifo_U_dcore_U_sub_fifo_n388), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n388));
   BUF_X32 FE_PHC2213_U_dfifo_U_dcore_U_sub_fifo_n427 (.Z(FE_PHN2213_U_dfifo_U_dcore_U_sub_fifo_n427), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n427));
   BUF_X32 FE_PHC2211_U_dfifo_U_dcore_U_sub_fifo_n386 (.Z(FE_PHN2211_U_dfifo_U_dcore_U_sub_fifo_n386), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n386));
   BUF_X32 FE_PHC2209_U_dfifo_U_dcore_U_sub_fifo_n368 (.Z(FE_PHN2209_U_dfifo_U_dcore_U_sub_fifo_n368), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n368));
   BUF_X32 FE_PHC2208_U_dfifo_U_dcore_U_sub_fifo_n445 (.Z(FE_PHN2208_U_dfifo_U_dcore_U_sub_fifo_n445), 
	.A(FE_PHN4824_U_dfifo_U_dcore_U_sub_fifo_n445));
   BUF_X32 FE_PHC2207_U_dfifo_U_dcore_U_sub_fifo_n387 (.Z(FE_PHN2207_U_dfifo_U_dcore_U_sub_fifo_n387), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n387));
   BUF_X32 FE_PHC2206_U_dfifo_U_dcore_U_sub_fifo_n432 (.Z(FE_PHN2206_U_dfifo_U_dcore_U_sub_fifo_n432), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n432));
   BUF_X32 FE_PHC2205_U_dfifo_U_dcore_U_sub_fifo_n314 (.Z(FE_PHN2205_U_dfifo_U_dcore_U_sub_fifo_n314), 
	.A(FE_PHN4889_U_dfifo_U_dcore_U_sub_fifo_n314));
   BUF_X32 FE_PHC2204_U_dfifo_U_dcore_U_sub_fifo_n394 (.Z(FE_PHN2204_U_dfifo_U_dcore_U_sub_fifo_n394), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n394));
   BUF_X32 FE_PHC2203_U_dfifo_U_dcore_U_sub_fifo_n435 (.Z(FE_PHN2203_U_dfifo_U_dcore_U_sub_fifo_n435), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n435));
   BUF_X32 FE_PHC2202_U_dfifo_U_dcore_U_sub_fifo_n373 (.Z(FE_PHN2202_U_dfifo_U_dcore_U_sub_fifo_n373), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n373));
   BUF_X32 FE_PHC2201_U_dfifo_U_dcore_U_sub_fifo_n434 (.Z(FE_PHN2201_U_dfifo_U_dcore_U_sub_fifo_n434), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n434));
   BUF_X32 FE_PHC2199_U_dfifo_U_dcore_U_sub_fifo_n423 (.Z(FE_PHN2199_U_dfifo_U_dcore_U_sub_fifo_n423), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n423));
   BUF_X32 FE_PHC2198_U_dfifo_U_dcore_U_sub_fifo_n433 (.Z(FE_PHN2198_U_dfifo_U_dcore_U_sub_fifo_n433), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n433));
   BUF_X32 FE_PHC2197_U_dfifo_U_dcore_U_sub_fifo_n426 (.Z(FE_PHN2197_U_dfifo_U_dcore_U_sub_fifo_n426), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n426));
   BUF_X32 FE_PHC2195_U_dfifo_U_dcore_U_sub_fifo_n428 (.Z(FE_PHN2195_U_dfifo_U_dcore_U_sub_fifo_n428), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n428));
   BUF_X32 FE_PHC2194_U_dfifo_U_dcore_U_sub_fifo_n437 (.Z(FE_PHN2194_U_dfifo_U_dcore_U_sub_fifo_n437), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n437));
   BUF_X32 FE_PHC2193_U_dfifo_U_dcore_U_sub_fifo_n421 (.Z(FE_PHN2193_U_dfifo_U_dcore_U_sub_fifo_n421), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n421));
   BUF_X32 FE_PHC2192_U_dfifo_U_dcore_U_sub_fifo_n384 (.Z(FE_PHN2192_U_dfifo_U_dcore_U_sub_fifo_n384), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n384));
   BUF_X32 FE_PHC2191_U_dfifo_U_dcore_U_sub_fifo_n436 (.Z(FE_PHN2191_U_dfifo_U_dcore_U_sub_fifo_n436), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n436));
   BUF_X32 FE_PHC2190_U_dfifo_U_dcore_U_sub_fifo_n379 (.Z(FE_PHN2190_U_dfifo_U_dcore_U_sub_fifo_n379), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n379));
   BUF_X32 FE_PHC2188_U_dfifo_U_dcore_U_sub_fifo_n385 (.Z(FE_PHN2188_U_dfifo_U_dcore_U_sub_fifo_n385), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n385));
   BUF_X32 FE_PHC2186_U_dfifo_U_dcore_U_sub_fifo_n431 (.Z(FE_PHN2186_U_dfifo_U_dcore_U_sub_fifo_n431), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n431));
   BUF_X32 FE_PHC2185_U_dfifo_U_dcore_U_sub_fifo_n380 (.Z(FE_PHN2185_U_dfifo_U_dcore_U_sub_fifo_n380), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n380));
   BUF_X32 FE_PHC2184_U_dfifo_U_dcore_U_sub_fifo_n366 (.Z(FE_PHN2184_U_dfifo_U_dcore_U_sub_fifo_n366), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n366));
   BUF_X32 FE_PHC2183_U_dfifo_U_dcore_U_sub_fifo_n429 (.Z(FE_PHN2183_U_dfifo_U_dcore_U_sub_fifo_n429), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n429));
   BUF_X32 FE_PHC2182_U_dfifo_U_dcore_U_sub_fifo_n365 (.Z(FE_PHN2182_U_dfifo_U_dcore_U_sub_fifo_n365), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n365));
   BUF_X32 FE_PHC2178_U_dfifo_U_dcore_U_sub_fifo_n382 (.Z(FE_PHN2178_U_dfifo_U_dcore_U_sub_fifo_n382), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n382));
   BUF_X32 FE_PHC2177_U_dfifo_U_dcore_U_sub_fifo_n424 (.Z(FE_PHN2177_U_dfifo_U_dcore_U_sub_fifo_n424), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n424));
   BUF_X32 FE_PHC2176_U_dfifo_U_dcore_U_sub_fifo_n389 (.Z(FE_PHN2176_U_dfifo_U_dcore_U_sub_fifo_n389), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n389));
   BUF_X32 FE_PHC2175_U_dfifo_U_dcore_U_sub_fifo_n317 (.Z(FE_PHN2175_U_dfifo_U_dcore_U_sub_fifo_n317), 
	.A(FE_PHN3788_U_dfifo_U_dcore_U_sub_fifo_n317));
   BUF_X32 FE_PHC2174_U_dfifo_U_dcore_U_sub_fifo_n390 (.Z(FE_PHN2174_U_dfifo_U_dcore_U_sub_fifo_n390), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n390));
   BUF_X32 FE_PHC2173_U_dfifo_U_dcore_U_sub_fifo_n391 (.Z(FE_PHN2173_U_dfifo_U_dcore_U_sub_fifo_n391), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n391));
   BUF_X32 FE_PHC2172_U_dfifo_U_dcore_U_sub_fifo_n425 (.Z(FE_PHN2172_U_dfifo_U_dcore_U_sub_fifo_n425), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n425));
   BUF_X32 FE_PHC2171_U_dfifo_U_dcore_U_sub_fifo_n419 (.Z(FE_PHN2171_U_dfifo_U_dcore_U_sub_fifo_n419), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n419));
   BUF_X32 FE_PHC2170_U_dfifo_U_dcore_U_sub_fifo_n383 (.Z(FE_PHN2170_U_dfifo_U_dcore_U_sub_fifo_n383), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n383));
   BUF_X32 FE_PHC2169_U_dfifo_U_dcore_U_sub_fifo_n392 (.Z(FE_PHN2169_U_dfifo_U_dcore_U_sub_fifo_n392), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n392));
   BUF_X32 FE_PHC2168_U_dfifo_U_dcore_U_sub_fifo_n393 (.Z(FE_PHN2168_U_dfifo_U_dcore_U_sub_fifo_n393), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n393));
   BUF_X32 FE_PHC2167_U_dfifo_U_dcore_U_sub_fifo_n321 (.Z(FE_PHN2167_U_dfifo_U_dcore_U_sub_fifo_n321), 
	.A(FE_PHN3794_U_dfifo_U_dcore_U_sub_fifo_n321));
   BUF_X32 FE_PHC2165_U_dfifo_U_dcore_U_sub_fifo_n413 (.Z(FE_PHN2165_U_dfifo_U_dcore_U_sub_fifo_n413), 
	.A(FE_PHN4856_U_dfifo_U_dcore_U_sub_fifo_n413));
   BUF_X32 FE_PHC2162_U_dfifo_U_dcore_U_sub_fifo_n395 (.Z(FE_PHN2162_U_dfifo_U_dcore_U_sub_fifo_n395), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n395));
   BUF_X32 FE_PHC2161_U_afifo_f_data2_7_ (.Z(FE_PHN2161_U_afifo_f_data2_7_), 
	.A(U_afifo_f_data2_7_));
   BUF_X32 FE_PHC2160_U_dfifo_U_dcore_U_sub_fifo_n313 (.Z(FE_PHN2160_U_dfifo_U_dcore_U_sub_fifo_n313), 
	.A(FE_PHN3748_U_dfifo_U_dcore_U_sub_fifo_n313));
   BUF_X32 FE_PHC2159_U_dfifo_U_dcore_U_sub_fifo_n363 (.Z(FE_PHN2159_U_dfifo_U_dcore_U_sub_fifo_n363), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n363));
   BUF_X32 FE_PHC2158_U_dfifo_U_dcore_U_sub_fifo_n401 (.Z(FE_PHN2158_U_dfifo_U_dcore_U_sub_fifo_n401), 
	.A(FE_PHN4806_U_dfifo_U_dcore_U_sub_fifo_n401));
   BUF_X32 FE_PHC2155_U_dfifo_U_dcore_U_sub_fifo_n420 (.Z(FE_PHN2155_U_dfifo_U_dcore_U_sub_fifo_n420), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n420));
   BUF_X32 FE_PHC2153_U_dfifo_U_dcore_U_sub_fifo_n416 (.Z(FE_PHN2153_U_dfifo_U_dcore_U_sub_fifo_n416), 
	.A(FE_PHN3752_U_dfifo_U_dcore_U_sub_fifo_n416));
   BUF_X32 FE_PHC2152_U_dfifo_U_dcore_U_sub_fifo_n333 (.Z(FE_PHN2152_U_dfifo_U_dcore_U_sub_fifo_n333), 
	.A(FE_PHN4769_U_dfifo_U_dcore_U_sub_fifo_n333));
   BUF_X32 FE_PHC2151_U_dfifo_U_dcore_U_sub_fifo_n361 (.Z(FE_PHN2151_U_dfifo_U_dcore_U_sub_fifo_n361), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n361));
   BUF_X32 FE_PHC2147_U_dfifo_U_dcore_U_sub_fifo_n443 (.Z(FE_PHN2147_U_dfifo_U_dcore_U_sub_fifo_n443), 
	.A(FE_PHN3727_U_dfifo_U_dcore_U_sub_fifo_n443));
   BUF_X32 FE_PHC2144_U_dfifo_U_dcore_U_sub_fifo_n326 (.Z(FE_PHN2144_U_dfifo_U_dcore_U_sub_fifo_n326), 
	.A(FE_PHN3732_U_dfifo_U_dcore_U_sub_fifo_n326));
   BUF_X32 FE_PHC2142_U_dfifo_U_dcore_U_sub_fifo_n315 (.Z(FE_PHN2142_U_dfifo_U_dcore_U_sub_fifo_n315), 
	.A(FE_PHN3754_U_dfifo_U_dcore_U_sub_fifo_n315));
   BUF_X32 FE_PHC2139_U_dfifo_U_dcore_U_sub_fifo_n405 (.Z(FE_PHN2139_U_dfifo_U_dcore_U_sub_fifo_n405), 
	.A(FE_PHN3711_U_dfifo_U_dcore_U_sub_fifo_n405));
   BUF_X32 FE_PHC2138_U_dfifo_U_dcore_U_sub_fifo_n403 (.Z(FE_PHN2138_U_dfifo_U_dcore_U_sub_fifo_n403), 
	.A(FE_PHN4768_U_dfifo_U_dcore_U_sub_fifo_n403));
   BUF_X32 FE_PHC2137_U_dfifo_U_dcore_U_sub_fifo_n322 (.Z(FE_PHN2137_U_dfifo_U_dcore_U_sub_fifo_n322), 
	.A(FE_PHN3674_U_dfifo_U_dcore_U_sub_fifo_n322));
   BUF_X32 FE_PHC2136_U_dfifo_U_dcore_U_sub_fifo_n411 (.Z(FE_PHN2136_U_dfifo_U_dcore_U_sub_fifo_n411), 
	.A(FE_PHN3721_U_dfifo_U_dcore_U_sub_fifo_n411));
   BUF_X32 FE_PHC2135_U_dfifo_U_dcore_U_sub_fifo_n402 (.Z(FE_PHN2135_U_dfifo_U_dcore_U_sub_fifo_n402), 
	.A(FE_PHN4744_U_dfifo_U_dcore_U_sub_fifo_n402));
   BUF_X32 FE_PHC2134_U_dfifo_U_dcore_U_sub_fifo_n325 (.Z(FE_PHN2134_U_dfifo_U_dcore_U_sub_fifo_n325), 
	.A(FE_PHN3741_U_dfifo_U_dcore_U_sub_fifo_n325));
   BUF_X32 FE_PHC2133_U_afifo_n3 (.Z(FE_PHN2133_U_afifo_n3), 
	.A(U_afifo_n3));
   BUF_X32 FE_PHC2132_U_dfifo_U_dcore_U_sub_fifo_n400 (.Z(FE_PHN2132_U_dfifo_U_dcore_U_sub_fifo_n400), 
	.A(FE_PHN3701_U_dfifo_U_dcore_U_sub_fifo_n400));
   BUF_X32 FE_PHC2131_U_dfifo_U_dcore_U_sub_fifo_n328 (.Z(FE_PHN2131_U_dfifo_U_dcore_U_sub_fifo_n328), 
	.A(FE_PHN3670_U_dfifo_U_dcore_U_sub_fifo_n328));
   BUF_X32 FE_PHC2130_U_dfifo_U_dcore_U_sub_fifo_n438 (.Z(FE_PHN2130_U_dfifo_U_dcore_U_sub_fifo_n438), 
	.A(FE_PHN3675_U_dfifo_U_dcore_U_sub_fifo_n438));
   BUF_X32 FE_PHC2129_U_dfifo_U_dcore_U_sub_fifo_n342 (.Z(FE_PHN2129_U_dfifo_U_dcore_U_sub_fifo_n342), 
	.A(FE_PHN3650_U_dfifo_U_dcore_U_sub_fifo_n342));
   BUF_X32 FE_PHC2128_U_dfifo_U_dcore_U_sub_fifo_n320 (.Z(FE_PHN2128_U_dfifo_U_dcore_U_sub_fifo_n320), 
	.A(FE_PHN4746_U_dfifo_U_dcore_U_sub_fifo_n320));
   BUF_X32 FE_PHC2127_U_dfifo_U_dcore_U_sub_fifo_n414 (.Z(FE_PHN2127_U_dfifo_U_dcore_U_sub_fifo_n414), 
	.A(FE_PHN3703_U_dfifo_U_dcore_U_sub_fifo_n414));
   BUF_X32 FE_PHC2126_U_dfifo_U_dcore_U_sub_fifo_n319 (.Z(FE_PHN2126_U_dfifo_U_dcore_U_sub_fifo_n319), 
	.A(FE_PHN3678_U_dfifo_U_dcore_U_sub_fifo_n319));
   BUF_X32 FE_PHC2124_U_dfifo_U_dcore_U_sub_fifo_n312 (.Z(FE_PHN2124_U_dfifo_U_dcore_U_sub_fifo_n312), 
	.A(FE_PHN3652_U_dfifo_U_dcore_U_sub_fifo_n312));
   BUF_X32 FE_PHC2123_U_dfifo_U_dcore_U_sub_fifo_n323 (.Z(FE_PHN2123_U_dfifo_U_dcore_U_sub_fifo_n323), 
	.A(FE_PHN3696_U_dfifo_U_dcore_U_sub_fifo_n323));
   BUF_X32 FE_PHC2122_U_dfifo_U_dcore_U_sub_fifo_n406 (.Z(FE_PHN2122_U_dfifo_U_dcore_U_sub_fifo_n406), 
	.A(FE_PHN3710_U_dfifo_U_dcore_U_sub_fifo_n406));
   BUF_X32 FE_PHC2121_U_dfifo_U_dcore_U_sub_fifo_n412 (.Z(FE_PHN2121_U_dfifo_U_dcore_U_sub_fifo_n412), 
	.A(FE_PHN4747_U_dfifo_U_dcore_U_sub_fifo_n412));
   BUF_X32 FE_PHC2119_U_dfifo_U_dcore_U_sub_fifo_n444 (.Z(FE_PHN2119_U_dfifo_U_dcore_U_sub_fifo_n444), 
	.A(FE_PHN3676_U_dfifo_U_dcore_U_sub_fifo_n444));
   BUF_X32 FE_PHC2118_U_dfifo_U_dcore_U_sub_fifo_n441 (.Z(FE_PHN2118_U_dfifo_U_dcore_U_sub_fifo_n441), 
	.A(FE_PHN3689_U_dfifo_U_dcore_U_sub_fifo_n441));
   BUF_X32 FE_PHC2117_U_dfifo_U_dcore_U_sub_fifo_n409 (.Z(FE_PHN2117_U_dfifo_U_dcore_U_sub_fifo_n409), 
	.A(FE_PHN3658_U_dfifo_U_dcore_U_sub_fifo_n409));
   BUF_X32 FE_PHC2116_U_dfifo_U_dcore_U_sub_fifo_n408 (.Z(FE_PHN2116_U_dfifo_U_dcore_U_sub_fifo_n408), 
	.A(FE_PHN3667_U_dfifo_U_dcore_U_sub_fifo_n408));
   BUF_X32 FE_PHC2115_U_dfifo_U_dcore_U_sub_fifo_n369 (.Z(FE_PHN2115_U_dfifo_U_dcore_U_sub_fifo_n369), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n369));
   BUF_X32 FE_PHC2113_U_dfifo_U_dcore_U_sub_fifo_n311 (.Z(FE_PHN2113_U_dfifo_U_dcore_U_sub_fifo_n311), 
	.A(FE_PHN3695_U_dfifo_U_dcore_U_sub_fifo_n311));
   BUF_X32 FE_PHC2112_U_dfifo_U_dcore_U_sub_fifo_n404 (.Z(FE_PHN2112_U_dfifo_U_dcore_U_sub_fifo_n404), 
	.A(FE_PHN3694_U_dfifo_U_dcore_U_sub_fifo_n404));
   BUF_X32 FE_PHC2111_U_dfifo_U_dcore_U_sub_fifo_n439 (.Z(FE_PHN2111_U_dfifo_U_dcore_U_sub_fifo_n439), 
	.A(FE_PHN3688_U_dfifo_U_dcore_U_sub_fifo_n439));
   BUF_X32 FE_PHC2110_U_dfifo_U_dcore_U_sub_fifo_n372 (.Z(FE_PHN2110_U_dfifo_U_dcore_U_sub_fifo_n372), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n372));
   BUF_X32 FE_PHC2108_U_dfifo_U_dcore_U_sub_fifo_n316 (.Z(FE_PHN2108_U_dfifo_U_dcore_U_sub_fifo_n316), 
	.A(FE_PHN4742_U_dfifo_U_dcore_U_sub_fifo_n316));
   BUF_X32 FE_PHC2026_U_afifo_U_acore_U_sub_fifo_n298 (.Z(FE_PHN2026_U_afifo_U_acore_U_sub_fifo_n298), 
	.A(U_afifo_U_acore_U_sub_fifo_n298));
   BUF_X32 FE_PHC2024_U_afifo_U_acore_U_sub_fifo_n223 (.Z(FE_PHN2024_U_afifo_U_acore_U_sub_fifo_n223), 
	.A(FE_PHN3504_U_afifo_U_acore_U_sub_fifo_n223));
   BUF_X32 FE_PHC2023_U_dfifo_U_dcore_U_sub_fifo_n264 (.Z(FE_PHN2023_U_dfifo_U_dcore_U_sub_fifo_n264), 
	.A(FE_PHN4281_U_dfifo_U_dcore_U_sub_fifo_n264));
   BUF_X32 FE_PHC2022_U_afifo_U_acore_U_sub_fifo_n275 (.Z(FE_PHN2022_U_afifo_U_acore_U_sub_fifo_n275), 
	.A(FE_PHN5117_U_afifo_U_acore_U_sub_fifo_n275));
   BUF_X32 FE_PHC2021_U_afifo_U_acore_U_sub_fifo_n250 (.Z(FE_PHN2021_U_afifo_U_acore_U_sub_fifo_n250), 
	.A(FE_PHN5118_U_afifo_U_acore_U_sub_fifo_n250));
   BUF_X32 FE_PHC2020_U_afifo_U_acore_U_sub_fifo_n218 (.Z(FE_PHN2020_U_afifo_U_acore_U_sub_fifo_n218), 
	.A(FE_PHN4973_U_afifo_U_acore_U_sub_fifo_n218));
   BUF_X32 FE_PHC2019_U_afifo_U_acore_U_sub_fifo_n176 (.Z(FE_PHN2019_U_afifo_U_acore_U_sub_fifo_n176), 
	.A(FE_PHN3306_U_afifo_U_acore_U_sub_fifo_n176));
   BUF_X32 FE_PHC2018_U_afifo_U_acore_U_sub_fifo_n196 (.Z(FE_PHN2018_U_afifo_U_acore_U_sub_fifo_n196), 
	.A(FE_PHN4203_U_afifo_U_acore_U_sub_fifo_n196));
   BUF_X32 FE_PHC2017_U_afifo_U_acore_U_sub_fifo_n175 (.Z(FE_PHN2017_U_afifo_U_acore_U_sub_fifo_n175), 
	.A(FE_PHN4065_U_afifo_U_acore_U_sub_fifo_n175));
   BUF_X32 FE_PHC2016_U_afifo_U_acore_U_sub_fifo_n311 (.Z(FE_PHN2016_U_afifo_U_acore_U_sub_fifo_n311), 
	.A(U_afifo_U_acore_U_sub_fifo_n311));
   BUF_X32 FE_PHC2015_U_afifo_U_acore_U_sub_fifo_n174 (.Z(FE_PHN2015_U_afifo_U_acore_U_sub_fifo_n174), 
	.A(FE_PHN3998_U_afifo_U_acore_U_sub_fifo_n174));
   BUF_X32 FE_PHC2014_U_afifo_U_acore_U_sub_fifo_n309 (.Z(FE_PHN2014_U_afifo_U_acore_U_sub_fifo_n309), 
	.A(FE_PHN5081_U_afifo_U_acore_U_sub_fifo_n309));
   BUF_X32 FE_PHC2013_U_afifo_U_acore_U_sub_fifo_n230 (.Z(FE_PHN2013_U_afifo_U_acore_U_sub_fifo_n230), 
	.A(FE_PHN4080_U_afifo_U_acore_U_sub_fifo_n230));
   BUF_X32 FE_PHC2012_U_afifo_U_acore_U_sub_fifo_n207 (.Z(FE_PHN2012_U_afifo_U_acore_U_sub_fifo_n207), 
	.A(FE_PHN4014_U_afifo_U_acore_U_sub_fifo_n207));
   BUF_X32 FE_PHC2011_U_afifo_U_acore_U_sub_fifo_n261 (.Z(FE_PHN2011_U_afifo_U_acore_U_sub_fifo_n261), 
	.A(FE_PHN3999_U_afifo_U_acore_U_sub_fifo_n261));
   BUF_X32 FE_PHC2010_U_afifo_U_acore_U_sub_fifo_n247 (.Z(FE_PHN2010_U_afifo_U_acore_U_sub_fifo_n247), 
	.A(FE_PHN4978_U_afifo_U_acore_U_sub_fifo_n247));
   BUF_X32 FE_PHC2009_U_afifo_U_acore_U_sub_fifo_n193 (.Z(FE_PHN2009_U_afifo_U_acore_U_sub_fifo_n193), 
	.A(FE_PHN3486_U_afifo_U_acore_U_sub_fifo_n193));
   BUF_X32 FE_PHC2008_U_afifo_U_acore_U_sub_fifo_n178 (.Z(FE_PHN2008_U_afifo_U_acore_U_sub_fifo_n178), 
	.A(FE_PHN4066_U_afifo_U_acore_U_sub_fifo_n178));
   BUF_X32 FE_PHC2007_U_afifo_U_acore_U_sub_fifo_n202 (.Z(FE_PHN2007_U_afifo_U_acore_U_sub_fifo_n202), 
	.A(FE_PHN4996_U_afifo_U_acore_U_sub_fifo_n202));
   BUF_X32 FE_PHC2006_U_afifo_U_acore_U_sub_fifo_n201 (.Z(FE_PHN2006_U_afifo_U_acore_U_sub_fifo_n201), 
	.A(FE_PHN3301_U_afifo_U_acore_U_sub_fifo_n201));
   BUF_X32 FE_PHC2005_U_afifo_U_acore_U_sub_fifo_n244 (.Z(FE_PHN2005_U_afifo_U_acore_U_sub_fifo_n244), 
	.A(FE_PHN3978_U_afifo_U_acore_U_sub_fifo_n244));
   BUF_X32 FE_PHC2004_U_dfifo_U_dcore_U_sub_fifo_n378 (.Z(FE_PHN2004_U_dfifo_U_dcore_U_sub_fifo_n378), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n378));
   BUF_X32 FE_PHC2003_U_afifo_U_acore_U_sub_fifo_n293 (.Z(FE_PHN2003_U_afifo_U_acore_U_sub_fifo_n293), 
	.A(U_afifo_U_acore_U_sub_fifo_n293));
   BUF_X32 FE_PHC2002_U_afifo_U_acore_U_sub_fifo_n313 (.Z(FE_PHN2002_U_afifo_U_acore_U_sub_fifo_n313), 
	.A(U_afifo_U_acore_U_sub_fifo_n313));
   BUF_X32 FE_PHC2001_U_afifo_U_acore_U_sub_fifo_n195 (.Z(FE_PHN2001_U_afifo_U_acore_U_sub_fifo_n195), 
	.A(FE_PHN4011_U_afifo_U_acore_U_sub_fifo_n195));
   BUF_X32 FE_PHC2000_U_afifo_U_acore_U_sub_fifo_n263 (.Z(FE_PHN2000_U_afifo_U_acore_U_sub_fifo_n263), 
	.A(FE_PHN4100_U_afifo_U_acore_U_sub_fifo_n263));
   BUF_X32 FE_PHC1999_U_afifo_U_acore_U_sub_fifo_n229 (.Z(FE_PHN1999_U_afifo_U_acore_U_sub_fifo_n229), 
	.A(FE_PHN4951_U_afifo_U_acore_U_sub_fifo_n229));
   BUF_X32 FE_PHC1998_U_afifo_U_acore_U_sub_fifo_n299 (.Z(FE_PHN1998_U_afifo_U_acore_U_sub_fifo_n299), 
	.A(U_afifo_U_acore_U_sub_fifo_n299));
   BUF_X32 FE_PHC1997_U_dfifo_U_dcore_U_sub_fifo_n375 (.Z(FE_PHN1997_U_dfifo_U_dcore_U_sub_fifo_n375), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n375));
   BUF_X32 FE_PHC1996_U_afifo_U_acore_U_sub_fifo_n217 (.Z(FE_PHN1996_U_afifo_U_acore_U_sub_fifo_n217), 
	.A(FE_PHN3914_U_afifo_U_acore_U_sub_fifo_n217));
   BUF_X32 FE_PHC1995_U_afifo_U_acore_U_sub_fifo_n251 (.Z(FE_PHN1995_U_afifo_U_acore_U_sub_fifo_n251), 
	.A(FE_PHN5098_U_afifo_U_acore_U_sub_fifo_n251));
   BUF_X32 FE_PHC1994_U_afifo_U_acore_U_sub_fifo_n206 (.Z(FE_PHN1994_U_afifo_U_acore_U_sub_fifo_n206), 
	.A(FE_PHN3302_U_afifo_U_acore_U_sub_fifo_n206));
   BUF_X32 FE_PHC1993_U_afifo_U_acore_U_sub_fifo_n225 (.Z(FE_PHN1993_U_afifo_U_acore_U_sub_fifo_n225), 
	.A(FE_PHN3945_U_afifo_U_acore_U_sub_fifo_n225));
   BUF_X32 FE_PHC1992_U_afifo_U_acore_U_sub_fifo_n303 (.Z(FE_PHN1992_U_afifo_U_acore_U_sub_fifo_n303), 
	.A(U_afifo_U_acore_U_sub_fifo_n303));
   BUF_X32 FE_PHC1991_U_afifo_U_acore_U_sub_fifo_n260 (.Z(FE_PHN1991_U_afifo_U_acore_U_sub_fifo_n260), 
	.A(FE_PHN5164_U_afifo_U_acore_U_sub_fifo_n260));
   BUF_X32 FE_PHC1990_U_dfifo_U_dcore_U_sub_fifo_n377 (.Z(FE_PHN1990_U_dfifo_U_dcore_U_sub_fifo_n377), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n377));
   BUF_X32 FE_PHC1989_U_afifo_U_acore_U_sub_fifo_n233 (.Z(FE_PHN1989_U_afifo_U_acore_U_sub_fifo_n233), 
	.A(FE_PHN3956_U_afifo_U_acore_U_sub_fifo_n233));
   BUF_X32 FE_PHC1988_U_afifo_U_acore_U_sub_fifo_n187 (.Z(FE_PHN1988_U_afifo_U_acore_U_sub_fifo_n187), 
	.A(FE_PHN5005_U_afifo_U_acore_U_sub_fifo_n187));
   BUF_X32 FE_PHC1987_U_afifo_U_acore_U_sub_fifo_n184 (.Z(FE_PHN1987_U_afifo_U_acore_U_sub_fifo_n184), 
	.A(FE_PHN5020_U_afifo_U_acore_U_sub_fifo_n184));
   BUF_X32 FE_PHC1986_U_afifo_U_acore_U_sub_fifo_n255 (.Z(FE_PHN1986_U_afifo_U_acore_U_sub_fifo_n255), 
	.A(FE_PHN5048_U_afifo_U_acore_U_sub_fifo_n255));
   BUF_X32 FE_PHC1985_U_afifo_U_acore_U_sub_fifo_n285 (.Z(FE_PHN1985_U_afifo_U_acore_U_sub_fifo_n285), 
	.A(FE_PHN5007_U_afifo_U_acore_U_sub_fifo_n285));
   BUF_X32 FE_PHC1984_U_afifo_U_acore_U_sub_fifo_n291 (.Z(FE_PHN1984_U_afifo_U_acore_U_sub_fifo_n291), 
	.A(FE_PHN4127_U_afifo_U_acore_U_sub_fifo_n291));
   BUF_X32 FE_PHC1982_U_afifo_U_acore_U_sub_fifo_n242 (.Z(FE_PHN1982_U_afifo_U_acore_U_sub_fifo_n242), 
	.A(FE_PHN4009_U_afifo_U_acore_U_sub_fifo_n242));
   BUF_X32 FE_PHC1981_U_afifo_U_acore_U_sub_fifo_n281 (.Z(FE_PHN1981_U_afifo_U_acore_U_sub_fifo_n281), 
	.A(FE_PHN3955_U_afifo_U_acore_U_sub_fifo_n281));
   BUF_X32 FE_PHC1980_U_afifo_U_acore_U_sub_fifo_n236 (.Z(FE_PHN1980_U_afifo_U_acore_U_sub_fifo_n236), 
	.A(FE_PHN5133_U_afifo_U_acore_U_sub_fifo_n236));
   BUF_X32 FE_PHC1979_U_afifo_U_acore_U_sub_fifo_n239 (.Z(FE_PHN1979_U_afifo_U_acore_U_sub_fifo_n239), 
	.A(FE_PHN3940_U_afifo_U_acore_U_sub_fifo_n239));
   BUF_X32 FE_PHC1977_U_afifo_U_acore_U_sub_fifo_n304 (.Z(FE_PHN1977_U_afifo_U_acore_U_sub_fifo_n304), 
	.A(FE_PHN4019_U_afifo_U_acore_U_sub_fifo_n304));
   BUF_X32 FE_PHC1976_U_afifo_U_acore_U_sub_fifo_n240 (.Z(FE_PHN1976_U_afifo_U_acore_U_sub_fifo_n240), 
	.A(FE_PHN4964_U_afifo_U_acore_U_sub_fifo_n240));
   BUF_X32 FE_PHC1975_U_afifo_U_acore_U_sub_fifo_n188 (.Z(FE_PHN1975_U_afifo_U_acore_U_sub_fifo_n188), 
	.A(FE_PHN5143_U_afifo_U_acore_U_sub_fifo_n188));
   BUF_X32 FE_PHC1974_U_afifo_U_acore_U_sub_fifo_n220 (.Z(FE_PHN1974_U_afifo_U_acore_U_sub_fifo_n220), 
	.A(FE_PHN5111_U_afifo_U_acore_U_sub_fifo_n220));
   BUF_X32 FE_PHC1973_U_afifo_U_acore_U_sub_fifo_n238 (.Z(FE_PHN1973_U_afifo_U_acore_U_sub_fifo_n238), 
	.A(FE_PHN3995_U_afifo_U_acore_U_sub_fifo_n238));
   BUF_X32 FE_PHC1972_U_afifo_U_acore_U_sub_fifo_n320 (.Z(FE_PHN1972_U_afifo_U_acore_U_sub_fifo_n320), 
	.A(FE_PHN4877_U_afifo_U_acore_U_sub_fifo_n320));
   BUF_X32 FE_PHC1971_U_afifo_U_acore_U_sub_fifo_n282 (.Z(FE_PHN1971_U_afifo_U_acore_U_sub_fifo_n282), 
	.A(FE_PHN5165_U_afifo_U_acore_U_sub_fifo_n282));
   BUF_X32 FE_PHC1969_U_dfifo_U_dcore_U_sub_fifo_n349 (.Z(FE_PHN1969_U_dfifo_U_dcore_U_sub_fifo_n349), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n349));
   BUF_X32 FE_PHC1968_U_dfifo_U_dcore_U_sub_fifo_n364 (.Z(FE_PHN1968_U_dfifo_U_dcore_U_sub_fifo_n364), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n364));
   BUF_X32 FE_PHC1966_U_afifo_U_acore_U_sub_fifo_n267 (.Z(FE_PHN1966_U_afifo_U_acore_U_sub_fifo_n267), 
	.A(FE_PHN4819_U_afifo_U_acore_U_sub_fifo_n267));
   BUF_X32 FE_PHC1965_U_dfifo_U_dcore_U_sub_fifo_n352 (.Z(FE_PHN1965_U_dfifo_U_dcore_U_sub_fifo_n352), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n352));
   BUF_X32 FE_PHC1964_U_dfifo_U_dcore_U_sub_fifo_n330 (.Z(FE_PHN1964_U_dfifo_U_dcore_U_sub_fifo_n330), 
	.A(FE_PHN3804_U_dfifo_U_dcore_U_sub_fifo_n330));
   BUF_X32 FE_PHC1963_U_dfifo_U_dcore_U_sub_fifo_n360 (.Z(FE_PHN1963_U_dfifo_U_dcore_U_sub_fifo_n360), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n360));
   BUF_X32 FE_PHC1962_U_afifo_U_acore_U_sub_fifo_n272 (.Z(FE_PHN1962_U_afifo_U_acore_U_sub_fifo_n272), 
	.A(FE_PHN3813_U_afifo_U_acore_U_sub_fifo_n272));
   BUF_X32 FE_PHC1961_U_dfifo_U_dcore_U_sub_fifo_n346 (.Z(FE_PHN1961_U_dfifo_U_dcore_U_sub_fifo_n346), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n346));
   BUF_X32 FE_PHC1960_U_dfifo_U_dcore_U_sub_fifo_n351 (.Z(FE_PHN1960_U_dfifo_U_dcore_U_sub_fifo_n351), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n351));
   BUF_X32 FE_PHC1959_U_afifo_U_acore_U_sub_fifo_n266 (.Z(FE_PHN1959_U_afifo_U_acore_U_sub_fifo_n266), 
	.A(FE_PHN4793_U_afifo_U_acore_U_sub_fifo_n266));
   BUF_X32 FE_PHC1958_U_dfifo_U_dcore_U_sub_fifo_n367 (.Z(FE_PHN1958_U_dfifo_U_dcore_U_sub_fifo_n367), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n367));
   BUF_X32 FE_PHC1957_U_dfifo_U_dcore_U_sub_fifo_n347 (.Z(FE_PHN1957_U_dfifo_U_dcore_U_sub_fifo_n347), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n347));
   BUF_X32 FE_PHC1956_U_dfifo_U_dcore_U_sub_fifo_n407 (.Z(FE_PHN1956_U_dfifo_U_dcore_U_sub_fifo_n407), 
	.A(FE_PHN3750_U_dfifo_U_dcore_U_sub_fifo_n407));
   BUF_X32 FE_PHC1955_U_dfifo_U_dcore_U_sub_fifo_n358 (.Z(FE_PHN1955_U_dfifo_U_dcore_U_sub_fifo_n358), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n358));
   BUF_X32 FE_PHC1954_U_dfifo_U_dcore_U_sub_fifo_n398 (.Z(FE_PHN1954_U_dfifo_U_dcore_U_sub_fifo_n398), 
	.A(FE_PHN4765_U_dfifo_U_dcore_U_sub_fifo_n398));
   BUF_X32 FE_PHC1953_U_dfifo_U_dcore_U_sub_fifo_n415 (.Z(FE_PHN1953_U_dfifo_U_dcore_U_sub_fifo_n415), 
	.A(FE_PHN3801_U_dfifo_U_dcore_U_sub_fifo_n415));
   BUF_X32 FE_PHC1952_U_dfifo_U_dcore_U_sub_fifo_n348 (.Z(FE_PHN1952_U_dfifo_U_dcore_U_sub_fifo_n348), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n348));
   BUF_X32 FE_PHC1951_U_dfifo_U_dcore_U_sub_fifo_n318 (.Z(FE_PHN1951_U_dfifo_U_dcore_U_sub_fifo_n318), 
	.A(FE_PHN3728_U_dfifo_U_dcore_U_sub_fifo_n318));
   BUF_X32 FE_PHC1950_U_afifo_U_acore_U_sub_fifo_n269 (.Z(FE_PHN1950_U_afifo_U_acore_U_sub_fifo_n269), 
	.A(FE_PHN4758_U_afifo_U_acore_U_sub_fifo_n269));
   BUF_X32 FE_PHC1949_U_dfifo_U_dcore_U_sub_fifo_n345 (.Z(FE_PHN1949_U_dfifo_U_dcore_U_sub_fifo_n345), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n345));
   BUF_X32 FE_PHC1948_U_afifo_U_acore_U_sub_fifo_n270 (.Z(FE_PHN1948_U_afifo_U_acore_U_sub_fifo_n270), 
	.A(FE_PHN3772_U_afifo_U_acore_U_sub_fifo_n270));
   BUF_X32 FE_PHC1947_U_dfifo_U_dcore_U_sub_fifo_n397 (.Z(FE_PHN1947_U_dfifo_U_dcore_U_sub_fifo_n397), 
	.A(FE_PHN4766_U_dfifo_U_dcore_U_sub_fifo_n397));
   BUF_X32 FE_PHC1946_U_dfifo_U_dcore_U_sub_fifo_n362 (.Z(FE_PHN1946_U_dfifo_U_dcore_U_sub_fifo_n362), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n362));
   BUF_X32 FE_PHC1945_U_dfifo_U_dcore_U_sub_fifo_n355 (.Z(FE_PHN1945_U_dfifo_U_dcore_U_sub_fifo_n355), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n355));
   BUF_X32 FE_PHC1944_U_dfifo_U_dcore_U_sub_fifo_n399 (.Z(FE_PHN1944_U_dfifo_U_dcore_U_sub_fifo_n399), 
	.A(FE_PHN3706_U_dfifo_U_dcore_U_sub_fifo_n399));
   BUF_X32 FE_PHC1943_U_dfifo_U_dcore_U_sub_fifo_n357 (.Z(FE_PHN1943_U_dfifo_U_dcore_U_sub_fifo_n357), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n357));
   BUF_X32 FE_PHC1942_U_dfifo_U_dcore_U_sub_fifo_n371 (.Z(FE_PHN1942_U_dfifo_U_dcore_U_sub_fifo_n371), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n371));
   BUF_X32 FE_PHC1941_U_dfifo_U_dcore_U_sub_fifo_n353 (.Z(FE_PHN1941_U_dfifo_U_dcore_U_sub_fifo_n353), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n353));
   BUF_X32 FE_PHC1940_U_dfifo_U_dcore_U_sub_fifo_n341 (.Z(FE_PHN1940_U_dfifo_U_dcore_U_sub_fifo_n341), 
	.A(FE_PHN3668_U_dfifo_U_dcore_U_sub_fifo_n341));
   BUF_X32 FE_PHC1939_U_dfifo_U_dcore_U_sub_fifo_n327 (.Z(FE_PHN1939_U_dfifo_U_dcore_U_sub_fifo_n327), 
	.A(FE_PHN4751_U_dfifo_U_dcore_U_sub_fifo_n327));
   BUF_X32 FE_PHC1938_U_dfifo_U_dcore_U_sub_fifo_n417 (.Z(FE_PHN1938_U_dfifo_U_dcore_U_sub_fifo_n417), 
	.A(FE_PHN3743_U_dfifo_U_dcore_U_sub_fifo_n417));
   BUF_X32 FE_PHC1937_U_dfifo_U_dcore_U_sub_fifo_n340 (.Z(FE_PHN1937_U_dfifo_U_dcore_U_sub_fifo_n340), 
	.A(FE_PHN4740_U_dfifo_U_dcore_U_sub_fifo_n340));
   BUF_X32 FE_PHC1936_U_dfifo_U_dcore_U_sub_fifo_n324 (.Z(FE_PHN1936_U_dfifo_U_dcore_U_sub_fifo_n324), 
	.A(FE_PHN3742_U_dfifo_U_dcore_U_sub_fifo_n324));
   BUF_X32 FE_PHC1935_U_dfifo_U_dcore_U_sub_fifo_n440 (.Z(FE_PHN1935_U_dfifo_U_dcore_U_sub_fifo_n440), 
	.A(FE_PHN4752_U_dfifo_U_dcore_U_sub_fifo_n440));
   BUF_X32 FE_PHC1933_U_dfifo_U_dcore_U_sub_fifo_n343 (.Z(FE_PHN1933_U_dfifo_U_dcore_U_sub_fifo_n343), 
	.A(FE_PHN3679_U_dfifo_U_dcore_U_sub_fifo_n343));
   BUF_X32 FE_PHC1932_U_dfifo_U_dcore_U_sub_fifo_n334 (.Z(FE_PHN1932_U_dfifo_U_dcore_U_sub_fifo_n334), 
	.A(FE_PHN3691_U_dfifo_U_dcore_U_sub_fifo_n334));
   BUF_X32 FE_PHC1931_U_dfifo_U_dcore_U_sub_fifo_n442 (.Z(FE_PHN1931_U_dfifo_U_dcore_U_sub_fifo_n442), 
	.A(FE_PHN4755_U_dfifo_U_dcore_U_sub_fifo_n442));
   BUF_X32 FE_PHC1930_U_dfifo_U_dcore_U_sub_fifo_n418 (.Z(FE_PHN1930_U_dfifo_U_dcore_U_sub_fifo_n418), 
	.A(FE_PHN3685_U_dfifo_U_dcore_U_sub_fifo_n418));
   BUF_X32 FE_PHC1929_U_dfifo_U_dcore_U_sub_fifo_n446 (.Z(FE_PHN1929_U_dfifo_U_dcore_U_sub_fifo_n446), 
	.A(FE_PHN4738_U_dfifo_U_dcore_U_sub_fifo_n446));
   BUF_X32 FE_PHC1928_U_dfifo_U_dcore_U_sub_fifo_n359 (.Z(FE_PHN1928_U_dfifo_U_dcore_U_sub_fifo_n359), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n359));
   BUF_X32 FE_PHC1927_U_dfifo_U_dcore_U_sub_fifo_n356 (.Z(FE_PHN1927_U_dfifo_U_dcore_U_sub_fifo_n356), 
	.A(FE_PHN4754_U_dfifo_U_dcore_U_sub_fifo_n356));
   BUF_X32 FE_PHC1926_U_dfifo_U_dcore_U_sub_fifo_n410 (.Z(FE_PHN1926_U_dfifo_U_dcore_U_sub_fifo_n410), 
	.A(FE_PHN3664_U_dfifo_U_dcore_U_sub_fifo_n410));
   BUF_X32 FE_PHC1925_U_dfifo_U_dcore_U_sub_fifo_n331 (.Z(FE_PHN1925_U_dfifo_U_dcore_U_sub_fifo_n331), 
	.A(FE_PHN3693_U_dfifo_U_dcore_U_sub_fifo_n331));
   BUF_X32 FE_PHC1924_U_dfifo_U_dcore_U_sub_fifo_n370 (.Z(FE_PHN1924_U_dfifo_U_dcore_U_sub_fifo_n370), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n370));
   BUF_X32 FE_PHC1923_U_dfifo_U_dcore_U_sub_fifo_n335 (.Z(FE_PHN1923_U_dfifo_U_dcore_U_sub_fifo_n335), 
	.A(FE_PHN3656_U_dfifo_U_dcore_U_sub_fifo_n335));
   BUF_X32 FE_PHC1922_U_dfifo_U_dcore_U_sub_fifo_n354 (.Z(FE_PHN1922_U_dfifo_U_dcore_U_sub_fifo_n354), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n354));
   BUF_X32 FE_PHC1907_U_afifo_m_data_in_7_ (.Z(FE_PHN1907_U_afifo_m_data_in_7_), 
	.A(U_afifo_m_data_in[7]));
   BUF_X32 FE_PHC1904_U_ctl_n141 (.Z(FE_PHN1904_U_ctl_n141), 
	.A(FE_PHN3271_U_ctl_n141));
   BUF_X32 FE_PHC1886_U_afifo_f_data2_38_ (.Z(FE_PHN1886_U_afifo_f_data2_38_), 
	.A(U_afifo_f_data2_38_));
   BUF_X32 FE_PHC1885_U_afifo_f_data2_44_ (.Z(FE_PHN1885_U_afifo_f_data2_44_), 
	.A(U_afifo_f_data2_44_));
   BUF_X32 FE_PHC1884_U_afifo_f_data2_42_ (.Z(FE_PHN1884_U_afifo_f_data2_42_), 
	.A(U_afifo_f_data2_42_));
   BUF_X32 FE_PHC1883_U_afifo_f_data2_31_ (.Z(FE_PHN1883_U_afifo_f_data2_31_), 
	.A(U_afifo_f_data2_31_));
   BUF_X32 FE_PHC1882_U_afifo_f_data2_18_ (.Z(FE_PHN1882_U_afifo_f_data2_18_), 
	.A(U_afifo_f_data2_18_));
   BUF_X32 FE_PHC1881_U_afifo_f_data2_5_ (.Z(FE_PHN1881_U_afifo_f_data2_5_), 
	.A(U_afifo_f_data2_5_));
   BUF_X32 FE_PHC1880_U_afifo_f_data2_20_ (.Z(FE_PHN1880_U_afifo_f_data2_20_), 
	.A(U_afifo_f_data2_20_));
   BUF_X32 FE_PHC1879_U_afifo_f_data2_0_ (.Z(FE_PHN1879_U_afifo_f_data2_0_), 
	.A(U_afifo_f_data2_0_));
   BUF_X32 FE_PHC1878_U_afifo_f_data2_37_ (.Z(FE_PHN1878_U_afifo_f_data2_37_), 
	.A(U_afifo_f_data2_37_));
   BUF_X32 FE_PHC1877_U_afifo_f_data2_6_ (.Z(FE_PHN1877_U_afifo_f_data2_6_), 
	.A(U_afifo_f_data2_6_));
   BUF_X32 FE_PHC1876_U_afifo_f_data2_24_ (.Z(FE_PHN1876_U_afifo_f_data2_24_), 
	.A(U_afifo_f_data2_24_));
   BUF_X32 FE_PHC1874_U_afifo_f_data2_23_ (.Z(FE_PHN1874_U_afifo_f_data2_23_), 
	.A(U_afifo_f_data2_23_));
   BUF_X32 FE_PHC1873_U_afifo_f_data2_26_ (.Z(FE_PHN1873_U_afifo_f_data2_26_), 
	.A(U_afifo_f_data2_26_));
   BUF_X32 FE_PHC1872_U_afifo_f_data2_43_ (.Z(FE_PHN1872_U_afifo_f_data2_43_), 
	.A(U_afifo_f_data2_43_));
   BUF_X32 FE_PHC1871_U_afifo_f_data2_39_ (.Z(FE_PHN1871_U_afifo_f_data2_39_), 
	.A(U_afifo_f_data2_39_));
   BUF_X32 FE_PHC1870_U_afifo_f_data2_35_ (.Z(FE_PHN1870_U_afifo_f_data2_35_), 
	.A(U_afifo_f_data2_35_));
   BUF_X32 FE_PHC1869_U_afifo_f_data2_40_ (.Z(FE_PHN1869_U_afifo_f_data2_40_), 
	.A(U_afifo_f_data2_40_));
   BUF_X32 FE_PHC1867_U_afifo_f_data2_27_ (.Z(FE_PHN1867_U_afifo_f_data2_27_), 
	.A(U_afifo_f_data2_27_));
   BUF_X32 FE_PHC1866_U_afifo_f_data2_29_ (.Z(FE_PHN1866_U_afifo_f_data2_29_), 
	.A(U_afifo_f_data2_29_));
   BUF_X32 FE_PHC1865_U_afifo_f_data2_25_ (.Z(FE_PHN1865_U_afifo_f_data2_25_), 
	.A(U_afifo_f_data2_25_));
   BUF_X32 FE_PHC1864_U_afifo_f_data2_22_ (.Z(FE_PHN1864_U_afifo_f_data2_22_), 
	.A(U_afifo_f_data2_22_));
   BUF_X32 FE_PHC1863_U_afifo_f_data2_32_ (.Z(FE_PHN1863_U_afifo_f_data2_32_), 
	.A(U_afifo_f_data2_32_));
   BUF_X32 FE_PHC1862_U_afifo_f_data2_2_ (.Z(FE_PHN1862_U_afifo_f_data2_2_), 
	.A(U_afifo_f_data2_2_));
   BUF_X32 FE_PHC1861_U_afifo_f_data2_30_ (.Z(FE_PHN1861_U_afifo_f_data2_30_), 
	.A(U_afifo_f_data2_30_));
   BUF_X32 FE_PHC1860_U_afifo_f_data2_19_ (.Z(FE_PHN1860_U_afifo_f_data2_19_), 
	.A(U_afifo_f_data2_19_));
   BUF_X32 FE_PHC1859_U_afifo_f_data2_36_ (.Z(FE_PHN1859_U_afifo_f_data2_36_), 
	.A(U_afifo_f_data2_36_));
   BUF_X32 FE_PHC1858_U_afifo_f_data2_28_ (.Z(FE_PHN1858_U_afifo_f_data2_28_), 
	.A(U_afifo_f_data2_28_));
   BUF_X32 FE_PHC1857_U_afifo_f_data2_34_ (.Z(FE_PHN1857_U_afifo_f_data2_34_), 
	.A(U_afifo_f_data2_34_));
   BUF_X32 FE_PHC1856_U_afifo_f_data2_33_ (.Z(FE_PHN1856_U_afifo_f_data2_33_), 
	.A(U_afifo_f_data2_33_));
   BUF_X32 FE_PHC1853_U_afifo_f_data2_21_ (.Z(FE_PHN1853_U_afifo_f_data2_21_), 
	.A(U_afifo_f_data2_21_));
   CLKBUF_X1 FE_PHC1852_U_afifo_U_acore_n100 (.Z(FE_PHN1852_U_afifo_U_acore_n100), 
	.A(U_afifo_U_acore_n100));
   BUF_X32 FE_PHC1851_U_afifo_U_acore_n96 (.Z(FE_PHN1851_U_afifo_U_acore_n96), 
	.A(U_afifo_U_acore_n96));
   CLKBUF_X1 FE_PHC1850_U_afifo_U_acore_n98 (.Z(FE_PHN1850_U_afifo_U_acore_n98), 
	.A(U_afifo_U_acore_n98));
   BUF_X32 FE_PHC1849_U_afifo_U_acore_n207 (.Z(FE_PHN1849_U_afifo_U_acore_n207), 
	.A(U_afifo_U_acore_n207));
   CLKBUF_X1 FE_PHC1847_U_afifo_U_acore_n181 (.Z(FE_PHN1847_U_afifo_U_acore_n181), 
	.A(U_afifo_U_acore_n181));
   CLKBUF_X1 FE_PHC1844_U_afifo_U_acore_n201 (.Z(FE_PHN1844_U_afifo_U_acore_n201), 
	.A(U_afifo_U_acore_n201));
   BUF_X32 FE_PHC1843_U_afifo_U_acore_U_sub_fifo_n126 (.Z(FE_PHN1843_U_afifo_U_acore_U_sub_fifo_n126), 
	.A(U_afifo_U_acore_U_sub_fifo_n126));
   BUF_X32 FE_PHC1842_U_dfifo_U_dcore_U_sub_fifo_n451 (.Z(FE_PHN1842_U_dfifo_U_dcore_U_sub_fifo_n451), 
	.A(FE_PHN4299_U_dfifo_U_dcore_U_sub_fifo_n451));
   BUF_X32 FE_PHC1841_U_afifo_U_acore_n184 (.Z(FE_PHN1841_U_afifo_U_acore_n184), 
	.A(U_afifo_U_acore_n184));
   CLKBUF_X1 FE_PHC1840_U_afifo_U_acore_n194 (.Z(FE_PHN1840_U_afifo_U_acore_n194), 
	.A(U_afifo_U_acore_n194));
   BUF_X32 FE_PHC1839_U_afifo_U_acore_n203 (.Z(FE_PHN1839_U_afifo_U_acore_n203), 
	.A(U_afifo_U_acore_n203));
   BUF_X32 FE_PHC1838_n37 (.Z(FE_PHN1838_n37), 
	.A(n37));
   BUF_X32 FE_PHC1837_U_afifo_U_acore_n102 (.Z(FE_PHN1837_U_afifo_U_acore_n102), 
	.A(U_afifo_U_acore_n102));
   BUF_X32 FE_PHC1836_U_afifo_U_acore_n210 (.Z(FE_PHN1836_U_afifo_U_acore_n210), 
	.A(U_afifo_U_acore_n210));
   BUF_X32 FE_PHC1835_U_afifo_U_acore_n197 (.Z(FE_PHN1835_U_afifo_U_acore_n197), 
	.A(U_afifo_U_acore_n197));
   BUF_X32 FE_PHC1834_U_afifo_U_acore_n177 (.Z(FE_PHN1834_U_afifo_U_acore_n177), 
	.A(U_afifo_U_acore_n177));
   BUF_X32 FE_PHC1833_U_afifo_U_acore_U_sub_fifo_n133 (.Z(FE_PHN1833_U_afifo_U_acore_U_sub_fifo_n133), 
	.A(U_afifo_U_acore_U_sub_fifo_n133));
   BUF_X32 FE_PHC1832_U_afifo_U_acore_U_sub_fifo_n129 (.Z(FE_PHN1832_U_afifo_U_acore_U_sub_fifo_n129), 
	.A(U_afifo_U_acore_U_sub_fifo_n129));
   BUF_X32 FE_PHC1831_U_afifo_U_acore_U_sub_fifo_n115 (.Z(FE_PHN1831_U_afifo_U_acore_U_sub_fifo_n115), 
	.A(U_afifo_U_acore_U_sub_fifo_n115));
   BUF_X32 FE_PHC1830_U_afifo_U_acore_U_sub_fifo_n148 (.Z(FE_PHN1830_U_afifo_U_acore_U_sub_fifo_n148), 
	.A(U_afifo_U_acore_U_sub_fifo_n148));
   BUF_X32 FE_PHC1829_U_afifo_U_acore_U_sub_fifo_n273 (.Z(FE_PHN1829_U_afifo_U_acore_U_sub_fifo_n273), 
	.A(FE_PHN5009_U_afifo_U_acore_U_sub_fifo_n273));
   BUF_X32 FE_PHC1828_U_afifo_U_acore_U_sub_fifo_n130 (.Z(FE_PHN1828_U_afifo_U_acore_U_sub_fifo_n130), 
	.A(U_afifo_U_acore_U_sub_fifo_n130));
   BUF_X32 FE_PHC1827_U_afifo_U_acore_U_sub_fifo_n125 (.Z(FE_PHN1827_U_afifo_U_acore_U_sub_fifo_n125), 
	.A(U_afifo_U_acore_U_sub_fifo_n125));
   BUF_X32 FE_PHC1826_U_afifo_U_acore_U_sub_fifo_n134 (.Z(FE_PHN1826_U_afifo_U_acore_U_sub_fifo_n134), 
	.A(U_afifo_U_acore_U_sub_fifo_n134));
   BUF_X32 FE_PHC1825_U_afifo_U_acore_U_sub_fifo_n106 (.Z(FE_PHN1825_U_afifo_U_acore_U_sub_fifo_n106), 
	.A(U_afifo_U_acore_U_sub_fifo_n106));
   BUF_X32 FE_PHC1824_U_afifo_U_acore_U_sub_fifo_n314 (.Z(FE_PHN1824_U_afifo_U_acore_U_sub_fifo_n314), 
	.A(FE_PHN4113_U_afifo_U_acore_U_sub_fifo_n314));
   BUF_X32 FE_PHC1823_U_afifo_U_acore_U_sub_fifo_n264 (.Z(FE_PHN1823_U_afifo_U_acore_U_sub_fifo_n264), 
	.A(FE_PHN5071_U_afifo_U_acore_U_sub_fifo_n264));
   BUF_X32 FE_PHC1822_U_afifo_U_acore_U_sub_fifo_n122 (.Z(FE_PHN1822_U_afifo_U_acore_U_sub_fifo_n122), 
	.A(U_afifo_U_acore_U_sub_fifo_n122));
   BUF_X32 FE_PHC1821_U_afifo_U_acore_U_sub_fifo_n136 (.Z(FE_PHN1821_U_afifo_U_acore_U_sub_fifo_n136), 
	.A(U_afifo_U_acore_U_sub_fifo_n136));
   BUF_X32 FE_PHC1820_U_afifo_U_acore_U_sub_fifo_n139 (.Z(FE_PHN1820_U_afifo_U_acore_U_sub_fifo_n139), 
	.A(U_afifo_U_acore_U_sub_fifo_n139));
   BUF_X32 FE_PHC1819_U_afifo_U_acore_U_sub_fifo_n219 (.Z(FE_PHN1819_U_afifo_U_acore_U_sub_fifo_n219), 
	.A(FE_PHN3494_U_afifo_U_acore_U_sub_fifo_n219));
   BUF_X32 FE_PHC1818_U_afifo_m_data_in_27_ (.Z(FE_PHN1818_U_afifo_m_data_in_27_), 
	.A(U_afifo_m_data_in[27]));
   BUF_X32 FE_PHC1817_U_afifo_f_data2_41_ (.Z(FE_PHN1817_U_afifo_f_data2_41_), 
	.A(U_afifo_f_data2_41_));
   BUF_X32 FE_PHC1816_U_afifo_U_acore_U_sub_fifo_n102 (.Z(FE_PHN1816_U_afifo_U_acore_U_sub_fifo_n102), 
	.A(U_afifo_U_acore_U_sub_fifo_n102));
   BUF_X32 FE_PHC1815_U_afifo_U_acore_U_sub_fifo_n143 (.Z(FE_PHN1815_U_afifo_U_acore_U_sub_fifo_n143), 
	.A(U_afifo_U_acore_U_sub_fifo_n143));
   BUF_X32 FE_PHC1814_U_afifo_U_acore_U_sub_fifo_n138 (.Z(FE_PHN1814_U_afifo_U_acore_U_sub_fifo_n138), 
	.A(U_afifo_U_acore_U_sub_fifo_n138));
   BUF_X32 FE_PHC1813_U_afifo_U_acore_U_sub_fifo_n216 (.Z(FE_PHN1813_U_afifo_U_acore_U_sub_fifo_n216), 
	.A(FE_PHN3984_U_afifo_U_acore_U_sub_fifo_n216));
   BUF_X32 FE_PHC1812_U_afifo_U_acore_U_sub_fifo_n123 (.Z(FE_PHN1812_U_afifo_U_acore_U_sub_fifo_n123), 
	.A(U_afifo_U_acore_U_sub_fifo_n123));
   BUF_X32 FE_PHC1811_U_afifo_U_acore_U_sub_fifo_n214 (.Z(FE_PHN1811_U_afifo_U_acore_U_sub_fifo_n214), 
	.A(FE_PHN4858_U_afifo_U_acore_U_sub_fifo_n214));
   BUF_X32 FE_PHC1810_U_afifo_U_acore_U_sub_fifo_n121 (.Z(FE_PHN1810_U_afifo_U_acore_U_sub_fifo_n121), 
	.A(U_afifo_U_acore_U_sub_fifo_n121));
   BUF_X32 FE_PHC1808_U_afifo_U_acore_U_sub_fifo_n140 (.Z(FE_PHN1808_U_afifo_U_acore_U_sub_fifo_n140), 
	.A(U_afifo_U_acore_U_sub_fifo_n140));
   BUF_X32 FE_PHC1807_U_afifo_U_acore_U_sub_fifo_n317 (.Z(FE_PHN1807_U_afifo_U_acore_U_sub_fifo_n317), 
	.A(FE_PHN4112_U_afifo_U_acore_U_sub_fifo_n317));
   BUF_X32 FE_PHC1806_U_afifo_U_acore_U_sub_fifo_n128 (.Z(FE_PHN1806_U_afifo_U_acore_U_sub_fifo_n128), 
	.A(U_afifo_U_acore_U_sub_fifo_n128));
   BUF_X32 FE_PHC1805_U_afifo_U_acore_U_sub_fifo_n127 (.Z(FE_PHN1805_U_afifo_U_acore_U_sub_fifo_n127), 
	.A(U_afifo_U_acore_U_sub_fifo_n127));
   BUF_X32 FE_PHC1804_U_afifo_U_acore_U_sub_fifo_n146 (.Z(FE_PHN1804_U_afifo_U_acore_U_sub_fifo_n146), 
	.A(U_afifo_U_acore_U_sub_fifo_n146));
   BUF_X32 FE_PHC1803_U_afifo_U_acore_U_sub_fifo_n277 (.Z(FE_PHN1803_U_afifo_U_acore_U_sub_fifo_n277), 
	.A(FE_PHN4981_U_afifo_U_acore_U_sub_fifo_n277));
   BUF_X32 FE_PHC1802_U_dfifo_U_dcore_U_sub_fifo_n80 (.Z(FE_PHN1802_U_dfifo_U_dcore_U_sub_fifo_n80), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n80));
   BUF_X32 FE_PHC1801_U_afifo_U_acore_U_sub_fifo_n108 (.Z(FE_PHN1801_U_afifo_U_acore_U_sub_fifo_n108), 
	.A(U_afifo_U_acore_U_sub_fifo_n108));
   BUF_X32 FE_PHC1800_U_afifo_U_acore_U_sub_fifo_n145 (.Z(FE_PHN1800_U_afifo_U_acore_U_sub_fifo_n145), 
	.A(U_afifo_U_acore_U_sub_fifo_n145));
   BUF_X32 FE_PHC1799_U_afifo_U_acore_U_sub_fifo_n135 (.Z(FE_PHN1799_U_afifo_U_acore_U_sub_fifo_n135), 
	.A(U_afifo_U_acore_U_sub_fifo_n135));
   BUF_X32 FE_PHC1798_n27 (.Z(FE_PHN1798_n27), 
	.A(n27));
   BUF_X32 FE_PHC1797_U_afifo_U_acore_U_sub_fifo_n131 (.Z(FE_PHN1797_U_afifo_U_acore_U_sub_fifo_n131), 
	.A(U_afifo_U_acore_U_sub_fifo_n131));
   BUF_X32 FE_PHC1796_U_afifo_U_acore_U_sub_fifo_n120 (.Z(FE_PHN1796_U_afifo_U_acore_U_sub_fifo_n120), 
	.A(U_afifo_U_acore_U_sub_fifo_n120));
   BUF_X32 FE_PHC1795_U_dfifo_U_dcore_U_sub_fifo_n82 (.Z(FE_PHN1795_U_dfifo_U_dcore_U_sub_fifo_n82), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n82));
   BUF_X32 FE_PHC1794_U_afifo_U_acore_U_sub_fifo_n222 (.Z(FE_PHN1794_U_afifo_U_acore_U_sub_fifo_n222), 
	.A(FE_PHN4936_U_afifo_U_acore_U_sub_fifo_n222));
   BUF_X32 FE_PHC1793_U_afifo_U_acore_U_sub_fifo_n104 (.Z(FE_PHN1793_U_afifo_U_acore_U_sub_fifo_n104), 
	.A(U_afifo_U_acore_U_sub_fifo_n104));
   BUF_X32 FE_PHC1792_U_afifo_U_acore_U_sub_fifo_n124 (.Z(FE_PHN1792_U_afifo_U_acore_U_sub_fifo_n124), 
	.A(U_afifo_U_acore_U_sub_fifo_n124));
   BUF_X32 FE_PHC1791_U_dfifo_U_dcore_U_sub_fifo_n55 (.Z(FE_PHN1791_U_dfifo_U_dcore_U_sub_fifo_n55), 
	.A(FE_PHN4321_U_dfifo_U_dcore_U_sub_fifo_n55));
   BUF_X32 FE_PHC1790_U_dfifo_U_dcore_U_sub_fifo_n79 (.Z(FE_PHN1790_U_dfifo_U_dcore_U_sub_fifo_n79), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n79));
   BUF_X32 FE_PHC1789_U_afifo_m_data_in_28_ (.Z(FE_PHN1789_U_afifo_m_data_in_28_), 
	.A(U_afifo_m_data_in[28]));
   BUF_X32 FE_PHC1788_U_dfifo_U_dcore_U_sub_fifo_n81 (.Z(FE_PHN1788_U_dfifo_U_dcore_U_sub_fifo_n81), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n81));
   BUF_X32 FE_PHC1787_U_dfifo_U_dcore_U_sub_fifo_n63 (.Z(FE_PHN1787_U_dfifo_U_dcore_U_sub_fifo_n63), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n63));
   BUF_X32 FE_PHC1786_U_afifo_m_data_in_19_ (.Z(FE_PHN1786_U_afifo_m_data_in_19_), 
	.A(U_afifo_m_data_in[19]));
   BUF_X32 FE_PHC1785_U_dfifo_U_dcore_U_sub_fifo_n62 (.Z(FE_PHN1785_U_dfifo_U_dcore_U_sub_fifo_n62), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n62));
   BUF_X32 FE_PHC1784_U_afifo_U_acore_U_sub_fifo_n268 (.Z(FE_PHN1784_U_afifo_U_acore_U_sub_fifo_n268), 
	.A(FE_PHN3837_U_afifo_U_acore_U_sub_fifo_n268));
   BUF_X32 FE_PHC1783_U_afifo_m_data_in_33_ (.Z(FE_PHN1783_U_afifo_m_data_in_33_), 
	.A(U_afifo_m_data_in[33]));
   BUF_X32 FE_PHC1782_U_dfifo_U_dcore_U_sub_fifo_n73 (.Z(FE_PHN1782_U_dfifo_U_dcore_U_sub_fifo_n73), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n73));
   BUF_X32 FE_PHC1781_U_dfifo_U_dcore_U_sub_fifo_n69 (.Z(FE_PHN1781_U_dfifo_U_dcore_U_sub_fifo_n69), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n69));
   BUF_X32 FE_PHC1780_U_dfifo_U_dcore_U_sub_fifo_n329 (.Z(FE_PHN1780_U_dfifo_U_dcore_U_sub_fifo_n329), 
	.A(FE_PHN3809_U_dfifo_U_dcore_U_sub_fifo_n329));
   BUF_X32 FE_PHC1779_U_dfifo_U_dcore_U_sub_fifo_n78 (.Z(FE_PHN1779_U_dfifo_U_dcore_U_sub_fifo_n78), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n78));
   BUF_X32 FE_PHC1778_U_dfifo_U_dcore_U_sub_fifo_n65 (.Z(FE_PHN1778_U_dfifo_U_dcore_U_sub_fifo_n65), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n65));
   BUF_X32 FE_PHC1777_n25 (.Z(FE_PHN1777_n25), 
	.A(n25));
   BUF_X32 FE_PHC1776_U_dfifo_U_dcore_U_sub_fifo_n71 (.Z(FE_PHN1776_U_dfifo_U_dcore_U_sub_fifo_n71), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n71));
   BUF_X32 FE_PHC1775_U_dfifo_U_dcore_U_sub_fifo_n70 (.Z(FE_PHN1775_U_dfifo_U_dcore_U_sub_fifo_n70), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n70));
   BUF_X32 FE_PHC1774_U_dfifo_U_dcore_U_sub_fifo_n59 (.Z(FE_PHN1774_U_dfifo_U_dcore_U_sub_fifo_n59), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n59));
   BUF_X32 FE_PHC1773_U_dfifo_U_dcore_U_sub_fifo_n64 (.Z(FE_PHN1773_U_dfifo_U_dcore_U_sub_fifo_n64), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n64));
   BUF_X32 FE_PHC1772_U_dfifo_U_dcore_U_sub_fifo_n72 (.Z(FE_PHN1772_U_dfifo_U_dcore_U_sub_fifo_n72), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n72));
   BUF_X32 FE_PHC1771_U_dfifo_U_dcore_U_sub_fifo_n60 (.Z(FE_PHN1771_U_dfifo_U_dcore_U_sub_fifo_n60), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n60));
   BUF_X32 FE_PHC1770_U_dfifo_U_dcore_U_sub_fifo_n338 (.Z(FE_PHN1770_U_dfifo_U_dcore_U_sub_fifo_n338), 
	.A(FE_PHN4832_U_dfifo_U_dcore_U_sub_fifo_n338));
   BUF_X32 FE_PHC1769_U_afifo_m_data_in_20_ (.Z(FE_PHN1769_U_afifo_m_data_in_20_), 
	.A(U_afifo_m_data_in[20]));
   BUF_X32 FE_PHC1768_U_dfifo_U_dcore_U_sub_fifo_n61 (.Z(FE_PHN1768_U_dfifo_U_dcore_U_sub_fifo_n61), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n61));
   BUF_X32 FE_PHC1767_U_dfifo_U_dcore_U_sub_fifo_n58 (.Z(FE_PHN1767_U_dfifo_U_dcore_U_sub_fifo_n58), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n58));
   BUF_X32 FE_PHC1766_U_dfifo_U_dcore_U_sub_fifo_n68 (.Z(FE_PHN1766_U_dfifo_U_dcore_U_sub_fifo_n68), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n68));
   BUF_X32 FE_PHC1765_U_dfifo_U_dcore_U_sub_fifo_n66 (.Z(FE_PHN1765_U_dfifo_U_dcore_U_sub_fifo_n66), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n66));
   BUF_X32 FE_PHC1764_U_dfifo_U_dcore_U_sub_fifo_n67 (.Z(FE_PHN1764_U_dfifo_U_dcore_U_sub_fifo_n67), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n67));
   BUF_X32 FE_PHC1763_U_afifo_m_data_in_31_ (.Z(FE_PHN1763_U_afifo_m_data_in_31_), 
	.A(U_afifo_m_data_in[31]));
   BUF_X32 FE_PHC1762_n39 (.Z(FE_PHN1762_n39), 
	.A(n39));
   BUF_X32 FE_PHC1761_U_dfifo_U_dcore_U_sub_fifo_n344 (.Z(FE_PHN1761_U_dfifo_U_dcore_U_sub_fifo_n344), 
	.A(FE_PHN4770_U_dfifo_U_dcore_U_sub_fifo_n344));
   BUF_X32 FE_PHC1760_U_dfifo_U_dcore_U_sub_fifo_n76 (.Z(FE_PHN1760_U_dfifo_U_dcore_U_sub_fifo_n76), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n76));
   BUF_X32 FE_PHC1758_U_dfifo_U_dcore_U_sub_fifo_n332 (.Z(FE_PHN1758_U_dfifo_U_dcore_U_sub_fifo_n332), 
	.A(FE_PHN3677_U_dfifo_U_dcore_U_sub_fifo_n332));
   BUF_X32 FE_PHC1757_U_afifo_f_core_ready (.Z(FE_PHN1757_U_afifo_f_core_ready), 
	.A(U_afifo_f_core_ready));
   BUF_X32 FE_PHC1756_U_dfifo_U_dcore_U_sub_fifo_n339 (.Z(FE_PHN1756_U_dfifo_U_dcore_U_sub_fifo_n339), 
	.A(FE_PHN3705_U_dfifo_U_dcore_U_sub_fifo_n339));
   BUF_X32 FE_PHC1755_U_dfifo_U_dcore_U_sub_fifo_n74 (.Z(FE_PHN1755_U_dfifo_U_dcore_U_sub_fifo_n74), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n74));
   BUF_X32 FE_PHC1754_U_dfifo_U_dcore_U_sub_fifo_n75 (.Z(FE_PHN1754_U_dfifo_U_dcore_U_sub_fifo_n75), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n75));
   BUF_X32 FE_PHC1753_U_dfifo_U_dcore_U_sub_fifo_n77 (.Z(FE_PHN1753_U_dfifo_U_dcore_U_sub_fifo_n77), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n77));
   BUF_X32 FE_PHC1752_U_dfifo_U_dcore_U_sub_fifo_n336 (.Z(FE_PHN1752_U_dfifo_U_dcore_U_sub_fifo_n336), 
	.A(FE_PHN3649_U_dfifo_U_dcore_U_sub_fifo_n336));
   BUF_X32 FE_PHC1750_U_afifo_m_data_in_30_ (.Z(FE_PHN1750_U_afifo_m_data_in_30_), 
	.A(U_afifo_m_data_in[30]));
   BUF_X32 FE_PHC1749_U_afifo_m_data_in_21_ (.Z(FE_PHN1749_U_afifo_m_data_in_21_), 
	.A(U_afifo_m_data_in[21]));
   BUF_X32 FE_PHC1691_U_afifo_n10 (.Z(FE_PHN1691_U_afifo_n10), 
	.A(U_afifo_n10));
   BUF_X32 FE_PHC1689_n29 (.Z(FE_PHN1689_n29), 
	.A(n29));
   BUF_X32 FE_PHC1688_U_afifo_m_data_in_24_ (.Z(FE_PHN1688_U_afifo_m_data_in_24_), 
	.A(U_afifo_m_data_in[24]));
   BUF_X32 FE_PHC1687_U_afifo_m_data_in_2_ (.Z(FE_PHN1687_U_afifo_m_data_in_2_), 
	.A(U_afifo_m_data_in[2]));
   BUF_X32 FE_PHC1686_U_afifo_m_data_in_43_ (.Z(FE_PHN1686_U_afifo_m_data_in_43_), 
	.A(U_afifo_m_data_in[43]));
   BUF_X32 FE_PHC1685_U_afifo_m_data_in_23_ (.Z(FE_PHN1685_U_afifo_m_data_in_23_), 
	.A(U_afifo_m_data_in[23]));
   BUF_X32 FE_PHC1684_U_ctl_n120 (.Z(FE_PHN1684_U_ctl_n120), 
	.A(FE_PHN3203_U_ctl_n120));
   BUF_X32 FE_PHC1681_U_ctl_n117 (.Z(FE_PHN1681_U_ctl_n117), 
	.A(FE_PHN3207_U_ctl_n117));
   BUF_X32 FE_PHC1680_U_afifo_m_data_in_49_ (.Z(FE_PHN1680_U_afifo_m_data_in_49_), 
	.A(FE_PHN3471_U_afifo_m_data_in_49_));
   BUF_X32 FE_PHC1679_U_rbuf_n82 (.Z(FE_PHN1679_U_rbuf_n82), 
	.A(FE_PHN3281_U_rbuf_n82));
   BUF_X32 FE_PHC1678_U_rbuf_n84 (.Z(FE_PHN1678_U_rbuf_n84), 
	.A(FE_PHN3280_U_rbuf_n84));
   BUF_X32 FE_PHC1677_U_rbuf_n85 (.Z(FE_PHN1677_U_rbuf_n85), 
	.A(FE_PHN3279_U_rbuf_n85));
   BUF_X32 FE_PHC1676_U_rbuf_n71 (.Z(FE_PHN1676_U_rbuf_n71), 
	.A(FE_PHN3272_U_rbuf_n71));
   BUF_X32 FE_PHC1675_U_ctl_n421 (.Z(FE_PHN1675_U_ctl_n421), 
	.A(U_ctl_n421));
   BUF_X16 FE_PHC1660_U_dfifo_U_dcore_n_empty (.Z(FE_PHN1660_U_dfifo_U_dcore_n_empty), 
	.A(U_dfifo_U_dcore_n_empty));
   BUF_X32 FE_PHC1650_U_dfifo_U_dcore_n169 (.Z(FE_PHN1650_U_dfifo_U_dcore_n169), 
	.A(U_dfifo_U_dcore_n169));
   BUF_X32 FE_PHC1635_U_afifo_U_acore_U_sub_fifo_n323 (.Z(FE_PHN1635_U_afifo_U_acore_U_sub_fifo_n323), 
	.A(U_afifo_U_acore_U_sub_fifo_n323));
   BUF_X32 FE_PHC1630_U_dfifo_U_dcore_n145 (.Z(FE_PHN1630_U_dfifo_U_dcore_n145), 
	.A(FE_PHN4780_U_dfifo_U_dcore_n145));
   BUF_X32 FE_PHC1622_U_afifo_m_data_in_15_ (.Z(FE_PHN1622_U_afifo_m_data_in_15_), 
	.A(U_afifo_m_data_in[15]));
   BUF_X32 FE_PHC1621_U_afifo_m_data_in_17_ (.Z(FE_PHN1621_U_afifo_m_data_in_17_), 
	.A(U_afifo_m_data_in[17]));
   BUF_X32 FE_PHC1620_U_afifo_m_data_in_16_ (.Z(FE_PHN1620_U_afifo_m_data_in_16_), 
	.A(U_afifo_m_data_in[16]));
   BUF_X32 FE_PHC1619_U_afifo_n14 (.Z(FE_PHN1619_U_afifo_n14), 
	.A(U_afifo_n14));
   BUF_X32 FE_PHC1618_U_afifo_m_data_in_14_ (.Z(FE_PHN1618_U_afifo_m_data_in_14_), 
	.A(FE_PHN3225_U_afifo_m_data_in_14_));
   BUF_X32 FE_PHC1616_U_afifo_m_data_in_48_ (.Z(FE_PHN1616_U_afifo_m_data_in_48_), 
	.A(U_afifo_m_data_in[48]));
   BUF_X32 FE_PHC1611_U_ctl_n137 (.Z(FE_PHN1611_U_ctl_n137), 
	.A(FE_PHN3150_U_ctl_n137));
   BUF_X32 FE_PHC1609_U_ctl_n140 (.Z(FE_PHN1609_U_ctl_n140), 
	.A(FE_PHN3149_U_ctl_n140));
   BUF_X32 FE_PHC1607_U_afifo_n5 (.Z(FE_PHN1607_U_afifo_n5), 
	.A(U_afifo_n5));
   BUF_X32 FE_PHC1605_U_ctl_n118 (.Z(FE_PHN1605_U_ctl_n118), 
	.A(U_ctl_n118));
   BUF_X32 FE_PHC1604_U_ctl_n106 (.Z(FE_PHN1604_U_ctl_n106), 
	.A(FE_PHN3144_U_ctl_n106));
   BUF_X32 FE_PHC1595_U_dfifo_U_dcore_U_sub_fifo_count_0_ (.Z(FE_PHN1595_U_dfifo_U_dcore_U_sub_fifo_count_0_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_count_0_));
   BUF_X32 FE_PHC1592_U_afifo_U_acore_U_sub_fifo_out_ptr_0_ (.Z(FE_PHN1592_U_afifo_U_acore_U_sub_fifo_out_ptr_0_), 
	.A(U_afifo_U_acore_U_sub_fifo_out_ptr_0_));
   BUF_X8 FE_PHC1591_U_dfifo_U_dcore_U_sub_fifo_n242 (.Z(FE_PHN1591_U_dfifo_U_dcore_U_sub_fifo_n242), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n242));
   BUF_X32 FE_PHC1584_U_dfifo_U_dcore_U_sub_fifo_n18 (.Z(FE_PHN1584_U_dfifo_U_dcore_U_sub_fifo_n18), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n18));
   BUF_X32 FE_PHC1579_U_dfifo_U_dcore_n168 (.Z(FE_PHN1579_U_dfifo_U_dcore_n168), 
	.A(U_dfifo_U_dcore_n168));
   BUF_X32 FE_PHC1564_U_afifo_U_acore_n186 (.Z(FE_PHN1564_U_afifo_U_acore_n186), 
	.A(U_afifo_U_acore_n186));
   BUF_X32 FE_PHC1563_U_afifo_U_acore_n192 (.Z(FE_PHN1563_U_afifo_U_acore_n192), 
	.A(U_afifo_U_acore_n192));
   BUF_X32 FE_PHC1562_U_dfifo_U_dcore_n186 (.Z(FE_PHN1562_U_dfifo_U_dcore_n186), 
	.A(FE_PHN3338_U_dfifo_U_dcore_n186));
   BUF_X32 FE_PHC1561_U_afifo_U_acore_n205 (.Z(FE_PHN1561_U_afifo_U_acore_n205), 
	.A(U_afifo_U_acore_n205));
   BUF_X32 FE_PHC1560_U_afifo_U_acore_n175 (.Z(FE_PHN1560_U_afifo_U_acore_n175), 
	.A(U_afifo_U_acore_n175));
   BUF_X32 FE_PHC1558_U_afifo_U_acore_n190 (.Z(FE_PHN1558_U_afifo_U_acore_n190), 
	.A(U_afifo_U_acore_n190));
   BUF_X32 FE_PHC1556_U_dfifo_U_dcore_U_sub_fifo_n83 (.Z(FE_PHN1556_U_dfifo_U_dcore_U_sub_fifo_n83), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n83));
   BUF_X32 FE_PHC1554_U_afifo_U_acore_n179 (.Z(FE_PHN1554_U_afifo_U_acore_n179), 
	.A(U_afifo_U_acore_n179));
   BUF_X32 FE_PHC1553_U_afifo_U_acore_U_sub_fifo_n209 (.Z(FE_PHN1553_U_afifo_U_acore_U_sub_fifo_n209), 
	.A(FE_PHN5153_U_afifo_U_acore_U_sub_fifo_n209));
   BUF_X32 FE_PHC1552_U_afifo_U_acore_n80 (.Z(FE_PHN1552_U_afifo_U_acore_n80), 
	.A(U_afifo_U_acore_n80));
   BUF_X32 FE_PHC1550_U_dfifo_U_dcore_n193 (.Z(FE_PHN1550_U_dfifo_U_dcore_n193), 
	.A(FE_PHN3351_U_dfifo_U_dcore_n193));
   BUF_X32 FE_PHC1547_U_dfifo_U_dcore_n194 (.Z(FE_PHN1547_U_dfifo_U_dcore_n194), 
	.A(FE_PHN3417_U_dfifo_U_dcore_n194));
   BUF_X32 FE_PHC1546_U_dfifo_U_dcore_U_sub_fifo_n125 (.Z(FE_PHN1546_U_dfifo_U_dcore_U_sub_fifo_n125), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n125));
   BUF_X32 FE_PHC1545_U_dfifo_U_dcore_U_sub_fifo_n123 (.Z(FE_PHN1545_U_dfifo_U_dcore_U_sub_fifo_n123), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n123));
   BUF_X32 FE_PHC1544_U_dfifo_U_dcore_n201 (.Z(FE_PHN1544_U_dfifo_U_dcore_n201), 
	.A(U_dfifo_U_dcore_n201));
   BUF_X32 FE_PHC1543_U_dfifo_U_dcore_U_sub_fifo_n120 (.Z(FE_PHN1543_U_dfifo_U_dcore_U_sub_fifo_n120), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n120));
   BUF_X32 FE_PHC1542_U_dfifo_U_dcore_U_sub_fifo_n122 (.Z(FE_PHN1542_U_dfifo_U_dcore_U_sub_fifo_n122), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n122));
   BUF_X32 FE_PHC1541_U_dfifo_U_dcore_U_sub_fifo_n118 (.Z(FE_PHN1541_U_dfifo_U_dcore_U_sub_fifo_n118), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n118));
   BUF_X32 FE_PHC1540_U_dfifo_U_dcore_U_sub_fifo_n124 (.Z(FE_PHN1540_U_dfifo_U_dcore_U_sub_fifo_n124), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n124));
   BUF_X32 FE_PHC1539_U_dfifo_U_dcore_U_sub_fifo_n119 (.Z(FE_PHN1539_U_dfifo_U_dcore_U_sub_fifo_n119), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n119));
   BUF_X32 FE_PHC1527_U_afifo_n152 (.Z(FE_PHN1527_U_afifo_n152), 
	.A(U_afifo_n152));
   BUF_X32 FE_PHC1525_n17 (.Z(FE_PHN1525_n17), 
	.A(n17));
   BUF_X32 FE_PHC1515_U_afifo_m_data_in_29_ (.Z(FE_PHN1515_U_afifo_m_data_in_29_), 
	.A(U_afifo_m_data_in[29]));
   BUF_X32 FE_PHC1513_U_afifo_m_data_in_38_ (.Z(FE_PHN1513_U_afifo_m_data_in_38_), 
	.A(U_afifo_m_data_in[38]));
   BUF_X32 FE_PHC1511_U_ctl_n130 (.Z(FE_PHN1511_U_ctl_n130), 
	.A(FE_PHN3151_U_ctl_n130));
   BUF_X32 FE_PHC1510_U_ctl_n128 (.Z(FE_PHN1510_U_ctl_n128), 
	.A(FE_PHN3146_U_ctl_n128));
   BUF_X32 FE_PHC1509_U_ctl_n129 (.Z(FE_PHN1509_U_ctl_n129), 
	.A(FE_PHN3148_U_ctl_n129));
   BUF_X32 FE_PHC1507_U_ctl_n131 (.Z(FE_PHN1507_U_ctl_n131), 
	.A(FE_PHN3147_U_ctl_n131));
   BUF_X32 FE_PHC1506_U_ctl_n394 (.Z(FE_PHN1506_U_ctl_n394), 
	.A(U_ctl_n394));
   BUF_X32 FE_PHC1505_U_ctl_n119 (.Z(FE_PHN1505_U_ctl_n119), 
	.A(FE_PHN3095_U_ctl_n119));
   BUF_X8 FE_PHC1498_U_dfifo_U_dcore_n203 (.Z(FE_PHN1498_U_dfifo_U_dcore_n203), 
	.A(U_dfifo_U_dcore_n203));
   BUF_X32 FE_PHC1474_U_afifo_U_acore_U_sub_fifo_n315 (.Z(FE_PHN1474_U_afifo_U_acore_U_sub_fifo_n315), 
	.A(FE_PHN5037_U_afifo_U_acore_U_sub_fifo_n315));
   BUF_X32 FE_PHC1471_U_afifo_U_acore_U_sub_fifo_n324 (.Z(FE_PHN1471_U_afifo_U_acore_U_sub_fifo_n324), 
	.A(U_afifo_U_acore_U_sub_fifo_n324));
   BUF_X32 FE_PHC1467_U_dfifo_U_dcore_n188 (.Z(FE_PHN1467_U_dfifo_U_dcore_n188), 
	.A(FE_PHN3334_U_dfifo_U_dcore_n188));
   BUF_X32 FE_PHC1466_U_dfifo_U_dcore_n187 (.Z(FE_PHN1466_U_dfifo_U_dcore_n187), 
	.A(U_dfifo_U_dcore_n187));
   BUF_X32 FE_PHC1465_U_dfifo_U_dcore_n192 (.Z(FE_PHN1465_U_dfifo_U_dcore_n192), 
	.A(FE_PHN3368_U_dfifo_U_dcore_n192));
   BUF_X32 FE_PHC1464_U_dfifo_U_dcore_n191 (.Z(FE_PHN1464_U_dfifo_U_dcore_n191), 
	.A(FE_PHN3329_U_dfifo_U_dcore_n191));
   BUF_X32 FE_PHC1460_U_dfifo_U_dcore_U_sub_fifo_n447 (.Z(FE_PHN1460_U_dfifo_U_dcore_U_sub_fifo_n447), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n447));
   BUF_X32 FE_PHC1459_U_dfifo_U_dcore_n189 (.Z(FE_PHN1459_U_dfifo_U_dcore_n189), 
	.A(FE_PHN3341_U_dfifo_U_dcore_n189));
   BUF_X32 FE_PHC1458_U_dfifo_U_dcore_n190 (.Z(FE_PHN1458_U_dfifo_U_dcore_n190), 
	.A(U_dfifo_U_dcore_n190));
   BUF_X32 FE_PHC1454_U_dfifo_U_dcore_n197 (.Z(FE_PHN1454_U_dfifo_U_dcore_n197), 
	.A(FE_PHN3332_U_dfifo_U_dcore_n197));
   BUF_X32 FE_PHC1453_U_dfifo_U_dcore_n196 (.Z(FE_PHN1453_U_dfifo_U_dcore_n196), 
	.A(U_dfifo_U_dcore_n196));
   BUF_X32 FE_PHC1452_U_dfifo_U_dcore_n195 (.Z(FE_PHN1452_U_dfifo_U_dcore_n195), 
	.A(FE_PHN3398_U_dfifo_U_dcore_n195));
   BUF_X32 FE_PHC1451_U_dfifo_U_dcore_n198 (.Z(FE_PHN1451_U_dfifo_U_dcore_n198), 
	.A(U_dfifo_U_dcore_n198));
   BUF_X32 FE_PHC1446_U_dfifo_U_dcore_n173 (.Z(FE_PHN1446_U_dfifo_U_dcore_n173), 
	.A(U_dfifo_U_dcore_n173));
   BUF_X32 FE_PHC1443_U_dfifo_U_dcore_n182 (.Z(FE_PHN1443_U_dfifo_U_dcore_n182), 
	.A(FE_PHN3339_U_dfifo_U_dcore_n182));
   BUF_X32 FE_PHC1442_U_dfifo_U_dcore_n172 (.Z(FE_PHN1442_U_dfifo_U_dcore_n172), 
	.A(U_dfifo_U_dcore_n172));
   BUF_X32 FE_PHC1441_U_dfifo_U_dcore_n181 (.Z(FE_PHN1441_U_dfifo_U_dcore_n181), 
	.A(FE_PHN3354_U_dfifo_U_dcore_n181));
   BUF_X32 FE_PHC1440_U_dfifo_U_dcore_n174 (.Z(FE_PHN1440_U_dfifo_U_dcore_n174), 
	.A(U_dfifo_U_dcore_n174));
   BUF_X32 FE_PHC1439_U_dfifo_U_dcore_n171 (.Z(FE_PHN1439_U_dfifo_U_dcore_n171), 
	.A(U_dfifo_U_dcore_n171));
   BUF_X32 FE_PHC1438_U_dfifo_U_dcore_n176 (.Z(FE_PHN1438_U_dfifo_U_dcore_n176), 
	.A(FE_PHN3358_U_dfifo_U_dcore_n176));
   BUF_X32 FE_PHC1437_U_dfifo_U_dcore_n175 (.Z(FE_PHN1437_U_dfifo_U_dcore_n175), 
	.A(U_dfifo_U_dcore_n175));
   BUF_X32 FE_PHC1436_U_dfifo_U_dcore_n179 (.Z(FE_PHN1436_U_dfifo_U_dcore_n179), 
	.A(FE_PHN3330_U_dfifo_U_dcore_n179));
   BUF_X32 FE_PHC1435_U_dfifo_U_dcore_n184 (.Z(FE_PHN1435_U_dfifo_U_dcore_n184), 
	.A(FE_PHN3363_U_dfifo_U_dcore_n184));
   BUF_X32 FE_PHC1434_U_dfifo_U_dcore_n183 (.Z(FE_PHN1434_U_dfifo_U_dcore_n183), 
	.A(U_dfifo_U_dcore_n183));
   BUF_X32 FE_PHC1432_n13 (.Z(FE_PHN1432_n13), 
	.A(n13));
   BUF_X16 FE_PHC1423_U_dfifo_U_dcore_m_sf_full (.Z(FE_PHN1423_U_dfifo_U_dcore_m_sf_full), 
	.A(U_dfifo_U_dcore_m_sf_full));
   BUF_X32 FE_PHC1422_U_dfifo_U_dcore_U_sub_fifo_count_1_ (.Z(FE_PHN1422_U_dfifo_U_dcore_U_sub_fifo_count_1_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_count_1_));
   BUF_X32 FE_PHC1417_U_dfifo_U_dcore_f_buf_data_1_ (.Z(FE_PHN1417_U_dfifo_U_dcore_f_buf_data_1_), 
	.A(U_dfifo_U_dcore_f_buf_data_1_));
   CLKBUF_X1 FE_PHC1408_U_afifo_U_acore_n173 (.Z(FE_PHN1408_U_afifo_U_acore_n173), 
	.A(U_afifo_U_acore_n173));
   BUF_X32 FE_PHC1406_U_afifo_U_acore_n76 (.Z(FE_PHN1406_U_afifo_U_acore_n76), 
	.A(U_afifo_U_acore_n76));
   BUF_X32 FE_PHC1405_U_afifo_U_acore_n90 (.Z(FE_PHN1405_U_afifo_U_acore_n90), 
	.A(U_afifo_U_acore_n90));
   BUF_X32 FE_PHC1404_U_afifo_U_acore_n92 (.Z(FE_PHN1404_U_afifo_U_acore_n92), 
	.A(U_afifo_U_acore_n92));
   BUF_X32 FE_PHC1374_U_afifo_m_data_in_12_ (.Z(FE_PHN1374_U_afifo_m_data_in_12_), 
	.A(FE_PHN3213_U_afifo_m_data_in_12_));
   BUF_X32 FE_PHC1373_U_afifo_m_data_in_42_ (.Z(FE_PHN1373_U_afifo_m_data_in_42_), 
	.A(U_afifo_m_data_in[42]));
   BUF_X32 FE_PHC1370_U_ctl_n122 (.Z(FE_PHN1370_U_ctl_n122), 
	.A(FE_PHN3062_U_ctl_n122));
   BUF_X32 FE_PHC1368_U_ctl_n136 (.Z(FE_PHN1368_U_ctl_n136), 
	.A(FE_PHN3469_U_ctl_n136));
   CLKBUF_X1 FE_PHC1342_U_ctl_n101 (.Z(FE_PHN1342_U_ctl_n101), 
	.A(U_ctl_n101));
   BUF_X32 FE_PHC1332_U_afifo_U_acore_n141 (.Z(FE_PHN1332_U_afifo_U_acore_n141), 
	.A(U_afifo_U_acore_n141));
   BUF_X32 FE_PHC1330_U_afifo_U_acore_n142 (.Z(FE_PHN1330_U_afifo_U_acore_n142), 
	.A(FE_PHN3267_U_afifo_U_acore_n142));
   BUF_X32 FE_PHC1327_U_afifo_U_acore_n144 (.Z(FE_PHN1327_U_afifo_U_acore_n144), 
	.A(FE_PHN3265_U_afifo_U_acore_n144));
   BUF_X32 FE_PHC1325_U_afifo_U_acore_n138 (.Z(FE_PHN1325_U_afifo_U_acore_n138), 
	.A(FE_PHN3264_U_afifo_U_acore_n138));
   BUF_X32 FE_PHC1324_U_afifo_U_acore_n139 (.Z(FE_PHN1324_U_afifo_U_acore_n139), 
	.A(U_afifo_U_acore_n139));
   BUF_X16 FE_PHC1319_U_afifo_U_acore_n134 (.Z(FE_PHN1319_U_afifo_U_acore_n134), 
	.A(U_afifo_U_acore_n134));
   BUF_X32 FE_PHC1318_U_afifo_U_acore_n140 (.Z(FE_PHN1318_U_afifo_U_acore_n140), 
	.A(U_afifo_U_acore_n140));
   BUF_X32 FE_PHC1317_U_afifo_U_acore_n136 (.Z(FE_PHN1317_U_afifo_U_acore_n136), 
	.A(U_afifo_U_acore_n136));
   BUF_X16 FE_PHC1316_U_afifo_U_acore_n135 (.Z(FE_PHN1316_U_afifo_U_acore_n135), 
	.A(U_afifo_U_acore_n135));
   BUF_X16 FE_PHC1314_U_afifo_U_acore_n133 (.Z(FE_PHN1314_U_afifo_U_acore_n133), 
	.A(U_afifo_U_acore_n133));
   BUF_X32 FE_PHC1313_U_afifo_U_acore_n148 (.Z(FE_PHN1313_U_afifo_U_acore_n148), 
	.A(U_afifo_U_acore_n148));
   BUF_X32 FE_PHC1312_U_afifo_U_acore_n105 (.Z(FE_PHN1312_U_afifo_U_acore_n105), 
	.A(U_afifo_U_acore_n105));
   BUF_X32 FE_PHC1309_U_afifo_U_acore_n121 (.Z(FE_PHN1309_U_afifo_U_acore_n121), 
	.A(FE_PHN3254_U_afifo_U_acore_n121));
   BUF_X32 FE_PHC1308_U_afifo_U_acore_n137 (.Z(FE_PHN1308_U_afifo_U_acore_n137), 
	.A(U_afifo_U_acore_n137));
   BUF_X32 FE_PHC1307_U_afifo_U_acore_n110 (.Z(FE_PHN1307_U_afifo_U_acore_n110), 
	.A(U_afifo_U_acore_n110));
   BUF_X32 FE_PHC1305_U_afifo_U_acore_n151 (.Z(FE_PHN1305_U_afifo_U_acore_n151), 
	.A(U_afifo_U_acore_n151));
   BUF_X32 FE_PHC1304_U_afifo_U_acore_n115 (.Z(FE_PHN1304_U_afifo_U_acore_n115), 
	.A(FE_PHN3253_U_afifo_U_acore_n115));
   BUF_X32 FE_PHC1302_U_afifo_U_acore_n118 (.Z(FE_PHN1302_U_afifo_U_acore_n118), 
	.A(U_afifo_U_acore_n118));
   BUF_X32 FE_PHC1301_U_afifo_U_acore_n147 (.Z(FE_PHN1301_U_afifo_U_acore_n147), 
	.A(FE_PHN3251_U_afifo_U_acore_n147));
   BUF_X32 FE_PHC1298_U_afifo_U_acore_n111 (.Z(FE_PHN1298_U_afifo_U_acore_n111), 
	.A(U_afifo_U_acore_n111));
   BUF_X32 FE_PHC1297_U_afifo_U_acore_n114 (.Z(FE_PHN1297_U_afifo_U_acore_n114), 
	.A(U_afifo_U_acore_n114));
   BUF_X32 FE_PHC1296_U_afifo_U_acore_n152 (.Z(FE_PHN1296_U_afifo_U_acore_n152), 
	.A(U_afifo_U_acore_n152));
   BUF_X32 FE_PHC1293_U_afifo_U_acore_n112 (.Z(FE_PHN1293_U_afifo_U_acore_n112), 
	.A(U_afifo_U_acore_n112));
   BUF_X32 FE_PHC1290_U_afifo_U_acore_n149 (.Z(FE_PHN1290_U_afifo_U_acore_n149), 
	.A(U_afifo_U_acore_n149));
   BUF_X32 FE_PHC1289_U_afifo_U_acore_n109 (.Z(FE_PHN1289_U_afifo_U_acore_n109), 
	.A(U_afifo_U_acore_n109));
   BUF_X32 FE_PHC1286_U_afifo_U_acore_n108 (.Z(FE_PHN1286_U_afifo_U_acore_n108), 
	.A(U_afifo_U_acore_n108));
   BUF_X32 FE_PHC1285_U_afifo_U_acore_n117 (.Z(FE_PHN1285_U_afifo_U_acore_n117), 
	.A(U_afifo_U_acore_n117));
   BUF_X32 FE_PHC1284_U_afifo_U_acore_n146 (.Z(FE_PHN1284_U_afifo_U_acore_n146), 
	.A(U_afifo_U_acore_n146));
   BUF_X32 FE_PHC1282_U_afifo_U_acore_n154 (.Z(FE_PHN1282_U_afifo_U_acore_n154), 
	.A(U_afifo_U_acore_n154));
   BUF_X32 FE_PHC1281_U_afifo_U_acore_n130 (.Z(FE_PHN1281_U_afifo_U_acore_n130), 
	.A(U_afifo_U_acore_n130));
   BUF_X32 FE_PHC1280_U_afifo_U_acore_n107 (.Z(FE_PHN1280_U_afifo_U_acore_n107), 
	.A(U_afifo_U_acore_n107));
   BUF_X32 FE_PHC1278_U_afifo_U_acore_n106 (.Z(FE_PHN1278_U_afifo_U_acore_n106), 
	.A(U_afifo_U_acore_n106));
   BUF_X32 FE_PHC1277_U_afifo_U_acore_n113 (.Z(FE_PHN1277_U_afifo_U_acore_n113), 
	.A(U_afifo_U_acore_n113));
   BUF_X32 FE_PHC1276_U_afifo_U_acore_n150 (.Z(FE_PHN1276_U_afifo_U_acore_n150), 
	.A(U_afifo_U_acore_n150));
   BUF_X32 FE_PHC1274_U_afifo_U_acore_n126 (.Z(FE_PHN1274_U_afifo_U_acore_n126), 
	.A(U_afifo_U_acore_n126));
   BUF_X32 FE_PHC1273_U_afifo_U_acore_n128 (.Z(FE_PHN1273_U_afifo_U_acore_n128), 
	.A(U_afifo_U_acore_n128));
   BUF_X32 FE_PHC1272_U_afifo_U_acore_n116 (.Z(FE_PHN1272_U_afifo_U_acore_n116), 
	.A(U_afifo_U_acore_n116));
   BUF_X32 FE_PHC1270_U_afifo_U_acore_n131 (.Z(FE_PHN1270_U_afifo_U_acore_n131), 
	.A(U_afifo_U_acore_n131));
   BUF_X32 FE_PHC1267_U_afifo_U_acore_n127 (.Z(FE_PHN1267_U_afifo_U_acore_n127), 
	.A(U_afifo_U_acore_n127));
   BUF_X32 FE_PHC1266_U_afifo_U_acore_n120 (.Z(FE_PHN1266_U_afifo_U_acore_n120), 
	.A(U_afifo_U_acore_n120));
   BUF_X32 FE_PHC1265_U_afifo_U_acore_n145 (.Z(FE_PHN1265_U_afifo_U_acore_n145), 
	.A(U_afifo_U_acore_n145));
   BUF_X32 FE_PHC1264_U_afifo_U_acore_n132 (.Z(FE_PHN1264_U_afifo_U_acore_n132), 
	.A(U_afifo_U_acore_n132));
   BUF_X32 FE_PHC1263_U_afifo_U_acore_n124 (.Z(FE_PHN1263_U_afifo_U_acore_n124), 
	.A(U_afifo_U_acore_n124));
   BUF_X32 FE_PHC1261_U_afifo_U_acore_n129 (.Z(FE_PHN1261_U_afifo_U_acore_n129), 
	.A(U_afifo_U_acore_n129));
   BUF_X32 FE_PHC1260_U_afifo_U_acore_n123 (.Z(FE_PHN1260_U_afifo_U_acore_n123), 
	.A(U_afifo_U_acore_n123));
   BUF_X32 FE_PHC1259_U_afifo_U_acore_n122 (.Z(FE_PHN1259_U_afifo_U_acore_n122), 
	.A(U_afifo_U_acore_n122));
   BUF_X32 FE_PHC1258_U_afifo_U_acore_n125 (.Z(FE_PHN1258_U_afifo_U_acore_n125), 
	.A(U_afifo_U_acore_n125));
   BUF_X32 FE_PHC1257_U_afifo_U_acore_n119 (.Z(FE_PHN1257_U_afifo_U_acore_n119), 
	.A(U_afifo_U_acore_n119));
   BUF_X32 FE_PHC1250_U_dfifo_U_dcore_n200 (.Z(FE_PHN1250_U_dfifo_U_dcore_n200), 
	.A(FE_PHN3438_U_dfifo_U_dcore_n200));
   BUF_X32 FE_PHC1248_U_dfifo_U_dcore_n199 (.Z(FE_PHN1248_U_dfifo_U_dcore_n199), 
	.A(U_dfifo_U_dcore_n199));
   BUF_X32 FE_PHC1246_U_dfifo_U_dcore_n170 (.Z(FE_PHN1246_U_dfifo_U_dcore_n170), 
	.A(U_dfifo_U_dcore_n170));
   BUF_X32 FE_PHC1245_U_dfifo_U_dcore_n177 (.Z(FE_PHN1245_U_dfifo_U_dcore_n177), 
	.A(U_dfifo_U_dcore_n177));
   BUF_X32 FE_PHC1244_U_dfifo_U_dcore_n185 (.Z(FE_PHN1244_U_dfifo_U_dcore_n185), 
	.A(U_dfifo_U_dcore_n185));
   BUF_X32 FE_PHC1239_U_afifo_m_data_in_5_ (.Z(FE_PHN1239_U_afifo_m_data_in_5_), 
	.A(U_afifo_m_data_in[5]));
   BUF_X32 FE_PHC1238_U_afifo_m_data_in_4_ (.Z(FE_PHN1238_U_afifo_m_data_in_4_), 
	.A(FE_PHN3210_U_afifo_m_data_in_4_));
   BUF_X32 FE_PHC1233_U_ctl_n125 (.Z(FE_PHN1233_U_ctl_n125), 
	.A(FE_PHN3145_U_ctl_n125));
   BUF_X32 FE_PHC1232_U_ctl_n124 (.Z(FE_PHN1232_U_ctl_n124), 
	.A(FE_PHN3014_U_ctl_n124));
   BUF_X32 FE_PHC1231_U_rbuf_n88 (.Z(FE_PHN1231_U_rbuf_n88), 
	.A(U_rbuf_n88));
   BUF_X32 FE_PHC1229_U_ctl_n138 (.Z(FE_PHN1229_U_ctl_n138), 
	.A(FE_PHN3042_U_ctl_n138));
   CLKBUF_X1 FE_PHC1226_U_ctl_n102 (.Z(FE_PHN1226_U_ctl_n102), 
	.A(U_ctl_n102));
   BUF_X8 FE_PHC1225_U_ctl_n104 (.Z(FE_PHN1225_U_ctl_n104), 
	.A(U_ctl_n104));
   BUF_X32 FE_PHC1223_U_afifo_U_acore_U_sub_fifo_n171 (.Z(FE_PHN1223_U_afifo_U_acore_U_sub_fifo_n171), 
	.A(U_afifo_U_acore_U_sub_fifo_n171));
   BUF_X32 FE_PHC1197_U_afifo_U_acore_n72 (.Z(FE_PHN1197_U_afifo_U_acore_n72), 
	.A(U_afifo_U_acore_n72));
   BUF_X32 FE_PHC1194_U_afifo_U_acore_n74 (.Z(FE_PHN1194_U_afifo_U_acore_n74), 
	.A(U_afifo_U_acore_n74));
   BUF_X32 FE_PHC1193_U_afifo_U_acore_n88 (.Z(FE_PHN1193_U_afifo_U_acore_n88), 
	.A(U_afifo_U_acore_n88));
   BUF_X32 FE_PHC1192_U_afifo_U_acore_n68 (.Z(FE_PHN1192_U_afifo_U_acore_n68), 
	.A(U_afifo_U_acore_n68));
   BUF_X32 FE_PHC1191_U_afifo_U_acore_n78 (.Z(FE_PHN1191_U_afifo_U_acore_n78), 
	.A(U_afifo_U_acore_n78));
   BUF_X32 FE_PHC1190_U_afifo_U_acore_n84 (.Z(FE_PHN1190_U_afifo_U_acore_n84), 
	.A(U_afifo_U_acore_n84));
   BUF_X32 FE_PHC1189_U_afifo_U_acore_n167 (.Z(FE_PHN1189_U_afifo_U_acore_n167), 
	.A(U_afifo_U_acore_n167));
   BUF_X32 FE_PHC1188_U_afifo_U_acore_n86 (.Z(FE_PHN1188_U_afifo_U_acore_n86), 
	.A(U_afifo_U_acore_n86));
   BUF_X32 FE_PHC1187_U_afifo_U_acore_n82 (.Z(FE_PHN1187_U_afifo_U_acore_n82), 
	.A(U_afifo_U_acore_n82));
   BUF_X32 FE_PHC1186_U_afifo_U_acore_n70 (.Z(FE_PHN1186_U_afifo_U_acore_n70), 
	.A(U_afifo_U_acore_n70));
   BUF_X32 FE_PHC1184_U_dfifo_U_dcore_U_sub_fifo_n452 (.Z(FE_PHN1184_U_dfifo_U_dcore_U_sub_fifo_n452), 
	.A(FE_PHN4745_U_dfifo_U_dcore_U_sub_fifo_n452));
   BUF_X32 FE_PHC1182_U_dfifo_U_dcore_n143 (.Z(FE_PHN1182_U_dfifo_U_dcore_n143), 
	.A(FE_PHN3756_U_dfifo_U_dcore_n143));
   BUF_X32 FE_PHC1181_U_dfifo_U_dcore_n149 (.Z(FE_PHN1181_U_dfifo_U_dcore_n149), 
	.A(U_dfifo_U_dcore_n149));
   BUF_X32 FE_PHC1180_U_dfifo_U_dcore_n146 (.Z(FE_PHN1180_U_dfifo_U_dcore_n146), 
	.A(FE_PHN3655_U_dfifo_U_dcore_n146));
   BUF_X32 FE_PHC1179_U_dfifo_U_dcore_n142 (.Z(FE_PHN1179_U_dfifo_U_dcore_n142), 
	.A(U_dfifo_U_dcore_n142));
   BUF_X32 FE_PHC1178_U_afifo_m_data_in_32_ (.Z(FE_PHN1178_U_afifo_m_data_in_32_), 
	.A(U_afifo_m_data_in[32]));
   BUF_X32 FE_PHC1162_U_ctl_n139 (.Z(FE_PHN1162_U_ctl_n139), 
	.A(FE_PHN3269_U_ctl_n139));
   BUF_X32 FE_PHC1132_U_dfifo_n3 (.Z(FE_PHN1132_U_dfifo_n3), 
	.A(FE_PHN3284_U_dfifo_n3));
   BUF_X32 FE_PHC1125_U_dfifo_U_dcore_n180 (.Z(FE_PHN1125_U_dfifo_U_dcore_n180), 
	.A(FE_PHN3364_U_dfifo_U_dcore_n180));
   BUF_X32 FE_PHC1115_U_rbuf_n86 (.Z(FE_PHN1115_U_rbuf_n86), 
	.A(FE_PHN2998_U_rbuf_n86));
   BUF_X32 FE_PHC1114_U_rbuf_n79 (.Z(FE_PHN1114_U_rbuf_n79), 
	.A(FE_PHN2997_U_rbuf_n79));
   BUF_X32 FE_PHC1113_U_afifo_n49 (.Z(FE_PHN1113_U_afifo_n49), 
	.A(U_afifo_n49));
   BUF_X32 FE_PHC1112_U_rbuf_n75 (.Z(FE_PHN1112_U_rbuf_n75), 
	.A(FE_PHN2996_U_rbuf_n75));
   BUF_X32 FE_PHC1111_U_rbuf_n83 (.Z(FE_PHN1111_U_rbuf_n83), 
	.A(FE_PHN3025_U_rbuf_n83));
   BUF_X32 FE_PHC1110_U_rbuf_n80 (.Z(FE_PHN1110_U_rbuf_n80), 
	.A(FE_PHN3019_U_rbuf_n80));
   BUF_X32 FE_PHC1109_U_rbuf_n72 (.Z(FE_PHN1109_U_rbuf_n72), 
	.A(FE_PHN3023_U_rbuf_n72));
   BUF_X32 FE_PHC1108_U_rbuf_n77 (.Z(FE_PHN1108_U_rbuf_n77), 
	.A(FE_PHN3021_U_rbuf_n77));
   BUF_X32 FE_PHC1107_U_ctl_n134 (.Z(FE_PHN1107_U_ctl_n134), 
	.A(FE_PHN3154_U_ctl_n134));
   BUF_X32 FE_PHC1106_U_ctl_n133 (.Z(FE_PHN1106_U_ctl_n133), 
	.A(FE_PHN3155_U_ctl_n133));
   BUF_X32 FE_PHC1105_U_rbuf_n74 (.Z(FE_PHN1105_U_rbuf_n74), 
	.A(FE_PHN3015_U_rbuf_n74));
   BUF_X32 FE_PHC1104_U_rbuf_n78 (.Z(FE_PHN1104_U_rbuf_n78), 
	.A(FE_PHN2949_U_rbuf_n78));
   CLKBUF_X1 FE_PHC1102_U_ctl_n103 (.Z(FE_PHN1102_U_ctl_n103), 
	.A(U_ctl_n103));
   BUF_X8 FE_PHC1100_U_afifo_U_acore_U_sub_fifo_n325 (.Z(FE_PHN1100_U_afifo_U_acore_U_sub_fifo_n325), 
	.A(U_afifo_U_acore_U_sub_fifo_n325));
   BUF_X32 FE_PHC1084_U_dfifo_U_dcore_n154 (.Z(FE_PHN1084_U_dfifo_U_dcore_n154), 
	.A(FE_PHN4926_U_dfifo_U_dcore_n154));
   CLKBUF_X1 FE_PHC1079_U_ctl_n400 (.Z(FE_PHN1079_U_ctl_n400), 
	.A(U_ctl_n400));
   BUF_X32 FE_PHC1075_U_rbuf_n63 (.Z(FE_PHN1075_U_rbuf_n63), 
	.A(FE_PHN3027_U_rbuf_n63));
   BUF_X32 FE_PHC1074_U_rbuf_n64 (.Z(FE_PHN1074_U_rbuf_n64), 
	.A(FE_PHN3026_U_rbuf_n64));
   BUF_X32 FE_PHC1073_U_rbuf_n59 (.Z(FE_PHN1073_U_rbuf_n59), 
	.A(FE_PHN3022_U_rbuf_n59));
   BUF_X32 FE_PHC1072_U_rbuf_n65 (.Z(FE_PHN1072_U_rbuf_n65), 
	.A(FE_PHN3024_U_rbuf_n65));
   BUF_X32 FE_PHC1071_U_rbuf_n67 (.Z(FE_PHN1071_U_rbuf_n67), 
	.A(FE_PHN3007_U_rbuf_n67));
   BUF_X32 FE_PHC1070_U_rbuf_n60 (.Z(FE_PHN1070_U_rbuf_n60), 
	.A(FE_PHN3020_U_rbuf_n60));
   BUF_X32 FE_PHC1069_U_rbuf_n56 (.Z(FE_PHN1069_U_rbuf_n56), 
	.A(FE_PHN3008_U_rbuf_n56));
   BUF_X32 FE_PHC1068_U_rbuf_n61 (.Z(FE_PHN1068_U_rbuf_n61), 
	.A(FE_PHN3006_U_rbuf_n61));
   BUF_X32 FE_PHC1067_U_rbuf_n57 (.Z(FE_PHN1067_U_rbuf_n57), 
	.A(FE_PHN3004_U_rbuf_n57));
   BUF_X32 FE_PHC1066_U_rbuf_n70 (.Z(FE_PHN1066_U_rbuf_n70), 
	.A(FE_PHN3005_U_rbuf_n70));
   BUF_X32 FE_PHC1065_U_rbuf_n58 (.Z(FE_PHN1065_U_rbuf_n58), 
	.A(FE_PHN3003_U_rbuf_n58));
   BUF_X32 FE_PHC1049_U_afifo_U_acore_U_sub_fifo_n11 (.Z(FE_PHN1049_U_afifo_U_acore_U_sub_fifo_n11), 
	.A(U_afifo_U_acore_U_sub_fifo_n11));
   BUF_X32 FE_PHC1039_U_rbuf_n73 (.Z(FE_PHN1039_U_rbuf_n73), 
	.A(FE_PHN2999_U_rbuf_n73));
   CLKBUF_X1 FE_PHC1036_U_ctl_f_hiu_terminate (.Z(FE_PHN1036_U_ctl_f_hiu_terminate), 
	.A(U_ctl_f_hiu_terminate));
   BUF_X32 FE_PHC1027_U_afifo_n2 (.Z(FE_PHN1027_U_afifo_n2), 
	.A(U_afifo_n2));
   BUF_X32 FE_PHC1022_U_dfifo_U_dcore_n137 (.Z(FE_PHN1022_U_dfifo_U_dcore_n137), 
	.A(FE_PHN3130_U_dfifo_U_dcore_n137));
   BUF_X32 FE_PHC1021_U_dfifo_U_dcore_n138 (.Z(FE_PHN1021_U_dfifo_U_dcore_n138), 
	.A(FE_PHN3129_U_dfifo_U_dcore_n138));
   BUF_X32 FE_PHC1019_U_dfifo_U_dcore_n141 (.Z(FE_PHN1019_U_dfifo_U_dcore_n141), 
	.A(FE_PHN3131_U_dfifo_U_dcore_n141));
   BUF_X32 FE_PHC1018_U_dfifo_U_dcore_n134 (.Z(FE_PHN1018_U_dfifo_U_dcore_n134), 
	.A(U_dfifo_U_dcore_n134));
   BUF_X32 FE_PHC1011_U_ctl_n135 (.Z(FE_PHN1011_U_ctl_n135), 
	.A(FE_PHN3096_U_ctl_n135));
   BUF_X32 FE_PHC1002_U_ctl_n100 (.Z(FE_PHN1002_U_ctl_n100), 
	.A(U_ctl_n100));
   CLKBUF_X1 FE_PHC999_U_ctl_fr_wr_bcnt_0_ (.Z(FE_PHN999_U_ctl_fr_wr_bcnt_0_), 
	.A(U_ctl_fr_wr_bcnt_0_));
   CLKBUF_X1 FE_PHC993_U_afifo_U_acore_U_sub_fifo_n149 (.Z(FE_PHN993_U_afifo_U_acore_U_sub_fifo_n149), 
	.A(U_afifo_U_acore_U_sub_fifo_n149));
   BUF_X32 FE_PHC975_U_ctl_n132 (.Z(FE_PHN975_U_ctl_n132), 
	.A(FE_PHN2963_U_ctl_n132));
   BUF_X32 FE_PHC962_U_afifo_U_acore_n_afull (.Z(FE_PHN962_U_afifo_U_acore_n_afull), 
	.A(U_afifo_U_acore_n_afull));
   BUF_X32 FE_PHC956_U_dfifo_U_dcore_n147 (.Z(FE_PHN956_U_dfifo_U_dcore_n147), 
	.A(FE_PHN3716_U_dfifo_U_dcore_n147));
   BUF_X32 FE_PHC954_U_dfifo_U_dcore_n150 (.Z(FE_PHN954_U_dfifo_U_dcore_n150), 
	.A(FE_PHN4046_U_dfifo_U_dcore_n150));
   BUF_X32 FE_PHC950_U_afifo_n185 (.Z(FE_PHN950_U_afifo_n185), 
	.A(U_afifo_n185));
   BUF_X32 FE_PHC947_U_rbuf_n62 (.Z(FE_PHN947_U_rbuf_n62), 
	.A(FE_PHN2957_U_rbuf_n62));
   BUF_X32 FE_PHC930_U_rbuf_n76 (.Z(FE_PHN930_U_rbuf_n76), 
	.A(FE_PHN3017_U_rbuf_n76));
   BUF_X32 FE_PHC929_U_rbuf_n81 (.Z(FE_PHN929_U_rbuf_n81), 
	.A(FE_PHN3016_U_rbuf_n81));
   BUF_X32 FE_PHC923_U_dfifo_U_dcore_n167 (.Z(FE_PHN923_U_dfifo_U_dcore_n167), 
	.A(FE_PHN3266_U_dfifo_U_dcore_n167));
   BUF_X32 FE_PHC920_U_dfifo_U_dcore_n158 (.Z(FE_PHN920_U_dfifo_U_dcore_n158), 
	.A(U_dfifo_U_dcore_n158));
   BUF_X32 FE_PHC919_U_dfifo_U_dcore_n165 (.Z(FE_PHN919_U_dfifo_U_dcore_n165), 
	.A(U_dfifo_U_dcore_n165));
   BUF_X32 FE_PHC915_U_dfifo_U_dcore_n161 (.Z(FE_PHN915_U_dfifo_U_dcore_n161), 
	.A(U_dfifo_U_dcore_n161));
   BUF_X32 FE_PHC914_U_dfifo_U_dcore_n164 (.Z(FE_PHN914_U_dfifo_U_dcore_n164), 
	.A(U_dfifo_U_dcore_n164));
   BUF_X32 FE_PHC913_U_dfifo_U_dcore_n159 (.Z(FE_PHN913_U_dfifo_U_dcore_n159), 
	.A(U_dfifo_U_dcore_n159));
   BUF_X32 FE_PHC912_U_dfifo_U_dcore_n162 (.Z(FE_PHN912_U_dfifo_U_dcore_n162), 
	.A(U_dfifo_U_dcore_n162));
   BUF_X32 FE_PHC911_U_dfifo_U_dcore_n160 (.Z(FE_PHN911_U_dfifo_U_dcore_n160), 
	.A(U_dfifo_U_dcore_n160));
   BUF_X32 FE_PHC910_U_dfifo_U_dcore_n153 (.Z(FE_PHN910_U_dfifo_U_dcore_n153), 
	.A(FE_PHN5054_U_dfifo_U_dcore_n153));
   BUF_X32 FE_PHC909_U_dfifo_U_dcore_n152 (.Z(FE_PHN909_U_dfifo_U_dcore_n152), 
	.A(FE_PHN3965_U_dfifo_U_dcore_n152));
   BUF_X32 FE_PHC908_U_dfifo_U_dcore_n163 (.Z(FE_PHN908_U_dfifo_U_dcore_n163), 
	.A(U_dfifo_U_dcore_n163));
   BUF_X32 FE_PHC903_U_dfifo_U_dcore_n166 (.Z(FE_PHN903_U_dfifo_U_dcore_n166), 
	.A(U_dfifo_U_dcore_n166));
   BUF_X32 FE_PHC890_U_dfifo_U_dcore_n178 (.Z(FE_PHN890_U_dfifo_U_dcore_n178), 
	.A(FE_PHN3372_U_dfifo_U_dcore_n178));
   CLKBUF_X1 FE_PHC888_U_ctl_n150 (.Z(FE_PHN888_U_ctl_n150), 
	.A(U_ctl_n150));
   BUF_X32 FE_PHC885_U_ctl_n123 (.Z(FE_PHN885_U_ctl_n123), 
	.A(FE_PHN3270_U_ctl_n123));
   BUF_X32 FE_PHC876_U_rbuf_n68 (.Z(FE_PHN876_U_rbuf_n68), 
	.A(FE_PHN2934_U_rbuf_n68));
   BUF_X32 FE_PHC872_U_rbuf_n66 (.Z(FE_PHN872_U_rbuf_n66), 
	.A(FE_PHN2937_U_rbuf_n66));
   BUF_X16 FE_PHC868_U_afifo_U_acore_U_sub_fifo_n172 (.Z(FE_PHN868_U_afifo_U_acore_U_sub_fifo_n172), 
	.A(U_afifo_U_acore_U_sub_fifo_n172));
   BUF_X32 FE_PHC867_U_afifo_U_acore_U_sub_fifo_count_1_ (.Z(FE_PHN867_U_afifo_U_acore_U_sub_fifo_count_1_), 
	.A(U_afifo_U_acore_U_sub_fifo_count_1_));
   BUF_X32 FE_PHC861_U_dfifo_U_dcore_n144 (.Z(FE_PHN861_U_dfifo_U_dcore_n144), 
	.A(FE_PHN3789_U_dfifo_U_dcore_n144));
   BUF_X32 FE_PHC860_U_dfifo_U_dcore_n148 (.Z(FE_PHN860_U_dfifo_U_dcore_n148), 
	.A(FE_PHN3214_U_dfifo_U_dcore_n148));
   BUF_X32 FE_PHC858_U_dfifo_U_dcore_n140 (.Z(FE_PHN858_U_dfifo_U_dcore_n140), 
	.A(FE_PHN3428_U_dfifo_U_dcore_n140));
   BUF_X32 FE_PHC857_U_dfifo_U_dcore_n135 (.Z(FE_PHN857_U_dfifo_U_dcore_n135), 
	.A(FE_PHN3128_U_dfifo_U_dcore_n135));
   BUF_X32 FE_PHC848_U_ctl_n127 (.Z(FE_PHN848_U_ctl_n127), 
	.A(FE_PHN2933_U_ctl_n127));
   BUF_X32 FE_PHC828_U_rbuf_n69 (.Z(FE_PHN828_U_rbuf_n69), 
	.A(FE_PHN2938_U_rbuf_n69));
   BUF_X32 FE_PHC827_U_rbuf_n55 (.Z(FE_PHN827_U_rbuf_n55), 
	.A(FE_PHN2940_U_rbuf_n55));
   CLKBUF_X1 FE_PHC817_U_afifo_U_acore_n2 (.Z(FE_PHN817_U_afifo_U_acore_n2), 
	.A(U_afifo_U_acore_n2));
   BUF_X32 FE_PHC815_U_afifo_U_acore_n11 (.Z(FE_PHN815_U_afifo_U_acore_n11), 
	.A(U_afifo_U_acore_n11));
   BUF_X32 FE_PHC812_U_dfifo_U_dcore_n151 (.Z(FE_PHN812_U_dfifo_U_dcore_n151), 
	.A(FE_PHN4945_U_dfifo_U_dcore_n151));
   BUF_X32 FE_PHC811_U_dfifo_U_dcore_n156 (.Z(FE_PHN811_U_dfifo_U_dcore_n156), 
	.A(FE_PHN5016_U_dfifo_U_dcore_n156));
   BUF_X32 FE_PHC810_U_dfifo_U_dcore_n155 (.Z(FE_PHN810_U_dfifo_U_dcore_n155), 
	.A(FE_PHN4901_U_dfifo_U_dcore_n155));
   BUF_X32 FE_PHC809_U_dfifo_U_dcore_n157 (.Z(FE_PHN809_U_dfifo_U_dcore_n157), 
	.A(FE_PHN4928_U_dfifo_U_dcore_n157));
   BUF_X32 FE_PHC808_U_afifo_n65 (.Z(FE_PHN808_U_afifo_n65), 
	.A(U_afifo_n65));
   BUF_X32 FE_PHC798_U_afifo_n259 (.Z(FE_PHN798_U_afifo_n259), 
	.A(U_afifo_n259));
   BUF_X32 FE_PHC795_U_ctl_n180 (.Z(FE_PHN795_U_ctl_n180), 
	.A(U_ctl_n180));
   BUF_X32 FE_PHC789_U_dfifo_U_dcore_U_sub_fifo_n450 (.Z(FE_PHN789_U_dfifo_U_dcore_U_sub_fifo_n450), 
	.A(FE_PHN4812_U_dfifo_U_dcore_U_sub_fifo_n450));
   BUF_X32 FE_PHC785_U_dfifo_U_dcore_n136 (.Z(FE_PHN785_U_dfifo_U_dcore_n136), 
	.A(U_dfifo_U_dcore_n136));
   BUF_X32 FE_PHC784_U_dfifo_U_dcore_n139 (.Z(FE_PHN784_U_dfifo_U_dcore_n139), 
	.A(FE_PHN3132_U_dfifo_U_dcore_n139));
   BUF_X16 FE_PHC782_U_rbuf_n89 (.Z(FE_PHN782_U_rbuf_n89), 
	.A(U_rbuf_n89));
   BUF_X32 FE_PHC761_U_afifo_U_acore_f_push_req_n (.Z(FE_PHN761_U_afifo_U_acore_f_push_req_n), 
	.A(U_afifo_U_acore_f_push_req_n));
   BUF_X4 FE_PHC750_U_afifo_U_acore_n_obuf_empty (.Z(FE_PHN750_U_afifo_U_acore_n_obuf_empty), 
	.A(U_afifo_U_acore_n_obuf_empty));
   BUF_X32 FE_PHC747_U_ctl_n335 (.Z(FE_PHN747_U_ctl_n335), 
	.A(U_ctl_n335));
   BUF_X32 FE_PHC744_U_ctl_n105 (.Z(FE_PHN744_U_ctl_n105), 
	.A(FE_PHN3382_U_ctl_n105));
   BUF_X32 FE_PHC736_m_rb_overflow (.Z(FE_PHN736_m_rb_overflow), 
	.A(FE_PHN2924_m_rb_overflow));
   CLKBUF_X1 FE_PHC714_miu_burst_done (.Z(FE_PHN714_miu_burst_done), 
	.A(miu_burst_done));
   CLKBUF_X1 FE_PHC708_U_ctl_n418 (.Z(FE_PHN708_U_ctl_n418), 
	.A(U_ctl_n418));
   BUF_X32 FE_PHC700_U_ctl_n297 (.Z(FE_PHN700_U_ctl_n297), 
	.A(U_ctl_n297));
   BUF_X32 FE_PHC699_U_ctl_n382 (.Z(FE_PHN699_U_ctl_n382), 
	.A(FE_PHN2914_U_ctl_n382));
   BUF_X2 FE_PHC695_hsel_reg (.Z(FE_PHN695_hsel_reg), 
	.A(hsel_reg));
   BUF_X32 FE_PHC687_U_ctl_n422 (.Z(FE_PHN687_U_ctl_n422), 
	.A(U_ctl_n422));
   BUF_X32 FE_PHC682_U_ctl_n295 (.Z(FE_PHN682_U_ctl_n295), 
	.A(U_ctl_n295));
   BUF_X32 FE_PHC676_hiu_terminate (.Z(hiu_terminate), 
	.A(FE_PHN3002_hiu_terminate));
   BUF_X32 FE_PHC673_m_af_push1_n (.Z(FE_PHN673_m_af_push1_n), 
	.A(FE_PHN2908_m_af_push1_n));
   BUF_X4 FE_OFC296_n64 (.Z(FE_OFN296_n64), 
	.A(n64));
   BUF_X4 FE_OFC295_n61 (.Z(FE_OFN295_n61), 
	.A(n61));
   BUF_X4 FE_OFC294_n60 (.Z(FE_OFN294_n60), 
	.A(n60));
   BUF_X4 FE_OFC292_n56 (.Z(FE_OFN292_n56), 
	.A(n56));
   BUF_X4 FE_OFC291_n55 (.Z(FE_OFN291_n55), 
	.A(n55));
   BUF_X4 FE_OFC290_n53 (.Z(FE_OFN290_n53), 
	.A(n53));
   BUF_X4 FE_OFC289_U_dfifo_U_dcore_U_sub_fifo_n8 (.Z(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n8));
   BUF_X4 FE_OFC288_U_dfifo_U_dcore_U_sub_fifo_n9 (.Z(FE_OFN288_U_dfifo_U_dcore_U_sub_fifo_n9), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n9));
   BUF_X4 FE_OFC286_U_dfifo_U_dcore_U_sub_fifo_n10 (.Z(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n10));
   BUF_X4 FE_OFC282_U_dfifo_U_dcore_U_sub_fifo_n14 (.Z(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n14));
   BUF_X4 FE_OFC281_U_dfifo_U_dcore_U_sub_fifo_n15 (.Z(FE_OFN281_U_dfifo_U_dcore_U_sub_fifo_n15), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n15));
   BUF_X4 FE_OFC280_U_dfifo_U_dcore_U_sub_fifo_n16 (.Z(FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n16));
   BUF_X4 FE_OFC278_U_dfifo_U_dcore_U_sub_fifo_n231 (.Z(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n231));
   BUF_X4 FE_OFC275_U_dfifo_U_dcore_U_sub_fifo_n232 (.Z(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n232));
   BUF_X4 FE_OFC273_U_dfifo_U_dcore_U_sub_fifo_n234 (.Z(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n234));
   BUF_X4 FE_OFC271_U_dfifo_U_dcore_U_sub_fifo_n560 (.Z(FE_OFN271_U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n560));
   BUF_X4 FE_OFC267_U_dfifo_U_dcore_U_sub_fifo_n562 (.Z(FE_OFN267_U_dfifo_U_dcore_U_sub_fifo_n562), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n562));
   BUF_X4 FE_OFC265_U_dfifo_U_dcore_U_sub_fifo_n605 (.Z(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n605));
   BUF_X4 FE_OFC264_U_afifo_U_acore_U_sub_fifo_n152 (.Z(FE_OFN264_U_afifo_U_acore_U_sub_fifo_n152), 
	.A(U_afifo_U_acore_U_sub_fifo_n152));
   BUF_X4 FE_OFC263_U_afifo_U_acore_U_sub_fifo_n161 (.Z(FE_OFN263_U_afifo_U_acore_U_sub_fifo_n161), 
	.A(U_afifo_U_acore_U_sub_fifo_n161));
   BUF_X4 FE_OFC262_U_afifo_U_acore_U_sub_fifo_n161 (.Z(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.A(U_afifo_U_acore_U_sub_fifo_n161));
   BUF_X4 FE_OFC261_U_afifo_U_acore_U_sub_fifo_n163 (.Z(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A(U_afifo_U_acore_U_sub_fifo_n163));
   BUF_X4 FE_OFC260_U_afifo_U_acore_U_sub_fifo_n212 (.Z(FE_OFN260_U_afifo_U_acore_U_sub_fifo_n212), 
	.A(U_afifo_U_acore_U_sub_fifo_n212));
   BUF_X4 FE_OFC259_U_afifo_U_acore_U_sub_fifo_n369 (.Z(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.A(U_afifo_U_acore_U_sub_fifo_n369));
   BUF_X4 FE_OFC258_U_dfifo_U_dcore_n1 (.Z(FE_OFN258_U_dfifo_U_dcore_n1), 
	.A(U_dfifo_U_dcore_n1));
   BUF_X4 FE_OFC256_U_dfifo_U_dcore_n2 (.Z(FE_OFN256_U_dfifo_U_dcore_n2), 
	.A(U_dfifo_U_dcore_n2));
   BUF_X4 FE_OFC255_U_dfifo_U_dcore_n3 (.Z(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A(U_dfifo_U_dcore_n3));
   BUF_X4 FE_OFC252_U_dfifo_U_dcore_n127 (.Z(FE_OFN252_U_dfifo_U_dcore_n127), 
	.A(U_dfifo_U_dcore_n127));
   BUF_X4 FE_OFC250_U_afifo_U_acore_n1 (.Z(FE_OFN250_U_afifo_U_acore_n1), 
	.A(U_afifo_U_acore_n1));
   BUF_X4 FE_OFC247_U_afifo_U_acore_n211 (.Z(FE_OFN247_U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n211));
   BUF_X4 FE_OFC244_U_rbuf_n180 (.Z(FE_OFN244_U_rbuf_n180), 
	.A(U_rbuf_n180));
   BUF_X4 FE_OFC237_U_afifo_n54 (.Z(FE_OFN237_U_afifo_n54), 
	.A(U_afifo_n54));
   BUF_X4 FE_OFC236_U_afifo_n93 (.Z(FE_OFN236_U_afifo_n93), 
	.A(U_afifo_n98));
   BUF_X4 FE_OFC225_hiu_data_26_ (.Z(FE_OFN225_hiu_data_26_), 
	.A(hiu_data[26]));
   BUF_X4 FE_OFC210_hwrite_s (.Z(FE_OFN210_hwrite_s), 
	.A(hwrite));
   BUF_X4 FE_OFC207_U_afifo_U_acore_U_sub_fifo_n169 (.Z(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.A(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169));
   BUF_X4 FE_OFC206_U_afifo_U_acore_U_sub_fifo_n369 (.Z(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.A(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369));
   BUF_X4 FE_OFC203_U_afifo_U_acore_U_sub_fifo_n1 (.Z(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.A(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1));
   BUF_X4 FE_OFC202_U_afifo_U_acore_U_sub_fifo_n162 (.Z(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162), 
	.A(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   BUF_X4 FE_OFC197_U_afifo_U_acore_n38 (.Z(FE_OFN197_U_afifo_U_acore_n38), 
	.A(FE_OFN26_U_afifo_U_acore_n38));
   BUF_X4 FE_OFC196_HRESETn (.Z(FE_OFN196_HRESETn), 
	.A(FE_OFN28_HRESETn));
   BUF_X4 FE_OFC193_HRESETn (.Z(FE_OFN193_HRESETn), 
	.A(FE_OFN29_HRESETn));
   BUF_X4 FE_OFC176_HRESETn (.Z(FE_OFN176_HRESETn), 
	.A(FE_OFN42_HRESETn));
   BUF_X4 FE_OFC171_HRESETn (.Z(FE_OFN171_HRESETn), 
	.A(FE_OFN47_HRESETn));
   BUF_X4 FE_OFC170_HRESETn (.Z(FE_OFN170_HRESETn), 
	.A(FE_OFN47_HRESETn));
   BUF_X4 FE_OFC169_HRESETn (.Z(FE_OFN169_HRESETn), 
	.A(FE_OFN47_HRESETn));
   BUF_X4 FE_OFC168_HRESETn (.Z(FE_OFN168_HRESETn), 
	.A(FE_OFN47_HRESETn));
   BUF_X4 FE_OFC157_HRESETn (.Z(FE_OFN157_HRESETn), 
	.A(FE_OFN53_HRESETn));
   BUF_X4 FE_OFC156_HRESETn (.Z(FE_OFN156_HRESETn), 
	.A(FE_OFN54_HRESETn));
   BUF_X4 FE_OFC153_HRESETn (.Z(FE_OFN153_HRESETn), 
	.A(FE_OFN55_HRESETn));
   BUF_X4 FE_OFC150_HRESETn (.Z(FE_OFN150_HRESETn), 
	.A(FE_OFN58_HRESETn));
   BUF_X4 FE_OFC149_HRESETn (.Z(FE_OFN149_HRESETn), 
	.A(FE_OFN58_HRESETn));
   BUF_X4 FE_OFC143_HRESETn (.Z(FE_OFN143_HRESETn), 
	.A(FE_OFN62_HRESETn));
   BUF_X4 FE_OFC136_HRESETn (.Z(FE_OFN136_HRESETn), 
	.A(FE_OFN67_HRESETn));
   CLKBUF_X3 FE_OFC69_HRESETn (.Z(FE_OFN69_HRESETn), 
	.A(FE_OFN62_HRESETn));
   BUF_X8 FE_OFC67_HRESETn (.Z(FE_OFN67_HRESETn), 
	.A(FE_OFN42_HRESETn));
   BUF_X8 FE_OFC62_HRESETn (.Z(FE_OFN62_HRESETn), 
	.A(FE_OFN42_HRESETn));
   BUF_X8 FE_OFC58_HRESETn (.Z(FE_OFN58_HRESETn), 
	.A(FE_OFN29_HRESETn));
   CLKBUF_X3 FE_OFC54_HRESETn (.Z(FE_OFN54_HRESETn), 
	.A(FE_OFN43_HRESETn));
   BUF_X8 FE_OFC47_HRESETn (.Z(FE_OFN47_HRESETn), 
	.A(FE_OFN32_HRESETn));
   INV_X8 FE_OFC32_HRESETn (.ZN(FE_OFN32_HRESETn), 
	.A(hresetn));
   BUF_X4 FE_OFC26_U_afifo_U_acore_n38 (.Z(FE_OFN26_U_afifo_U_acore_n38), 
	.A(U_afifo_U_acore_n38));
   BUF_X4 FE_OFC7_U_afifo_U_acore_U_sub_fifo_n162 (.Z(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162), 
	.A(U_afifo_U_acore_U_sub_fifo_n162));
   BUF_X4 FE_OFC6_U_afifo_U_acore_U_sub_fifo_n1 (.Z(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.A(U_afifo_U_acore_U_sub_fifo_n1));
   BUF_X4 FE_OFC4_U_afifo_U_acore_U_sub_fifo_n169 (.Z(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.A(U_afifo_U_acore_U_sub_fifo_n169));
   NAND2_X2 U_afifo_U299 (.ZN(U_afifo_n259), 
	.A2(U_afifo_n153), 
	.A1(U_afifo_m_data_out_49));
   AND2_X4 U_afifo_U298 (.ZN(U_afifo_n156), 
	.A2(U_afifo_m_full), 
	.A1(U_afifo_m_pop_n));
   NAND2_X1 U_afifo_U297 (.ZN(U_afifo_n168), 
	.A2(U_afifo_m_afull), 
	.A1(U_afifo_m_pop_n));
   AOI22_X2 U_afifo_U293 (.ZN(U_afifo_n181), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN2161_U_afifo_f_data2_7_), 
	.A2(U_afifo_n98), 
	.A1(1'b0));
   INV_X4 U_afifo_U292 (.ZN(U_afifo_m_data_in[7]), 
	.A(U_afifo_n181));
   AOI21_X2 U_afifo_U291 (.ZN(U_afifo_n182), 
	.B2(U_afifo_n99), 
	.B1(1'b0), 
	.A(FE_PHN1527_U_afifo_n152));
   INV_X4 U_afifo_U290 (.ZN(U_afifo_m_data_in[8]), 
	.A(U_afifo_n182));
   OAI21_X2 U_afifo_U288 (.ZN(U_afifo_n51), 
	.B2(FE_PHN2567_U_afifo_n165), 
	.B1(1'b0), 
	.A(1'b1));
   OAI21_X2 U_afifo_U287 (.ZN(U_afifo_n16), 
	.B2(FE_PHN2638_U_afifo_n159), 
	.B1(1'b0), 
	.A(1'b1));
   OAI21_X2 U_afifo_U285 (.ZN(U_afifo_n52), 
	.B2(FE_PHN2575_U_afifo_n166), 
	.B1(1'b0), 
	.A(1'b1));
   OAI21_X2 U_afifo_U284 (.ZN(U_afifo_n17), 
	.B2(FE_PHN2558_U_afifo_n160), 
	.B1(1'b0), 
	.A(1'b1));
   NAND2_X2 U_afifo_U282 (.ZN(U_afifo_n173), 
	.A2(1'b1), 
	.A1(FE_PHN1881_U_afifo_f_data2_5_));
   NAND2_X2 U_afifo_U281 (.ZN(U_afifo_n154), 
	.A2(FE_PHN3390_U_afifo_n173), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U280 (.ZN(U_afifo_n3), 
	.B2(FE_PHN3481_U_afifo_n157), 
	.B1(FE_PHN1757_U_afifo_f_core_ready), 
	.A(1'b1));
   NAND2_X2 U_afifo_U279 (.ZN(U_afifo_n186), 
	.A2(FE_PHN1879_U_afifo_f_data2_0_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U278 (.ZN(U_afifo_n4), 
	.B2(U_afifo_n187), 
	.B1(1'b1), 
	.A(FE_PHN3458_U_afifo_n186));
   OAI21_X2 U_afifo_U276 (.ZN(U_afifo_n8), 
	.B2(FE_PHN2565_U_afifo_n191), 
	.B1(1'b0), 
	.A(1'b1));
   NAND2_X2 U_afifo_U275 (.ZN(U_afifo_n224), 
	.A2(FE_PHN1883_U_afifo_f_data2_31_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U274 (.ZN(U_afifo_n35), 
	.B2(U_afifo_n225), 
	.B1(1'b1), 
	.A(FE_PHN3403_U_afifo_n224));
   NAND2_X2 U_afifo_U273 (.ZN(U_afifo_n250), 
	.A2(FE_PHN1885_U_afifo_f_data2_44_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U272 (.ZN(U_afifo_n48), 
	.B2(1'b1), 
	.B1(1'b1), 
	.A(FE_PHN3400_U_afifo_n250));
   NAND2_X2 U_afifo_U271 (.ZN(U_afifo_n202), 
	.A2(FE_PHN1880_U_afifo_f_data2_20_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U270 (.ZN(U_afifo_n24), 
	.B2(U_afifo_n203), 
	.B1(1'b1), 
	.A(FE_PHN3441_U_afifo_n202));
   NAND2_X2 U_afifo_U269 (.ZN(U_afifo_n216), 
	.A2(FE_PHN1867_U_afifo_f_data2_27_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U268 (.ZN(U_afifo_n31), 
	.B2(U_afifo_n217), 
	.B1(1'b1), 
	.A(FE_PHN3393_U_afifo_n216));
   NAND2_X2 U_afifo_U267 (.ZN(U_afifo_n198), 
	.A2(FE_PHN1882_U_afifo_f_data2_18_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U266 (.ZN(U_afifo_n22), 
	.B2(U_ctl_n16), 
	.B1(1'b1), 
	.A(FE_PHN3435_U_afifo_n198));
   NAND2_X2 U_afifo_U265 (.ZN(U_afifo_n214), 
	.A2(FE_PHN1873_U_afifo_f_data2_26_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U264 (.ZN(U_afifo_n30), 
	.B2(U_afifo_n215), 
	.B1(1'b1), 
	.A(FE_PHN3388_U_afifo_n214));
   NAND2_X2 U_afifo_U263 (.ZN(U_afifo_n228), 
	.A2(FE_PHN1856_U_afifo_f_data2_33_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U262 (.ZN(U_afifo_n37), 
	.B2(U_afifo_n229), 
	.B1(1'b1), 
	.A(FE_PHN3385_U_afifo_n228));
   NAND2_X2 U_afifo_U261 (.ZN(U_afifo_n200), 
	.A2(FE_PHN1860_U_afifo_f_data2_19_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U260 (.ZN(U_afifo_n23), 
	.B2(U_afifo_n201), 
	.B1(1'b1), 
	.A(FE_PHN3397_U_afifo_n200));
   NAND2_X2 U_afifo_U259 (.ZN(U_afifo_n226), 
	.A2(FE_PHN1863_U_afifo_f_data2_32_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U258 (.ZN(U_afifo_n36), 
	.B2(U_afifo_n227), 
	.B1(1'b1), 
	.A(FE_PHN3422_U_afifo_n226));
   NAND2_X2 U_afifo_U257 (.ZN(U_afifo_n206), 
	.A2(FE_PHN1864_U_afifo_f_data2_22_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U256 (.ZN(U_afifo_n26), 
	.B2(U_afifo_n207), 
	.B1(1'b1), 
	.A(FE_PHN3420_U_afifo_n206));
   NAND2_X2 U_afifo_U255 (.ZN(U_afifo_n222), 
	.A2(FE_PHN1861_U_afifo_f_data2_30_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U254 (.ZN(U_afifo_n34), 
	.B2(U_afifo_n223), 
	.B1(1'b1), 
	.A(FE_PHN3392_U_afifo_n222));
   NAND2_X2 U_afifo_U253 (.ZN(U_afifo_n188), 
	.A2(FE_PHN1862_U_afifo_f_data2_2_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U252 (.ZN(U_afifo_n6), 
	.B2(hwrite), 
	.B1(1'b1), 
	.A(FE_PHN3425_U_afifo_n188));
   NAND2_X2 U_afifo_U251 (.ZN(U_afifo_n220), 
	.A2(FE_PHN1866_U_afifo_f_data2_29_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U250 (.ZN(U_afifo_n33), 
	.B2(U_afifo_n221), 
	.B1(1'b1), 
	.A(FE_PHN3429_U_afifo_n220));
   NAND2_X2 U_afifo_U249 (.ZN(U_afifo_n218), 
	.A2(FE_PHN1858_U_afifo_f_data2_28_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U248 (.ZN(U_afifo_n32), 
	.B2(U_afifo_n219), 
	.B1(1'b1), 
	.A(FE_PHN3404_U_afifo_n218));
   NAND2_X2 U_afifo_U247 (.ZN(U_afifo_n208), 
	.A2(FE_PHN1874_U_afifo_f_data2_23_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U246 (.ZN(U_afifo_n27), 
	.B2(U_afifo_n209), 
	.B1(1'b1), 
	.A(FE_PHN3436_U_afifo_n208));
   NAND2_X2 U_afifo_U245 (.ZN(U_afifo_n204), 
	.A2(FE_PHN1853_U_afifo_f_data2_21_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U244 (.ZN(U_afifo_n25), 
	.B2(U_afifo_n205), 
	.B1(1'b1), 
	.A(FE_PHN3413_U_afifo_n204));
   NAND2_X2 U_afifo_U243 (.ZN(U_afifo_n212), 
	.A2(FE_PHN1865_U_afifo_f_data2_25_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U242 (.ZN(U_afifo_n29), 
	.B2(U_afifo_n213), 
	.B1(1'b1), 
	.A(FE_PHN3439_U_afifo_n212));
   NAND2_X2 U_afifo_U241 (.ZN(U_afifo_n210), 
	.A2(FE_PHN1876_U_afifo_f_data2_24_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U240 (.ZN(U_afifo_n28), 
	.B2(U_afifo_n211), 
	.B1(1'b1), 
	.A(FE_PHN3434_U_afifo_n210));
   OAI21_X2 U_afifo_U238 (.ZN(U_afifo_n19), 
	.B2(U_afifo_n162), 
	.B1(1'b0), 
	.A(1'b1));
   OAI21_X2 U_afifo_U236 (.ZN(U_afifo_n18), 
	.B2(U_afifo_n161), 
	.B1(1'b0), 
	.A(1'b1));
   OAI21_X2 U_afifo_U234 (.ZN(U_afifo_n20), 
	.B2(U_afifo_n163), 
	.B1(1'b0), 
	.A(1'b1));
   NAND2_X2 U_afifo_U231 (.ZN(U_afifo_n234), 
	.A2(FE_PHN1859_U_afifo_f_data2_36_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U230 (.ZN(U_afifo_n40), 
	.B2(U_afifo_n235), 
	.B1(1'b1), 
	.A(FE_PHN3408_U_afifo_n234));
   NAND2_X2 U_afifo_U229 (.ZN(U_afifo_n238), 
	.A2(FE_PHN1886_U_afifo_f_data2_38_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U228 (.ZN(U_afifo_n42), 
	.B2(U_afifo_n239), 
	.B1(1'b1), 
	.A(FE_PHN3402_U_afifo_n238));
   NAND2_X2 U_afifo_U227 (.ZN(U_afifo_n246), 
	.A2(FE_PHN1884_U_afifo_f_data2_42_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U226 (.ZN(U_afifo_n46), 
	.B2(U_ctl_n227), 
	.B1(1'b1), 
	.A(FE_PHN3394_U_afifo_n246));
   NAND2_X2 U_afifo_U225 (.ZN(U_afifo_n248), 
	.A2(FE_PHN1872_U_afifo_f_data2_43_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U224 (.ZN(U_afifo_n47), 
	.B2(U_ctl_n230), 
	.B1(1'b1), 
	.A(FE_PHN3419_U_afifo_n248));
   NAND2_X2 U_afifo_U223 (.ZN(U_afifo_n230), 
	.A2(FE_PHN1857_U_afifo_f_data2_34_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U222 (.ZN(U_afifo_n38), 
	.B2(U_afifo_n231), 
	.B1(1'b1), 
	.A(FE_PHN3410_U_afifo_n230));
   NAND2_X2 U_afifo_U221 (.ZN(U_afifo_n240), 
	.A2(FE_PHN1871_U_afifo_f_data2_39_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U220 (.ZN(U_afifo_n43), 
	.B2(U_afifo_n241), 
	.B1(1'b1), 
	.A(FE_PHN3396_U_afifo_n240));
   NAND2_X2 U_afifo_U219 (.ZN(U_afifo_n244), 
	.A2(FE_PHN1817_U_afifo_f_data2_41_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U218 (.ZN(U_afifo_n45), 
	.B2(U_afifo_n245), 
	.B1(1'b1), 
	.A(FE_PHN3395_U_afifo_n244));
   NAND2_X2 U_afifo_U217 (.ZN(U_afifo_n232), 
	.A2(FE_PHN1870_U_afifo_f_data2_35_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U216 (.ZN(U_afifo_n39), 
	.B2(U_afifo_n233), 
	.B1(1'b1), 
	.A(FE_PHN3424_U_afifo_n232));
   NAND2_X2 U_afifo_U215 (.ZN(U_afifo_n242), 
	.A2(FE_PHN1869_U_afifo_f_data2_40_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U214 (.ZN(U_afifo_n44), 
	.B2(U_afifo_n243), 
	.B1(1'b1), 
	.A(FE_PHN3383_U_afifo_n242));
   NAND2_X2 U_afifo_U213 (.ZN(U_afifo_n236), 
	.A2(FE_PHN1878_U_afifo_f_data2_37_), 
	.A1(1'b1));
   OAI21_X2 U_afifo_U212 (.ZN(U_afifo_n41), 
	.B2(U_afifo_n237), 
	.B1(1'b1), 
	.A(FE_PHN3418_U_afifo_n236));
   NAND2_X2 U_afifo_U210 (.ZN(U_afifo_n171), 
	.A2(1'b1), 
	.A1(FE_PHN1877_U_afifo_f_data2_6_));
   NAND2_X2 U_afifo_U209 (.ZN(U_afifo_n155), 
	.A2(FE_PHN3381_U_afifo_n171), 
	.A1(1'b1));
   INV_X4 U_afifo_U208 (.ZN(U_afifo_n256), 
	.A(U_afifo_m_data_out_0_));
   NOR3_X2 U_afifo_U207 (.ZN(hiu_req[1]), 
	.A3(U_afifo_n256), 
	.A2(U_afifo_m_empty), 
	.A1(m_af_dummy_req));
   AOI21_X2 U_afifo_U206 (.ZN(m_af_ready), 
	.B2(U_afifo_f_push2_pending), 
	.B1(U_afifo_m_afull), 
	.A(U_afifo_n151));
   AOI22_X2 U_afifo_U205 (.ZN(U_afifo_n179), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1881_U_afifo_f_data2_5_), 
	.A2(U_afifo_n140), 
	.A1(m_af_data1_in_5_));
   INV_X4 U_afifo_U204 (.ZN(U_afifo_m_data_in[5]), 
	.A(U_afifo_n179));
   AOI22_X2 U_afifo_U203 (.ZN(U_afifo_n180), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1877_U_afifo_f_data2_6_), 
	.A2(FE_OFN236_U_afifo_n93), 
	.A1(1'b0));
   INV_X4 U_afifo_U202 (.ZN(U_afifo_m_data_in[6]), 
	.A(U_afifo_n180));
   OAI21_X2 U_afifo_U201 (.ZN(U_afifo_n_new_req), 
	.B2(U_afifo_n255), 
	.B1(U_afifo_m_aempty), 
	.A(U_afifo_n184));
   NAND2_X2 U_afifo_U200 (.ZN(U_afifo_n169), 
	.A2(U_afifo_n167), 
	.A1(U_afifo_n168));
   OAI21_X2 U_afifo_U199 (.ZN(U_afifo_n65), 
	.B2(U_afifo_n156), 
	.B1(FE_PHN950_U_afifo_n185), 
	.A(U_afifo_n169));
   NOR3_X2 U_afifo_U198 (.ZN(hiu_req[0]), 
	.A3(U_afifo_m_data_out_0_), 
	.A2(U_afifo_m_empty), 
	.A1(m_af_dummy_req));
   INV_X1 U_afifo_U197 (.ZN(U_afifo_n187), 
	.A(m_af_data1_in_0_));
   INV_X1 U_afifo_U196 (.ZN(U_afifo_n255), 
	.A(miu_burst_done));
   OAI21_X1 U_afifo_U195 (.ZN(U_afifo_n184), 
	.B2(U_afifo_m_empty), 
	.B1(miu_burst_done), 
	.A(FE_PHN950_U_afifo_n185));
   INV_X4 U_afifo_U194 (.ZN(m_af_dummy_req), 
	.A(FE_PHN798_U_afifo_n259));
   INV_X1 U_afifo_U189 (.ZN(U_afifo_n147), 
	.A(U_afifo_n54));
   INV_X1 U_afifo_U184 (.ZN(U_afifo_n140), 
	.A(U_afifo_n54));
   NAND2_X2 U_afifo_U182 (.ZN(U_afifo_n137), 
	.A2(FE_PHN1884_U_afifo_f_data2_42_), 
	.A1(U_afifo_n54));
   INV_X1 U_afifo_U156 (.ZN(U_afifo_n99), 
	.A(U_afifo_n54));
   INV_X1 U_afifo_U155 (.ZN(U_afifo_n98), 
	.A(U_afifo_n54));
   NAND2_X2 U_afifo_U145 (.ZN(U_afifo_n84), 
	.A2(FE_PHN1886_U_afifo_f_data2_38_), 
	.A1(U_afifo_n54));
   NAND2_X2 U_afifo_U139 (.ZN(U_afifo_n75), 
	.A2(FE_PHN1863_U_afifo_f_data2_32_), 
	.A1(FE_OFN237_U_afifo_n54));
   NAND2_X1 U_afifo_U125 (.ZN(U_afifo_n183), 
	.A2(U_afifo_f_push2_pending), 
	.A1(FE_PHN1757_U_afifo_f_core_ready));
   INV_X2 U_afifo_U123 (.ZN(U_afifo_n167), 
	.A(U_afifo_m_full));
   INV_X1 U_afifo_U122 (.ZN(U_afifo_n257), 
	.A(U_afifo_m_data_out_49));
   NAND2_X2 U_afifo_U121 (.ZN(U_afifo_m_pop_n), 
	.A2(FE_PHN798_U_afifo_n259), 
	.A1(miu_burst_done));
   OAI21_X1 U_afifo_U120 (.ZN(U_afifo_n2), 
	.B2(FE_PHN798_U_afifo_n259), 
	.B1(U_afifo_n255), 
	.A(U_afifo_n258));
   INV_X1 U_afifo_U116 (.ZN(U_afifo_n55), 
	.A(FE_PHN950_U_afifo_n185));
   NAND2_X2 U_afifo_U107 (.ZN(U_afifo_n85), 
	.A2(haddr[28]), 
	.A1(U_afifo_n147));
   AND2_X2 U_afifo_U103 (.ZN(U_afifo_m_data_in[45]), 
	.A2(haddr[0]), 
	.A1(U_afifo_n147));
   NAND2_X2 U_afifo_U96 (.ZN(U_afifo_n76), 
	.A2(haddr[22]), 
	.A1(U_afifo_n147));
   AND2_X2 U_afifo_U92 (.ZN(U_afifo_m_data_in[46]), 
	.A2(haddr[1]), 
	.A1(U_afifo_n140));
   AND2_X2 U_afifo_U91 (.ZN(U_afifo_m_data_in[11]), 
	.A2(U_afifo_n99), 
	.A1(m_af_data1_in_11_));
   NAND2_X2 U_afifo_U81 (.ZN(U_afifo_m_data_in[38]), 
	.A2(U_afifo_n84), 
	.A1(U_afifo_n85));
   NAND2_X2 U_afifo_U64 (.ZN(U_afifo_m_data_in[32]), 
	.A2(U_afifo_n75), 
	.A1(U_afifo_n76));
   NAND2_X2 U_afifo_U62 (.ZN(U_afifo_m_data_in[42]), 
	.A2(U_afifo_n137), 
	.A1(U_afifo_n138));
   AOI22_X2 U_afifo_U59 (.ZN(U_afifo_n192), 
	.B2(1'b1), 
	.B1(FE_PHN2161_U_afifo_f_data2_7_), 
	.A2(1'b0), 
	.A1(m_af_data2_in[7]));
   INV_X2 U_afifo_U58 (.ZN(U_afifo_n217), 
	.A(haddr[17]));
   INV_X2 U_afifo_U57 (.ZN(U_afifo_n205), 
	.A(haddr[11]));
   INV_X2 U_afifo_U56 (.ZN(U_afifo_n219), 
	.A(haddr[18]));
   INV_X2 U_afifo_U55 (.ZN(U_afifo_n207), 
	.A(haddr[12]));
   INV_X2 U_afifo_U54 (.ZN(U_afifo_n209), 
	.A(haddr[13]));
   INV_X2 U_afifo_U53 (.ZN(U_afifo_n201), 
	.A(haddr[9]));
   INV_X2 U_afifo_U52 (.ZN(U_afifo_n213), 
	.A(haddr[15]));
   INV_X2 U_afifo_U51 (.ZN(U_afifo_n215), 
	.A(haddr[16]));
   INV_X2 U_afifo_U50 (.ZN(U_afifo_n211), 
	.A(haddr[14]));
   INV_X2 U_afifo_U49 (.ZN(U_afifo_n203), 
	.A(haddr[10]));
   INV_X2 U_afifo_U48 (.ZN(U_afifo_n243), 
	.A(haddr[30]));
   INV_X2 U_afifo_U47 (.ZN(U_afifo_n245), 
	.A(haddr[31]));
   INV_X2 U_afifo_U46 (.ZN(U_afifo_n235), 
	.A(haddr[26]));
   INV_X2 U_afifo_U45 (.ZN(U_afifo_n237), 
	.A(haddr[27]));
   INV_X2 U_afifo_U44 (.ZN(U_afifo_n239), 
	.A(haddr[28]));
   INV_X2 U_afifo_U43 (.ZN(U_afifo_n241), 
	.A(haddr[29]));
   INV_X2 U_afifo_U42 (.ZN(U_afifo_n229), 
	.A(haddr[23]));
   INV_X2 U_afifo_U41 (.ZN(U_afifo_n225), 
	.A(haddr[21]));
   INV_X2 U_afifo_U40 (.ZN(U_afifo_n231), 
	.A(haddr[24]));
   INV_X2 U_afifo_U39 (.ZN(U_afifo_n223), 
	.A(haddr[20]));
   INV_X2 U_afifo_U38 (.ZN(U_afifo_n227), 
	.A(haddr[22]));
   INV_X2 U_afifo_U37 (.ZN(U_afifo_n233), 
	.A(haddr[25]));
   INV_X2 U_afifo_U36 (.ZN(U_afifo_n221), 
	.A(haddr[19]));
   OAI21_X1 U_afifo_U35 (.ZN(U_afifo_n258), 
	.B2(U_afifo_n257), 
	.B1(U_afifo_n255), 
	.A(FE_PHN3374_U_afifo_f_clr_pers));
   NAND2_X2 U_afifo_U33 (.ZN(U_afifo_n185), 
	.A2(U_afifo_n183), 
	.A1(U_afifo_n54));
   AND2_X2 U_afifo_U32 (.ZN(U_afifo_n152), 
	.A2(U_afifo_f_data2_8_), 
	.A1(U_afifo_n54));
   NAND2_X2 U_afifo_U29 (.ZN(U_afifo_n138), 
	.A2(hsize[0]), 
	.A1(U_afifo_n98));
   NOR2_X2 U_afifo_U28 (.ZN(U_afifo_m_data_in[49]), 
	.A2(FE_PHN3481_U_afifo_n157), 
	.A1(U_afifo_n54));
   INV_X4 U_afifo_U26 (.ZN(U_afifo_n54), 
	.A(U_afifo_n178));
   INV_X1 U_afifo_U25 (.ZN(U_afifo_m_data_in[13]), 
	.A(FE_PHN1113_U_afifo_n49));
   AOI22_X1 U_afifo_U24 (.ZN(U_afifo_n49), 
	.B2(m_af_data1_in_13_), 
	.B1(U_afifo_n178), 
	.A2(U_afifo_f_data2_13_), 
	.A1(U_afifo_n54));
   AOI22_X1 U_afifo_U22 (.ZN(U_afifo_n15), 
	.B2(U_afifo_n54), 
	.B1(U_afifo_f_data2_48_), 
	.A2(U_afifo_n147), 
	.A1(haddr[3]));
   INV_X1 U_afifo_U21 (.ZN(U_afifo_m_data_in[47]), 
	.A(FE_PHN1619_U_afifo_n14));
   AOI22_X1 U_afifo_U20 (.ZN(U_afifo_n14), 
	.B2(U_afifo_n54), 
	.B1(U_afifo_f_data2_47_), 
	.A2(U_afifo_n99), 
	.A1(haddr[2]));
   INV_X1 U_afifo_U19 (.ZN(U_afifo_m_data_in[14]), 
	.A(U_afifo_n13));
   AOI22_X1 U_afifo_U18 (.ZN(U_afifo_n13), 
	.B2(U_afifo_n54), 
	.B1(U_afifo_f_data2_14_), 
	.A2(U_afifo_n98), 
	.A1(haddr[4]));
   INV_X1 U_afifo_U17 (.ZN(U_afifo_m_data_in[15]), 
	.A(U_afifo_n11));
   AOI22_X1 U_afifo_U16 (.ZN(U_afifo_n11), 
	.B2(U_afifo_n54), 
	.B1(U_afifo_f_data2_15_), 
	.A2(U_afifo_n99), 
	.A1(haddr[5]));
   INV_X1 U_afifo_U15 (.ZN(U_afifo_m_data_in[18]), 
	.A(FE_PHN1691_U_afifo_n10));
   AOI22_X1 U_afifo_U14 (.ZN(U_afifo_n10), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1882_U_afifo_f_data2_18_), 
	.A2(U_afifo_n98), 
	.A1(haddr[8]));
   INV_X1 U_afifo_U13 (.ZN(U_afifo_m_data_in[43]), 
	.A(U_afifo_n9));
   AOI22_X1 U_afifo_U12 (.ZN(U_afifo_n9), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1872_U_afifo_f_data2_43_), 
	.A2(U_afifo_n98), 
	.A1(hsize[1]));
   INV_X1 U_afifo_U11 (.ZN(U_afifo_m_data_in[44]), 
	.A(U_afifo_n7));
   AOI22_X1 U_afifo_U10 (.ZN(U_afifo_n7), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1885_U_afifo_f_data2_44_), 
	.A2(U_afifo_n140), 
	.A1(1'b0));
   INV_X1 U_afifo_U9 (.ZN(U_afifo_m_data_in[0]), 
	.A(FE_PHN1607_U_afifo_n5));
   AOI22_X1 U_afifo_U8 (.ZN(U_afifo_n5), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1879_U_afifo_f_data2_0_), 
	.A2(U_afifo_n140), 
	.A1(m_af_data1_in_0_));
   INV_X1 U_afifo_U7 (.ZN(U_afifo_m_data_in[4]), 
	.A(U_afifo_n1));
   AOI22_X2 U_afifo_U6 (.ZN(U_afifo_n1), 
	.B2(m_af_data1_in_4_), 
	.B1(FE_OFN236_U_afifo_n93), 
	.A2(U_afifo_f_data2_4_), 
	.A1(U_afifo_n54));
   AND2_X4 U_afifo_U5 (.ZN(hiu_wrap_burst), 
	.A2(U_afifo_m_data_out_3), 
	.A1(FE_PHN798_U_afifo_n259));
   INV_X4 U_afifo_U3 (.ZN(U_afifo_n178), 
	.A(FE_PHN673_m_af_push1_n));
   DFFR_X2 U_afifo_f_data2_reg_8_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_n158), 
	.Q(U_afifo_f_data2_8_), 
	.D(U_afifo_n12), 
	.CK(HCLK__L5_N27));
   DFFR_X2 U_afifo_f_data2_reg_12_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_n159), 
	.Q(U_afifo_f_data2_12_), 
	.D(U_afifo_n16), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_f_data2_reg_13_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_n160), 
	.Q(U_afifo_f_data2_13_), 
	.D(FE_PHN5024_U_afifo_n17), 
	.CK(HCLK__L5_N27));
   DFFR_X2 U_afifo_f_data2_reg_47_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_n165), 
	.Q(U_afifo_f_data2_47_), 
	.D(U_afifo_n51), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_f_data2_reg_48_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_n166), 
	.Q(U_afifo_f_data2_48_), 
	.D(U_afifo_n52), 
	.CK(HCLK__L5_N27));
   DFFR_X2 U_afifo_f_data2_reg_4_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_n191), 
	.Q(U_afifo_f_data2_4_), 
	.D(U_afifo_n8), 
	.CK(HCLK__L5_N27));
   DFFS_X2 U_afifo_f_data2_reg_7_ (.SN(FE_OFN34_HRESETn), 
	.QN(U_afifo_f_data2_7_), 
	.D(FE_PHN4028_U_afifo_n192), 
	.CK(HCLK__L5_N27));
   DFFR_X1 U_afifo_f_new_req_reg (.RN(FE_OFN153_HRESETn), 
	.QN(m_af_new_req), 
	.D(FE_PHN3032_U_afifo_n_new_req), 
	.CK(HCLK__L5_N35));
   DFFS_X2 U_afifo_f_ready_reg (.SN(FE_OFN153_HRESETn), 
	.QN(U_afifo_n151), 
	.D(FE_PHN808_U_afifo_n65), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_afifo_f_clr_pers_reg (.RN(FE_OFN153_HRESETn), 
	.QN(U_afifo_n153), 
	.Q(U_afifo_f_clr_pers), 
	.D(FE_PHN1027_U_afifo_n2), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_afifo_f_push2_pending_reg (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_n157), 
	.Q(U_afifo_f_push2_pending), 
	.D(FE_PHN2133_U_afifo_n3), 
	.CK(HCLK__L5_N36));
   DFFS_X2 U_afifo_f_core_ready_reg (.SN(FE_OFN31_HRESETn), 
	.Q(U_afifo_f_core_ready), 
	.D(FE_PHN808_U_afifo_n65), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_f_data2_reg_0_ (.RN(FE_OFN34_HRESETn), 
	.Q(U_afifo_f_data2_0_), 
	.D(U_afifo_n4), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_f_data2_reg_2_ (.RN(FE_OFN34_HRESETn), 
	.Q(U_afifo_f_data2_2_), 
	.D(U_afifo_n6), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_f_data2_reg_5_ (.RN(FE_OFN34_HRESETn), 
	.Q(U_afifo_f_data2_5_), 
	.D(U_afifo_n154), 
	.CK(HCLK__L5_N27));
   DFFR_X1 U_afifo_f_data2_reg_6_ (.RN(FE_OFN34_HRESETn), 
	.Q(U_afifo_f_data2_6_), 
	.D(U_afifo_n155), 
	.CK(HCLK__L5_N27));
   DFFR_X1 U_afifo_f_data2_reg_14_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_n161), 
	.Q(U_afifo_f_data2_14_), 
	.D(FE_PHN2656_U_afifo_n18), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_f_data2_reg_15_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_n162), 
	.Q(U_afifo_f_data2_15_), 
	.D(FE_PHN2677_U_afifo_n19), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_f_data2_reg_16_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_n163), 
	.Q(U_afifo_f_data2_16_), 
	.D(FE_PHN2704_U_afifo_n20), 
	.CK(HCLK__L5_N27));
   DFFR_X1 U_afifo_f_data2_reg_17_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_n164), 
	.Q(U_afifo_f_data2_17_), 
	.D(U_afifo_n21), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_18_ (.RN(FE_OFN193_HRESETn), 
	.Q(U_afifo_f_data2_18_), 
	.D(U_afifo_n22), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_19_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_19_), 
	.D(U_afifo_n23), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_20_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_20_), 
	.D(U_afifo_n24), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_21_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_21_), 
	.D(U_afifo_n25), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_22_ (.RN(FE_OFN193_HRESETn), 
	.Q(U_afifo_f_data2_22_), 
	.D(U_afifo_n26), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_23_ (.RN(FE_OFN193_HRESETn), 
	.Q(U_afifo_f_data2_23_), 
	.D(U_afifo_n27), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_24_ (.RN(FE_OFN193_HRESETn), 
	.Q(U_afifo_f_data2_24_), 
	.D(U_afifo_n28), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_25_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_25_), 
	.D(U_afifo_n29), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_26_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_26_), 
	.D(U_afifo_n30), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_27_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_27_), 
	.D(U_afifo_n31), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_28_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_28_), 
	.D(U_afifo_n32), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_29_ (.RN(FE_OFN193_HRESETn), 
	.Q(U_afifo_f_data2_29_), 
	.D(U_afifo_n33), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_30_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_30_), 
	.D(U_afifo_n34), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_31_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_31_), 
	.D(U_afifo_n35), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_32_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_32_), 
	.D(U_afifo_n36), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_33_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_33_), 
	.D(U_afifo_n37), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_34_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_34_), 
	.D(U_afifo_n38), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_35_ (.RN(FE_OFN193_HRESETn), 
	.Q(U_afifo_f_data2_35_), 
	.D(U_afifo_n39), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_36_ (.RN(FE_OFN193_HRESETn), 
	.Q(U_afifo_f_data2_36_), 
	.D(U_afifo_n40), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_37_ (.RN(FE_OFN32_HRESETn), 
	.Q(U_afifo_f_data2_37_), 
	.D(U_afifo_n41), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_38_ (.RN(FE_OFN193_HRESETn), 
	.Q(U_afifo_f_data2_38_), 
	.D(U_afifo_n42), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_39_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_f_data2_39_), 
	.D(U_afifo_n43), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_40_ (.RN(FE_OFN32_HRESETn), 
	.Q(U_afifo_f_data2_40_), 
	.D(U_afifo_n44), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_41_ (.RN(FE_OFN32_HRESETn), 
	.Q(U_afifo_f_data2_41_), 
	.D(U_afifo_n45), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_42_ (.RN(FE_OFN34_HRESETn), 
	.Q(U_afifo_f_data2_42_), 
	.D(U_afifo_n46), 
	.CK(HCLK__L5_N27));
   DFFR_X1 U_afifo_f_data2_reg_43_ (.RN(FE_OFN32_HRESETn), 
	.Q(U_afifo_f_data2_43_), 
	.D(U_afifo_n47), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_f_data2_reg_44_ (.RN(FE_OFN32_HRESETn), 
	.Q(U_afifo_f_data2_44_), 
	.D(U_afifo_n48), 
	.CK(HCLK__L5_N39));
   OAI221_X1 U_dfifo_U26 (.ZN(U_dfifo_n3), 
	.C2(U_dfifo_n2), 
	.C1(U_ctl_n384), 
	.B2(U_dfifo_f_1st_half), 
	.B1(miu_pop_n), 
	.A(U_dfifo_m_data_out_1_));
   MUX2_X2 U_dfifo_U25 (.Z(hiu_data[8]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[8]), 
	.A(hiu_data[24]));
   MUX2_X2 U_dfifo_U24 (.Z(hiu_data[0]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[0]), 
	.A(hiu_data[16]));
   MUX2_X2 U_dfifo_U23 (.Z(hiu_data[9]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[9]), 
	.A(hiu_data[25]));
   MUX2_X2 U_dfifo_U22 (.Z(hiu_data[1]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[1]), 
	.A(hiu_data[17]));
   MUX2_X2 U_dfifo_U21 (.Z(hiu_data[10]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[10]), 
	.A(hiu_data[26]));
   MUX2_X2 U_dfifo_U20 (.Z(hiu_data[2]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[2]), 
	.A(hiu_data[18]));
   MUX2_X2 U_dfifo_U19 (.Z(hiu_data[12]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[12]), 
	.A(hiu_data[28]));
   MUX2_X2 U_dfifo_U18 (.Z(hiu_data[4]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[4]), 
	.A(hiu_data[20]));
   MUX2_X2 U_dfifo_U17 (.Z(hiu_data[11]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[11]), 
	.A(hiu_data[27]));
   MUX2_X2 U_dfifo_U16 (.Z(hiu_data[3]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[3]), 
	.A(hiu_data[19]));
   MUX2_X2 U_dfifo_U15 (.Z(hiu_data[13]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[13]), 
	.A(hiu_data[29]));
   MUX2_X2 U_dfifo_U14 (.Z(hiu_data[5]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[5]), 
	.A(hiu_data[21]));
   MUX2_X2 U_dfifo_U13 (.Z(hiu_data[15]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[15]), 
	.A(hiu_data[31]));
   MUX2_X2 U_dfifo_U12 (.Z(hiu_data[7]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[7]), 
	.A(hiu_data[23]));
   MUX2_X2 U_dfifo_U11 (.Z(hiu_data[14]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[14]), 
	.A(hiu_data[30]));
   MUX2_X2 U_dfifo_U10 (.Z(hiu_data[6]), 
	.S(U_dfifo_n4), 
	.B(U_dfifo_m_btm_data[6]), 
	.A(hiu_data[22]));
   NAND2_X2 U_dfifo_U8 (.ZN(U_dfifo_n4), 
	.A2(U_dfifo_n2), 
	.A1(U_dfifo_m_data_out_1_));
   AOI21_X2 U_dfifo_U7 (.ZN(U_dfifo_n5), 
	.B2(U_dfifo_m_data_out_1_), 
	.B1(U_dfifo_f_1st_half), 
	.A(miu_pop_n));
   AND2_X2 U_dfifo_U6 (.ZN(m_df_wr_term), 
	.A2(U_dfifo_m_data_out_0_), 
	.A1(U_dfifo_n5));
   AOI21_X2 U_dfifo_U5 (.ZN(m_df_ready), 
	.B2(m_df_push_n), 
	.B1(U_dfifo_m_afull), 
	.A(U_dfifo_m_full));
   DFFS_X2 U_dfifo_f_1st_half_reg (.SN(FE_OFN160_HRESETn), 
	.QN(U_dfifo_n2), 
	.Q(U_dfifo_f_1st_half), 
	.D(FE_PHN1132_U_dfifo_n3), 
	.CK(HCLK__L5_N6));
   INV_X4 U_rbuf_U215 (.ZN(U_rbuf_n177), 
	.A(U_rbuf_n161));
   AND3_X4 U_rbuf_U214 (.ZN(U_rbuf_n16), 
	.A3(U_rbuf_n160), 
	.A2(m_two_to_one), 
	.A1(n48));
   INV_X4 U_rbuf_U212 (.ZN(U_rbuf_n196), 
	.A(U_rbuf_n198));
   NOR2_X2 U_rbuf_U208 (.ZN(U_rbuf_n148), 
	.A2(U_rbuf_n17), 
	.A1(U_ctl_n324));
   NOR2_X2 U_rbuf_U207 (.ZN(U_rbuf_n154), 
	.A2(U_rbuf_n148), 
	.A1(miu_push_n));
   NAND2_X2 U_rbuf_U206 (.ZN(U_rbuf_n151), 
	.A2(U_rbuf_n154), 
	.A1(m_rb_pop_n));
   INV_X4 U_rbuf_U205 (.ZN(m_rb_overflow), 
	.A(U_rbuf_n151));
   NAND2_X2 U_rbuf_U204 (.ZN(U_rbuf_n125), 
	.A2(U_rbuf_n120), 
	.A1(m_double));
   NAND2_X2 U_rbuf_U203 (.ZN(U_rbuf_n126), 
	.A2(n48), 
	.A1(U_rbuf_n125));
   NAND2_X4 U_rbuf_U202 (.ZN(U_rbuf_n143), 
	.A2(U_rbuf_n126), 
	.A1(U_rbuf_n146));
   NAND2_X2 U_rbuf_U201 (.ZN(U_rbuf_n128), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[1]));
   OAI21_X2 U_rbuf_U200 (.ZN(hrdata[1]), 
	.B2(U_rbuf_n19), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n128));
   NAND2_X2 U_rbuf_U199 (.ZN(U_rbuf_n136), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[9]));
   OAI21_X2 U_rbuf_U198 (.ZN(hrdata[9]), 
	.B2(U_rbuf_n27), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n136));
   NAND2_X2 U_rbuf_U197 (.ZN(U_rbuf_n130), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[3]));
   OAI21_X2 U_rbuf_U196 (.ZN(hrdata[3]), 
	.B2(U_rbuf_n21), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n130));
   NAND2_X2 U_rbuf_U195 (.ZN(U_rbuf_n132), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[5]));
   OAI21_X2 U_rbuf_U194 (.ZN(hrdata[5]), 
	.B2(U_rbuf_n23), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n132));
   NAND2_X2 U_rbuf_U193 (.ZN(U_rbuf_n134), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[7]));
   OAI21_X2 U_rbuf_U192 (.ZN(hrdata[7]), 
	.B2(U_rbuf_n25), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n134));
   NAND2_X2 U_rbuf_U191 (.ZN(U_rbuf_n160), 
	.A2(big_endian), 
	.A1(m_double));
   NAND2_X2 U_rbuf_U188 (.ZN(U_rbuf_n39), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[29]));
   NAND2_X2 U_rbuf_U187 (.ZN(U_rbuf_n139), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[12]));
   OAI21_X2 U_rbuf_U186 (.ZN(hrdata[12]), 
	.B2(U_rbuf_n30), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n139));
   NAND2_X2 U_rbuf_U185 (.ZN(U_rbuf_n135), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[8]));
   OAI21_X2 U_rbuf_U184 (.ZN(hrdata[8]), 
	.B2(U_rbuf_n26), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n135));
   NAND2_X2 U_rbuf_U183 (.ZN(U_rbuf_n133), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[6]));
   OAI21_X2 U_rbuf_U182 (.ZN(hrdata[6]), 
	.B2(U_rbuf_n24), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n133));
   NAND2_X2 U_rbuf_U181 (.ZN(U_rbuf_n138), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[11]));
   OAI21_X2 U_rbuf_U180 (.ZN(hrdata[11]), 
	.B2(U_rbuf_n29), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n138));
   NAND2_X2 U_rbuf_U179 (.ZN(U_rbuf_n142), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[15]));
   NAND2_X2 U_rbuf_U178 (.ZN(U_rbuf_n131), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[4]));
   OAI21_X2 U_rbuf_U177 (.ZN(hrdata[4]), 
	.B2(U_rbuf_n22), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n131));
   NAND2_X2 U_rbuf_U176 (.ZN(U_rbuf_n129), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[2]));
   OAI21_X2 U_rbuf_U175 (.ZN(hrdata[2]), 
	.B2(U_rbuf_n20), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n129));
   NAND2_X2 U_rbuf_U174 (.ZN(U_rbuf_n127), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[0]));
   OAI21_X2 U_rbuf_U173 (.ZN(hrdata[0]), 
	.B2(U_rbuf_n18), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n127));
   NAND2_X2 U_rbuf_U172 (.ZN(U_rbuf_n140), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[13]));
   NAND2_X2 U_rbuf_U171 (.ZN(U_rbuf_n141), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[14]));
   OAI21_X2 U_rbuf_U170 (.ZN(hrdata[14]), 
	.B2(U_rbuf_n33), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n141));
   NAND2_X2 U_rbuf_U169 (.ZN(U_rbuf_n45), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[25]));
   NAND2_X2 U_rbuf_U168 (.ZN(U_rbuf_n44), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[9]));
   NAND3_X2 U_rbuf_U167 (.ZN(hrdata[25]), 
	.A3(U_rbuf_n43), 
	.A2(U_rbuf_n44), 
	.A1(U_rbuf_n45));
   NAND2_X2 U_rbuf_U166 (.ZN(U_rbuf_n54), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[17]));
   NAND2_X2 U_rbuf_U165 (.ZN(U_rbuf_n53), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[1]));
   NAND3_X2 U_rbuf_U164 (.ZN(hrdata[17]), 
	.A3(U_rbuf_n52), 
	.A2(U_rbuf_n53), 
	.A1(U_rbuf_n54));
   NAND2_X2 U_rbuf_U163 (.ZN(U_rbuf_n51), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[19]));
   NAND2_X2 U_rbuf_U162 (.ZN(U_rbuf_n50), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[3]));
   NAND3_X2 U_rbuf_U161 (.ZN(hrdata[19]), 
	.A3(U_rbuf_n49), 
	.A2(U_rbuf_n50), 
	.A1(U_rbuf_n51));
   NAND2_X2 U_rbuf_U160 (.ZN(U_rbuf_n48), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[21]));
   NAND2_X2 U_rbuf_U159 (.ZN(U_rbuf_n47), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[5]));
   NAND3_X2 U_rbuf_U158 (.ZN(hrdata[21]), 
	.A3(U_rbuf_n46), 
	.A2(U_rbuf_n47), 
	.A1(U_rbuf_n48));
   NAND2_X2 U_rbuf_U157 (.ZN(U_rbuf_n42), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[23]));
   NAND2_X2 U_rbuf_U156 (.ZN(U_rbuf_n41), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[7]));
   NAND3_X2 U_rbuf_U155 (.ZN(hrdata[23]), 
	.A3(U_rbuf_n40), 
	.A2(U_rbuf_n41), 
	.A1(U_rbuf_n42));
   NAND2_X2 U_rbuf_U154 (.ZN(U_rbuf_n137), 
	.A2(U_rbuf_n143), 
	.A1(miu_data[10]));
   NOR2_X2 U_rbuf_U153 (.ZN(U_rbuf_n149), 
	.A2(U_rbuf_f_rbuf_state_1_), 
	.A1(U_rbuf_n154));
   NAND2_X2 U_rbuf_U152 (.ZN(m_rb_ready), 
	.A2(U_rbuf_f_rbuf_state_0_), 
	.A1(U_rbuf_n149));
   NAND2_X2 U_rbuf_U151 (.ZN(U_rbuf_n116), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[16]));
   NAND2_X2 U_rbuf_U150 (.ZN(U_rbuf_n114), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[0]));
   NAND3_X2 U_rbuf_U149 (.ZN(hrdata[16]), 
	.A3(U_rbuf_n114), 
	.A2(U_rbuf_n115), 
	.A1(U_rbuf_n116));
   NAND2_X2 U_rbuf_U148 (.ZN(U_rbuf_n113), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[18]));
   NAND2_X2 U_rbuf_U147 (.ZN(U_rbuf_n111), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[2]));
   NAND3_X2 U_rbuf_U146 (.ZN(hrdata[18]), 
	.A3(U_rbuf_n111), 
	.A2(U_rbuf_n112), 
	.A1(U_rbuf_n113));
   NAND2_X2 U_rbuf_U145 (.ZN(U_rbuf_n101), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[27]));
   NAND2_X2 U_rbuf_U144 (.ZN(U_rbuf_n99), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[11]));
   NAND3_X2 U_rbuf_U143 (.ZN(hrdata[27]), 
	.A3(U_rbuf_n99), 
	.A2(U_rbuf_n100), 
	.A1(U_rbuf_n101));
   NAND2_X2 U_rbuf_U142 (.ZN(U_rbuf_n98), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[28]));
   NAND2_X2 U_rbuf_U141 (.ZN(U_rbuf_n96), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[12]));
   NAND3_X2 U_rbuf_U140 (.ZN(hrdata[28]), 
	.A3(U_rbuf_n96), 
	.A2(U_rbuf_n97), 
	.A1(U_rbuf_n98));
   NAND2_X2 U_rbuf_U139 (.ZN(U_rbuf_n104), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[24]));
   NAND2_X2 U_rbuf_U138 (.ZN(U_rbuf_n102), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[8]));
   NAND3_X2 U_rbuf_U137 (.ZN(hrdata[24]), 
	.A3(U_rbuf_n102), 
	.A2(U_rbuf_n103), 
	.A1(U_rbuf_n104));
   NAND2_X2 U_rbuf_U136 (.ZN(U_rbuf_n92), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[31]));
   NAND2_X2 U_rbuf_U135 (.ZN(U_rbuf_n90), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[15]));
   NAND3_X2 U_rbuf_U134 (.ZN(hrdata[31]), 
	.A3(U_rbuf_n90), 
	.A2(U_rbuf_n91), 
	.A1(U_rbuf_n92));
   NAND2_X2 U_rbuf_U133 (.ZN(U_rbuf_n110), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[20]));
   NAND2_X2 U_rbuf_U132 (.ZN(U_rbuf_n108), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[4]));
   NAND3_X2 U_rbuf_U131 (.ZN(hrdata[20]), 
	.A3(U_rbuf_n108), 
	.A2(U_rbuf_n109), 
	.A1(U_rbuf_n110));
   NAND2_X2 U_rbuf_U130 (.ZN(U_rbuf_n95), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[30]));
   NAND2_X2 U_rbuf_U129 (.ZN(U_rbuf_n93), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[14]));
   NAND3_X2 U_rbuf_U128 (.ZN(hrdata[30]), 
	.A3(U_rbuf_n93), 
	.A2(U_rbuf_n94), 
	.A1(U_rbuf_n95));
   NAND2_X2 U_rbuf_U127 (.ZN(U_rbuf_n107), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[22]));
   NAND2_X2 U_rbuf_U126 (.ZN(U_rbuf_n105), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[6]));
   NAND3_X2 U_rbuf_U125 (.ZN(hrdata[22]), 
	.A3(U_rbuf_n105), 
	.A2(U_rbuf_n106), 
	.A1(U_rbuf_n107));
   AOI21_X2 U_rbuf_U123 (.ZN(U_rbuf_n158), 
	.B2(U_rbuf_f_rbuf_state_0_), 
	.B1(U_rbuf_n157), 
	.A(U_rbuf_n156));
   INV_X4 U_rbuf_U122 (.ZN(U_rbuf_n159), 
	.A(m_rb_start));
   OAI211_X2 U_rbuf_U121 (.ZN(U_rbuf_n88), 
	.C2(U_rbuf_n158), 
	.C1(1'b1), 
	.B(m_rb_ready), 
	.A(U_rbuf_n159));
   NAND2_X1 U_rbuf_U119 (.ZN(U_rbuf_n123), 
	.A2(m_two_to_one), 
	.A1(m_double));
   OAI21_X2 U_rbuf_U117 (.ZN(U_rbuf_n55), 
	.B2(U_rbuf_n180), 
	.B1(U_rbuf_n181), 
	.A(U_rbuf_n162));
   OAI21_X2 U_rbuf_U116 (.ZN(U_rbuf_n66), 
	.B2(U_rbuf_n192), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n173));
   AOI22_X2 U_rbuf_U114 (.ZN(U_rbuf_n169), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_7_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[23]));
   OAI21_X2 U_rbuf_U113 (.ZN(U_rbuf_n62), 
	.B2(FE_PHN4635_U_rbuf_n188), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n169));
   OAI21_X2 U_rbuf_U111 (.ZN(U_rbuf_n65), 
	.B2(U_rbuf_n191), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n172));
   AOI22_X2 U_rbuf_U109 (.ZN(U_rbuf_n165), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_3_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[19]));
   OAI21_X2 U_rbuf_U108 (.ZN(U_rbuf_n58), 
	.B2(U_rbuf_n184), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n165));
   OAI21_X2 U_rbuf_U107 (.ZN(U_rbuf_n69), 
	.B2(U_rbuf_n195), 
	.B1(FE_OFN244_U_rbuf_n180), 
	.A(U_rbuf_n176));
   AOI22_X2 U_rbuf_U106 (.ZN(U_rbuf_n175), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_13_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[29]));
   OAI21_X2 U_rbuf_U105 (.ZN(U_rbuf_n68), 
	.B2(U_rbuf_n194), 
	.B1(U_rbuf_n180), 
	.A(FE_PHN4663_U_rbuf_n175));
   OAI21_X2 U_rbuf_U104 (.ZN(U_rbuf_n63), 
	.B2(U_rbuf_n189), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n170));
   OAI21_X2 U_rbuf_U102 (.ZN(U_rbuf_n64), 
	.B2(U_rbuf_n190), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n171));
   AOI22_X2 U_rbuf_U101 (.ZN(U_rbuf_n179), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_15_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[31]));
   OAI21_X2 U_rbuf_U100 (.ZN(U_rbuf_n70), 
	.B2(U_rbuf_n197), 
	.B1(U_rbuf_n180), 
	.A(FE_PHN4646_U_rbuf_n179));
   OAI21_X2 U_rbuf_U99 (.ZN(U_rbuf_n59), 
	.B2(U_rbuf_n185), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n166));
   AOI22_X2 U_rbuf_U98 (.ZN(U_rbuf_n164), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_2_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[18]));
   OAI21_X2 U_rbuf_U97 (.ZN(U_rbuf_n57), 
	.B2(U_rbuf_n183), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n164));
   AOI22_X2 U_rbuf_U95 (.ZN(U_rbuf_n163), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_1_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[17]));
   OAI21_X2 U_rbuf_U94 (.ZN(U_rbuf_n56), 
	.B2(FE_PHN4644_U_rbuf_n182), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n163));
   OAI21_X2 U_rbuf_U92 (.ZN(U_rbuf_n60), 
	.B2(U_rbuf_n186), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n167));
   AOI22_X2 U_rbuf_U90 (.ZN(U_rbuf_n174), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_12_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[28]));
   OAI21_X2 U_rbuf_U89 (.ZN(U_rbuf_n67), 
	.B2(U_rbuf_n193), 
	.B1(U_rbuf_n180), 
	.A(FE_PHN4647_U_rbuf_n174));
   AOI22_X2 U_rbuf_U87 (.ZN(U_rbuf_n168), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_6_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[22]));
   OAI21_X2 U_rbuf_U86 (.ZN(U_rbuf_n61), 
	.B2(U_rbuf_n187), 
	.B1(U_rbuf_n180), 
	.A(U_rbuf_n168));
   NOR2_X2 U_rbuf_U85 (.ZN(U_rbuf_n124), 
	.A2(U_rbuf_n34), 
	.A1(U_rbuf_n123));
   AOI22_X2 U_rbuf_U84 (.ZN(U_rbuf_n83), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n30), 
	.A2(U_rbuf_n193), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U83 (.ZN(U_rbuf_n84), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n31), 
	.A2(U_rbuf_n194), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U82 (.ZN(U_rbuf_n81), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n28), 
	.A2(U_rbuf_n191), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U81 (.ZN(U_rbuf_n85), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n33), 
	.A2(U_rbuf_n195), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U80 (.ZN(U_rbuf_n71), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n18), 
	.A2(U_rbuf_n181), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U79 (.ZN(U_rbuf_n86), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n32), 
	.A2(U_rbuf_n197), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U78 (.ZN(U_rbuf_n74), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n21), 
	.A2(U_rbuf_n184), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U77 (.ZN(U_rbuf_n79), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n26), 
	.A2(U_rbuf_n189), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U76 (.ZN(U_rbuf_n73), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n20), 
	.A2(U_rbuf_n183), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U75 (.ZN(U_rbuf_n80), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n27), 
	.A2(U_rbuf_n190), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U74 (.ZN(U_rbuf_n72), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n19), 
	.A2(FE_PHN4644_U_rbuf_n182), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U73 (.ZN(U_rbuf_n78), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n25), 
	.A2(FE_PHN4635_U_rbuf_n188), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U72 (.ZN(U_rbuf_n77), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n24), 
	.A2(U_rbuf_n187), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U71 (.ZN(U_rbuf_n75), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n22), 
	.A2(U_rbuf_n185), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U70 (.ZN(U_rbuf_n76), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n23), 
	.A2(U_rbuf_n186), 
	.A1(U_rbuf_n198));
   AOI22_X2 U_rbuf_U69 (.ZN(U_rbuf_n82), 
	.B2(U_rbuf_n196), 
	.B1(U_rbuf_n29), 
	.A2(U_rbuf_n192), 
	.A1(U_rbuf_n198));
   INV_X4 U_rbuf_U68 (.ZN(U_rbuf_n120), 
	.A(big_endian));
   NOR2_X2 U_rbuf_U67 (.ZN(U_rbuf_n198), 
	.A2(U_rbuf_n124), 
	.A1(miu_push_n));
   NAND2_X1 U_rbuf_U66 (.ZN(U_rbuf_n40), 
	.A2(U_rbuf_f_top_data_7_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U65 (.ZN(U_rbuf_n46), 
	.A2(U_rbuf_f_top_data_5_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U64 (.ZN(U_rbuf_n49), 
	.A2(U_rbuf_f_top_data_3_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U63 (.ZN(U_rbuf_n52), 
	.A2(U_rbuf_f_top_data_1_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U62 (.ZN(U_rbuf_n43), 
	.A2(U_rbuf_f_top_data_9_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U61 (.ZN(U_rbuf_n106), 
	.A2(U_rbuf_f_top_data_6_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U60 (.ZN(U_rbuf_n94), 
	.A2(U_rbuf_f_top_data_14_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U59 (.ZN(U_rbuf_n109), 
	.A2(U_rbuf_f_top_data_4_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U58 (.ZN(U_rbuf_n91), 
	.A2(U_rbuf_f_top_data_15_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U57 (.ZN(U_rbuf_n103), 
	.A2(U_rbuf_f_top_data_8_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U56 (.ZN(U_rbuf_n97), 
	.A2(U_rbuf_f_top_data_12_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U55 (.ZN(U_rbuf_n100), 
	.A2(U_rbuf_f_top_data_11_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U54 (.ZN(U_rbuf_n112), 
	.A2(U_rbuf_f_top_data_2_), 
	.A1(U_rbuf_n145));
   NAND2_X1 U_rbuf_U53 (.ZN(U_rbuf_n115), 
	.A2(U_rbuf_f_top_data_0_), 
	.A1(U_rbuf_n145));
   NAND2_X2 U_rbuf_U52 (.ZN(hrdata[15]), 
	.A2(U_rbuf_n142), 
	.A1(U_rbuf_n15));
   NAND3_X2 U_rbuf_U51 (.ZN(hrdata[26]), 
	.A3(U_rbuf_n7), 
	.A2(U_rbuf_n8), 
	.A1(U_rbuf_n9));
   NAND2_X2 U_rbuf_U50 (.ZN(U_rbuf_n7), 
	.A2(U_rbuf_f_top_data_10_), 
	.A1(U_rbuf_n145));
   NAND2_X2 U_rbuf_U49 (.ZN(U_rbuf_n8), 
	.A2(U_rbuf_n16), 
	.A1(miu_data[10]));
   NAND2_X2 U_rbuf_U48 (.ZN(U_rbuf_n9), 
	.A2(U_rbuf_n6), 
	.A1(miu_data[26]));
   NAND2_X2 U_rbuf_U47 (.ZN(U_rbuf_n180), 
	.A2(U_rbuf_n161), 
	.A1(m_two_to_one));
   NOR2_X2 U_rbuf_U46 (.ZN(U_rbuf_n178), 
	.A2(m_two_to_one), 
	.A1(miu_push_n));
   XOR2_X1 U_rbuf_U44 (.Z(U_rbuf_n34), 
	.B(big_endian), 
	.A(U_rbuf_f_1st_half));
   INV_X1 U_rbuf_U40 (.ZN(U_rbuf_n183), 
	.A(miu_data[2]));
   INV_X1 U_rbuf_U39 (.ZN(U_rbuf_n192), 
	.A(miu_data[11]));
   INV_X1 U_rbuf_U38 (.ZN(U_rbuf_n195), 
	.A(miu_data[14]));
   INV_X1 U_rbuf_U37 (.ZN(U_rbuf_n197), 
	.A(miu_data[15]));
   OAI21_X1 U_rbuf_U36 (.ZN(U_rbuf_n157), 
	.B2(m_rb_pop_n), 
	.B1(1'b0), 
	.A(U_rbuf_n154));
   INV_X1 U_rbuf_U35 (.ZN(U_rbuf_n189), 
	.A(miu_data[8]));
   INV_X1 U_rbuf_U34 (.ZN(U_rbuf_n185), 
	.A(miu_data[4]));
   INV_X1 U_rbuf_U33 (.ZN(U_rbuf_n194), 
	.A(miu_data[13]));
   OR2_X2 U_rbuf_U31 (.ZN(U_rbuf_n15), 
	.A2(U_rbuf_n32), 
	.A1(U_rbuf_n143));
   NOR3_X1 U_rbuf_U30 (.ZN(U_rbuf_n156), 
	.A3(U_rbuf_n35), 
	.A2(FE_PHN736_m_rb_overflow), 
	.A1(1'b0));
   INV_X4 U_rbuf_U28 (.ZN(U_rbuf_n6), 
	.A(U_rbuf_n146));
   OAI21_X2 U_rbuf_U27 (.ZN(hrdata[10]), 
	.B2(U_rbuf_n28), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n137));
   AOI22_X1 U_rbuf_U25 (.ZN(U_rbuf_n176), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_14_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[30]));
   AOI22_X1 U_rbuf_U24 (.ZN(U_rbuf_n173), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_11_), 
	.A2(U_rbuf_n178), 
	.A1(FE_PHN4664_miu_data_27_));
   AOI22_X1 U_rbuf_U23 (.ZN(U_rbuf_n172), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_10_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[26]));
   AOI22_X1 U_rbuf_U22 (.ZN(U_rbuf_n171), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_9_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[25]));
   AOI22_X1 U_rbuf_U21 (.ZN(U_rbuf_n170), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_8_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[24]));
   AOI22_X1 U_rbuf_U20 (.ZN(U_rbuf_n167), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_5_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[21]));
   AOI22_X1 U_rbuf_U19 (.ZN(U_rbuf_n166), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_4_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[20]));
   AOI22_X1 U_rbuf_U18 (.ZN(U_rbuf_n162), 
	.B2(U_rbuf_n177), 
	.B1(U_rbuf_f_top_data_0_), 
	.A2(U_rbuf_n178), 
	.A1(miu_data[16]));
   OAI211_X1 U_rbuf_U17 (.ZN(U_rbuf_n89), 
	.C2(U_rbuf_n17), 
	.C1(U_rbuf_n3), 
	.B(U_rbuf_n4), 
	.A(U_rbuf_n159));
   NAND2_X1 U_rbuf_U16 (.ZN(U_rbuf_n4), 
	.A2(U_rbuf_n17), 
	.A1(U_rbuf_n3));
   NOR2_X1 U_rbuf_U15 (.ZN(U_rbuf_n3), 
	.A2(U_ctl_n96), 
	.A1(miu_push_n));
   OR2_X1 U_rbuf_U13 (.ZN(U_rbuf_n146), 
	.A2(m_rb_sel_buf), 
	.A1(m_two_to_one));
   OAI21_X2 U_rbuf_U12 (.ZN(U_rbuf_n145), 
	.B2(U_ctl_n96), 
	.B1(U_rbuf_n160), 
	.A(n48));
   AOI21_X2 U_rbuf_U10 (.ZN(U_rbuf_n38), 
	.B2(U_rbuf_n16), 
	.B1(miu_data[13]), 
	.A(n50));
   NAND2_X2 U_rbuf_U9 (.ZN(hrdata[29]), 
	.A2(U_rbuf_n39), 
	.A1(U_rbuf_n38));
   OAI21_X2 U_rbuf_U8 (.ZN(hrdata[13]), 
	.B2(U_rbuf_n31), 
	.B1(U_rbuf_n143), 
	.A(U_rbuf_n140));
   DFFR_X2 U_rbuf_f_top_data_reg_0_ (.RN(FE_OFN30_HRESETn), 
	.Q(U_rbuf_f_top_data_0_), 
	.D(FE_PHN827_U_rbuf_n55), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_top_data_reg_1_ (.RN(FE_OFN54_HRESETn), 
	.Q(U_rbuf_f_top_data_1_), 
	.D(FE_PHN1069_U_rbuf_n56), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_top_data_reg_2_ (.RN(FE_OFN30_HRESETn), 
	.Q(U_rbuf_f_top_data_2_), 
	.D(FE_PHN1067_U_rbuf_n57), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_top_data_reg_3_ (.RN(FE_OFN30_HRESETn), 
	.Q(U_rbuf_f_top_data_3_), 
	.D(FE_PHN1065_U_rbuf_n58), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_top_data_reg_4_ (.RN(FE_OFN54_HRESETn), 
	.Q(U_rbuf_f_top_data_4_), 
	.D(FE_PHN1073_U_rbuf_n59), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_top_data_reg_5_ (.RN(FE_OFN51_HRESETn), 
	.Q(U_rbuf_f_top_data_5_), 
	.D(FE_PHN1070_U_rbuf_n60), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_top_data_reg_6_ (.RN(FE_OFN160_HRESETn), 
	.Q(U_rbuf_f_top_data_6_), 
	.D(FE_PHN1068_U_rbuf_n61), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_top_data_reg_7_ (.RN(FE_OFN51_HRESETn), 
	.Q(U_rbuf_f_top_data_7_), 
	.D(FE_PHN947_U_rbuf_n62), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_top_data_reg_8_ (.RN(FE_OFN54_HRESETn), 
	.Q(U_rbuf_f_top_data_8_), 
	.D(FE_PHN1075_U_rbuf_n63), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_top_data_reg_9_ (.RN(FE_OFN54_HRESETn), 
	.Q(U_rbuf_f_top_data_9_), 
	.D(FE_PHN1074_U_rbuf_n64), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_top_data_reg_10_ (.RN(FE_OFN51_HRESETn), 
	.Q(U_rbuf_f_top_data_10_), 
	.D(FE_PHN1072_U_rbuf_n65), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_top_data_reg_11_ (.RN(FE_OFN54_HRESETn), 
	.Q(U_rbuf_f_top_data_11_), 
	.D(FE_PHN872_U_rbuf_n66), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_top_data_reg_12_ (.RN(FE_OFN54_HRESETn), 
	.Q(U_rbuf_f_top_data_12_), 
	.D(FE_PHN1071_U_rbuf_n67), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_top_data_reg_13_ (.RN(FE_OFN54_HRESETn), 
	.Q(U_rbuf_f_top_data_13_), 
	.D(FE_PHN876_U_rbuf_n68), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_top_data_reg_14_ (.RN(FE_OFN54_HRESETn), 
	.Q(U_rbuf_f_top_data_14_), 
	.D(FE_PHN828_U_rbuf_n69), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_top_data_reg_15_ (.RN(FE_OFN30_HRESETn), 
	.Q(U_rbuf_f_top_data_15_), 
	.D(FE_PHN1066_U_rbuf_n70), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_btm_data_reg_0_ (.RN(FE_OFN30_HRESETn), 
	.QN(U_rbuf_n18), 
	.D(FE_PHN1676_U_rbuf_n71), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_btm_data_reg_1_ (.RN(FE_OFN54_HRESETn), 
	.QN(U_rbuf_n19), 
	.D(FE_PHN1109_U_rbuf_n72), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_btm_data_reg_2_ (.RN(FE_OFN28_HRESETn), 
	.QN(U_rbuf_n20), 
	.D(FE_PHN1039_U_rbuf_n73), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_btm_data_reg_3_ (.RN(FE_OFN30_HRESETn), 
	.QN(U_rbuf_n21), 
	.D(FE_PHN1105_U_rbuf_n74), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_btm_data_reg_4_ (.RN(FE_OFN28_HRESETn), 
	.QN(U_rbuf_n22), 
	.D(FE_PHN1112_U_rbuf_n75), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_btm_data_reg_5_ (.RN(FE_OFN30_HRESETn), 
	.QN(U_rbuf_n23), 
	.D(FE_PHN930_U_rbuf_n76), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_btm_data_reg_6_ (.RN(FE_OFN54_HRESETn), 
	.QN(U_rbuf_n24), 
	.D(FE_PHN1108_U_rbuf_n77), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_btm_data_reg_7_ (.RN(FE_OFN30_HRESETn), 
	.QN(U_rbuf_n25), 
	.D(FE_PHN1104_U_rbuf_n78), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_btm_data_reg_8_ (.RN(FE_OFN54_HRESETn), 
	.QN(U_rbuf_n26), 
	.D(FE_PHN1114_U_rbuf_n79), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_btm_data_reg_9_ (.RN(FE_OFN54_HRESETn), 
	.QN(U_rbuf_n27), 
	.D(FE_PHN1110_U_rbuf_n80), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_btm_data_reg_10_ (.RN(FE_OFN30_HRESETn), 
	.QN(U_rbuf_n28), 
	.D(FE_PHN929_U_rbuf_n81), 
	.CK(hclk));
   DFFR_X2 U_rbuf_f_btm_data_reg_11_ (.RN(FE_OFN54_HRESETn), 
	.QN(U_rbuf_n29), 
	.D(FE_PHN1679_U_rbuf_n82), 
	.CK(HCLK__L5_N5));
   DFFR_X2 U_rbuf_f_btm_data_reg_12_ (.RN(FE_OFN54_HRESETn), 
	.QN(U_rbuf_n30), 
	.D(FE_PHN1111_U_rbuf_n83), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_rbuf_f_btm_data_reg_13_ (.RN(FE_OFN54_HRESETn), 
	.QN(U_rbuf_n31), 
	.D(FE_PHN1678_U_rbuf_n84), 
	.CK(HCLK__L5_N5));
   DFFR_X2 U_rbuf_f_btm_data_reg_14_ (.RN(FE_OFN54_HRESETn), 
	.QN(U_rbuf_n33), 
	.D(FE_PHN1677_U_rbuf_n85), 
	.CK(HCLK__L5_N5));
   DFFR_X2 U_rbuf_f_btm_data_reg_15_ (.RN(FE_OFN30_HRESETn), 
	.QN(U_rbuf_n32), 
	.D(FE_PHN1115_U_rbuf_n86), 
	.CK(hclk));
   DFFR_X1 U_rbuf_f_rbuf_state_reg_1_ (.RN(FE_OFN153_HRESETn), 
	.QN(U_rbuf_n35), 
	.Q(U_rbuf_f_rbuf_state_1_), 
	.D(1'b0), 
	.CK(hclk));
   DFFR_X1 U_rbuf_f_rbuf_state_reg_0_ (.RN(FE_OFN153_HRESETn), 
	.Q(U_rbuf_f_rbuf_state_0_), 
	.D(FE_PHN1231_U_rbuf_n88), 
	.CK(hclk));
   DFFS_X2 U_rbuf_f_1st_half_reg (.SN(FE_OFN30_HRESETn), 
	.QN(U_rbuf_n17), 
	.Q(U_rbuf_f_1st_half), 
	.D(FE_PHN2930_U_rbuf_n89), 
	.CK(hclk));
   OAI21_X1 U_ctl_U457 (.ZN(U_ctl_n347), 
	.B2(U_ctl_n349), 
	.B1(U_rbuf_n120), 
	.A(m_two_to_one));
   NOR2_X1 U_ctl_U456 (.ZN(U_ctl_N89), 
	.A2(FE_PHN3141_U_ctl_n421), 
	.A1(htrans[1]));
   INV_X4 U_ctl_U455 (.ZN(U_ctl_n326), 
	.A(FE_PHN2913_U_ctl_n422));
   INV_X4 U_ctl_U452 (.ZN(U_ctl_n276), 
	.A(haddr[5]));
   NAND2_X2 U_ctl_U451 (.ZN(U_ctl_n418), 
	.A2(big_endian), 
	.A1(U_ctl_fd_wr_width));
   AND3_X4 U_ctl_U448 (.ZN(U_ctl_n318), 
	.A3(haddr[5]), 
	.A2(1'b1), 
	.A1(1'b1));
   MUX2_X2 U_ctl_U447 (.Z(m_df_data_in[25]), 
	.S(U_ctl_n364), 
	.B(hwdata[23]), 
	.A(hwdata[7]));
   MUX2_X2 U_ctl_U446 (.Z(m_df_data_in[18]), 
	.S(U_ctl_n364), 
	.B(hwdata[16]), 
	.A(hwdata[0]));
   MUX2_X2 U_ctl_U444 (.Z(m_df_data_in[33]), 
	.S(U_ctl_n364), 
	.B(hwdata[31]), 
	.A(hwdata[15]));
   MUX2_X2 U_ctl_U443 (.Z(m_df_data_in[26]), 
	.S(U_ctl_n364), 
	.B(hwdata[24]), 
	.A(hwdata[8]));
   NOR2_X2 U_ctl_U440 (.ZN(U_ctl_n248), 
	.A2(U_ctl_n346), 
	.A1(U_ctl_n63));
   NOR2_X2 U_ctl_U437 (.ZN(U_ctl_n325), 
	.A2(haddr[7]), 
	.A1(haddr[6]));
   NAND2_X2 U_ctl_U436 (.ZN(U_ctl_n201), 
	.A2(U_ctl_fd_miu_col_width_2_), 
	.A1(U_ctl_fd_miu_col_width_0_));
   NOR2_X2 U_ctl_U435 (.ZN(U_ctl_n202), 
	.A2(U_ctl_fd_miu_data_width_0_), 
	.A1(U_ctl_fd_miu_data_width_1_));
   INV_X4 U_ctl_U433 (.ZN(U_ctl_n288), 
	.A(haddr[2]));
   INV_X4 U_ctl_U432 (.ZN(U_ctl_n289), 
	.A(haddr[3]));
   NAND2_X2 U_ctl_U431 (.ZN(U_ctl_n269), 
	.A2(U_ctl_n289), 
	.A1(U_ctl_n288));
   NAND2_X2 U_ctl_U430 (.ZN(U_ctl_n329), 
	.A2(U_ctl_n276), 
	.A1(U_ctl_n267));
   INV_X4 U_ctl_U429 (.ZN(U_ctl_n227), 
	.A(hsize[0]));
   NAND2_X2 U_ctl_U428 (.ZN(U_ctl_n199), 
	.A2(hsize[1]), 
	.A1(U_ctl_n227));
   NAND2_X2 U_ctl_U427 (.ZN(U_ctl_n208), 
	.A2(1'b1), 
	.A1(U_ctl_n248));
   NOR2_X2 U_ctl_U426 (.ZN(U_ctl_n193), 
	.A2(haddr[4]), 
	.A1(haddr[7]));
   NAND3_X2 U_ctl_U425 (.ZN(U_ctl_n198), 
	.A3(U_ctl_n276), 
	.A2(U_ctl_n288), 
	.A1(U_ctl_n193));
   OAI211_X2 U_ctl_U424 (.ZN(U_ctl_n195), 
	.C2(U_ctl_n154), 
	.C1(U_ctl_fd_miu_col_width_1_), 
	.B(U_ctl_n194), 
	.A(U_ctl_n202));
   NOR2_X2 U_ctl_U423 (.ZN(U_ctl_n196), 
	.A2(U_ctl_n195), 
	.A1(haddr[3]));
   NAND2_X2 U_ctl_U422 (.ZN(U_ctl_n197), 
	.A2(U_ctl_n235), 
	.A1(U_ctl_n196));
   NOR2_X2 U_ctl_U421 (.ZN(U_ctl_n200), 
	.A2(U_ctl_n197), 
	.A1(U_ctl_n198));
   NAND2_X2 U_ctl_U420 (.ZN(U_ctl_n167), 
	.A2(U_ctl_n201), 
	.A1(U_ctl_n166));
   NOR2_X2 U_ctl_U418 (.ZN(U_ctl_n305), 
	.A2(U_ctl_f_bh_state_2_), 
	.A1(U_ctl_f_bh_state_1_));
   NAND2_X2 U_ctl_U417 (.ZN(U_ctl_n221), 
	.A2(U_ctl_n158), 
	.A1(U_ctl_n98));
   AOI21_X2 U_ctl_U416 (.ZN(U_ctl_n211), 
	.B2(U_ctl_n209), 
	.B1(miu_push_n), 
	.A(U_ctl_n221));
   NOR3_X2 U_ctl_U415 (.ZN(U_ctl_n336), 
	.A3(U_ctl_fd_amba_bcnt_2_), 
	.A2(U_ctl_fd_amba_bcnt_1_), 
	.A1(U_ctl_fd_amba_bcnt_0_));
   NOR2_X2 U_ctl_U414 (.ZN(U_ctl_n210), 
	.A2(U_ctl_fd_incr), 
	.A1(U_ctl_fd_amba_bcnt_3_));
   NAND2_X2 U_ctl_U413 (.ZN(U_ctl_n220), 
	.A2(U_ctl_n210), 
	.A1(U_ctl_n336));
   NAND3_X2 U_ctl_U412 (.ZN(U_ctl_n212), 
	.A3(U_ctl_n220), 
	.A2(U_ctl_n211), 
	.A1(hready));
   NAND2_X2 U_ctl_U411 (.ZN(m_rb_pop_n), 
	.A2(U_ctl_fd_rd_ready), 
	.A1(hready));
   NOR2_X2 U_ctl_U410 (.ZN(U_ctl_n341), 
	.A2(m_af_new_req), 
	.A1(U_ctl_fr_prv_1wrap_tm));
   NOR2_X2 U_ctl_U409 (.ZN(U_ctl_n214), 
	.A2(U_ctl_n186), 
	.A1(FE_PHN736_m_rb_overflow));
   NOR3_X2 U_ctl_U408 (.ZN(U_ctl_n308), 
	.A3(U_ctl_fr_wr_bcnt_3_), 
	.A2(U_ctl_fr_wr_bcnt_1_), 
	.A1(U_ctl_n339));
   INV_X4 U_ctl_U407 (.ZN(U_ctl_n292), 
	.A(U_ctl_n304));
   OAI211_X2 U_ctl_U406 (.ZN(U_ctl_n297), 
	.C2(U_ctl_f_bh_state_0_), 
	.C1(U_ctl_n214), 
	.B(U_ctl_n292), 
	.A(U_ctl_n305));
   INV_X4 U_ctl_U401 (.ZN(U_ctl_n403), 
	.A(hwdata[14]));
   INV_X4 U_ctl_U400 (.ZN(U_ctl_n402), 
	.A(hwdata[22]));
   NOR2_X2 U_ctl_U399 (.ZN(U_ctl_n168), 
	.A2(U_rbuf_n120), 
	.A1(U_ctl_n402));
   NOR2_X2 U_ctl_U398 (.ZN(U_ctl_n170), 
	.A2(U_ctl_n168), 
	.A1(U_ctl_n169));
   NOR2_X2 U_ctl_U397 (.ZN(U_ctl_n400), 
	.A2(U_ctl_n126), 
	.A1(U_ctl_n170));
   NOR2_X2 U_ctl_U396 (.ZN(U_ctl_n335), 
	.A2(big_endian), 
	.A1(U_ctl_n126));
   INV_X4 U_ctl_U395 (.ZN(U_ctl_n183), 
	.A(FE_PHN888_U_ctl_n150));
   NOR2_X2 U_ctl_U388 (.ZN(U_ctl_n251), 
	.A2(U_ctl_n346), 
	.A1(U_ctl_n398));
   NAND2_X2 U_ctl_U387 (.ZN(U_ctl_n252), 
	.A2(U_ctl_n250), 
	.A1(U_ctl_n251));
   NAND2_X2 U_ctl_U386 (.ZN(U_ctl_n180), 
	.A2(U_ctl_n252), 
	.A1(FE_PHN888_U_ctl_n150));
   NOR2_X2 U_ctl_U377 (.ZN(m_af_data2_in[7]), 
	.A2(U_ctl_n173), 
	.A1(U_ctl_n89));
   NAND2_X2 U_ctl_U376 (.ZN(U_ctl_n382), 
	.A2(hready), 
	.A1(U_ctl_n251));
   INV_X4 U_ctl_U375 (.ZN(U_ctl_n337), 
	.A(FE_PHN699_U_ctl_n382));
   OAI21_X2 U_ctl_U374 (.ZN(U_ctl_n392), 
	.B2(1'b1), 
	.B1(U_ctl_n336), 
	.A(U_ctl_n337));
   AOI22_X2 U_ctl_U373 (.ZN(U_ctl_n394), 
	.B2(U_ctl_n392), 
	.B1(U_ctl_fd_amba_bcnt_3_), 
	.A2(1'b0), 
	.A1(1'b0));
   OAI21_X2 U_ctl_U372 (.ZN(U_ctl_n116), 
	.B2(1'b1), 
	.B1(U_ctl_fd_amba_bcnt_3_), 
	.A(FE_PHN1506_U_ctl_n394));
   NAND3_X2 U_ctl_U371 (.ZN(U_ctl_n364), 
	.A3(m_two_to_one), 
	.A2(big_endian), 
	.A1(U_ctl_n98));
   NOR3_X2 U_ctl_U357 (.ZN(U_ctl_n323), 
	.A3(1'b0), 
	.A2(1'b0), 
	.A1(FE_PHN699_U_ctl_n382));
   OAI21_X2 U_ctl_U355 (.ZN(U_ctl_n395), 
	.B2(U_ctl_n143), 
	.B1(1'b1), 
	.A(U_ctl_n337));
   NAND2_X2 U_ctl_U340 (.ZN(U_ctl_n349), 
	.A2(U_ctl_fd_haddr_1_), 
	.A1(U_ctl_fd_narrow_trans));
   AOI21_X2 U_ctl_U339 (.ZN(U_ctl_n375), 
	.B2(U_ctl_n349), 
	.B1(U_rbuf_n120), 
	.A(U_ctl_n347));
   AOI21_X2 U_ctl_U338 (.ZN(U_ctl_n348), 
	.B2(U_ctl_n349), 
	.B1(U_rbuf_n120), 
	.A(U_ctl_n96));
   OAI21_X2 U_ctl_U337 (.ZN(U_ctl_n374), 
	.B2(U_ctl_n349), 
	.B1(U_rbuf_n120), 
	.A(U_ctl_n348));
   AOI22_X2 U_ctl_U336 (.ZN(U_ctl_n350), 
	.B2(hwdata[8]), 
	.B1(U_ctl_n374), 
	.A2(hwdata[24]), 
	.A1(U_ctl_n375));
   INV_X4 U_ctl_U335 (.ZN(m_df_data_in[10]), 
	.A(U_ctl_n350));
   AOI22_X2 U_ctl_U334 (.ZN(U_ctl_n351), 
	.B2(hwdata[15]), 
	.B1(U_ctl_n374), 
	.A2(hwdata[31]), 
	.A1(U_ctl_n375));
   INV_X4 U_ctl_U333 (.ZN(m_df_data_in[17]), 
	.A(U_ctl_n351));
   NAND3_X2 U_ctl_U332 (.ZN(U_ctl_n294), 
	.A3(m_rb_ready), 
	.A2(m_af_ready), 
	.A1(m_df_ready));
   NAND2_X2 U_ctl_U331 (.ZN(hready_resp), 
	.A2(U_ctl_n151), 
	.A1(U_ctl_n294));
   AOI22_X2 U_ctl_U330 (.ZN(U_ctl_n376), 
	.B2(hwdata[7]), 
	.B1(U_ctl_n374), 
	.A2(hwdata[23]), 
	.A1(U_ctl_n375));
   INV_X4 U_ctl_U329 (.ZN(m_df_data_in[9]), 
	.A(U_ctl_n376));
   NAND4_X2 U_ctl_U328 (.ZN(FE_PHN676_hiu_terminate), 
	.A4(U_ctl_n293), 
	.A3(U_ctl_n306), 
	.A2(FE_PHN700_U_ctl_n297), 
	.A1(FE_PHN682_U_ctl_n295));
   NAND2_X2 U_ctl_U325 (.ZN(m_af_data1_in_5_), 
	.A2(U_ctl_n174), 
	.A1(1'b1));
   AOI22_X2 U_ctl_U321 (.ZN(U_ctl_n358), 
	.B2(hwdata[0]), 
	.B1(U_ctl_n374), 
	.A2(hwdata[16]), 
	.A1(U_ctl_n375));
   INV_X4 U_ctl_U320 (.ZN(m_df_data_in[2]), 
	.A(U_ctl_n358));
   INV_X4 U_ctl_U319 (.ZN(U_ctl_n363), 
	.A(U_ctl_n364));
   AOI22_X2 U_ctl_U318 (.ZN(m_df_data_in[24]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n402), 
	.A2(U_ctl_n371), 
	.A1(U_ctl_n363));
   INV_X4 U_ctl_U317 (.ZN(U_ctl_n373), 
	.A(U_ctl_n375));
   INV_X4 U_ctl_U316 (.ZN(U_ctl_n372), 
	.A(U_ctl_n374));
   OAI22_X2 U_ctl_U315 (.ZN(m_df_data_in[14]), 
	.B2(U_ctl_n360), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n359), 
	.A1(U_ctl_n373));
   OAI22_X2 U_ctl_U314 (.ZN(m_df_data_in[11]), 
	.B2(U_ctl_n353), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n352), 
	.A1(U_ctl_n373));
   OAI22_X2 U_ctl_U313 (.ZN(m_df_data_in[13]), 
	.B2(U_ctl_n357), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n356), 
	.A1(U_ctl_n373));
   OAI22_X2 U_ctl_U312 (.ZN(m_df_data_in[12]), 
	.B2(U_ctl_n355), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n354), 
	.A1(U_ctl_n373));
   OAI22_X2 U_ctl_U311 (.ZN(U_ctl_n119), 
	.B2(U_ctl_n143), 
	.B1(U_ctl_n337), 
	.A2(U_ctl_n395), 
	.A1(U_ctl_n323));
   AOI22_X2 U_ctl_U310 (.ZN(m_df_data_in[23]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n370), 
	.A2(U_ctl_n369), 
	.A1(U_ctl_n363));
   OAI22_X2 U_ctl_U309 (.ZN(m_df_data_in[16]), 
	.B2(U_ctl_n362), 
	.B1(U_ctl_n373), 
	.A2(U_ctl_n372), 
	.A1(U_ctl_n403));
   INV_X4 U_ctl_U308 (.ZN(U_ctl_n361), 
	.A(hwdata[29]));
   OAI22_X2 U_ctl_U307 (.ZN(m_df_data_in[15]), 
	.B2(U_ctl_n372), 
	.B1(U_ctl_n222), 
	.A2(U_ctl_n373), 
	.A1(U_ctl_n361));
   INV_X4 U_ctl_U306 (.ZN(U_ctl_n414), 
	.A(hwdata[18]));
   AOI22_X2 U_ctl_U305 (.ZN(m_df_data_in[20]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n414), 
	.A2(U_ctl_n366), 
	.A1(U_ctl_n363));
   INV_X4 U_ctl_U304 (.ZN(U_ctl_n417), 
	.A(hwdata[17]));
   AOI22_X2 U_ctl_U303 (.ZN(m_df_data_in[19]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n417), 
	.A2(U_ctl_n365), 
	.A1(U_ctl_n363));
   INV_X4 U_ctl_U302 (.ZN(U_ctl_n408), 
	.A(hwdata[20]));
   AOI22_X2 U_ctl_U301 (.ZN(m_df_data_in[22]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n408), 
	.A2(U_ctl_n368), 
	.A1(U_ctl_n363));
   INV_X4 U_ctl_U300 (.ZN(U_ctl_n411), 
	.A(hwdata[19]));
   AOI22_X2 U_ctl_U299 (.ZN(m_df_data_in[21]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n411), 
	.A2(U_ctl_n367), 
	.A1(U_ctl_n363));
   AOI22_X2 U_ctl_U298 (.ZN(U_ctl_n391), 
	.B2(U_ctl_fd_rd_ready), 
	.B1(FE_PHN3141_U_ctl_n421), 
	.A2(U_ctl_n337), 
	.A1(m_af_data1_in_2_));
   INV_X4 U_ctl_U297 (.ZN(U_ctl_n106), 
	.A(U_ctl_n391));
   OAI22_X2 U_ctl_U296 (.ZN(m_df_data_in[8]), 
	.B2(U_ctl_n371), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n373), 
	.A1(U_ctl_n402));
   OAI22_X2 U_ctl_U293 (.ZN(m_df_data_in[5]), 
	.B2(U_ctl_n367), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n411), 
	.A1(U_ctl_n373));
   OAI22_X2 U_ctl_U292 (.ZN(m_df_data_in[4]), 
	.B2(U_ctl_n366), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n414), 
	.A1(U_ctl_n373));
   OAI22_X2 U_ctl_U291 (.ZN(m_df_data_in[7]), 
	.B2(U_ctl_n369), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n373), 
	.A1(U_ctl_n370));
   OAI22_X2 U_ctl_U290 (.ZN(m_df_data_in[6]), 
	.B2(U_ctl_n368), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n408), 
	.A1(U_ctl_n373));
   OAI22_X2 U_ctl_U289 (.ZN(m_df_data_in[3]), 
	.B2(U_ctl_n365), 
	.B1(U_ctl_n372), 
	.A2(U_ctl_n417), 
	.A1(U_ctl_n373));
   OAI22_X2 U_ctl_U287 (.ZN(U_ctl_n401), 
	.B2(U_ctl_n326), 
	.B1(U_ctl_fd_miu_data_width_1_), 
	.A2(FE_PHN1079_U_ctl_n400), 
	.A1(FE_PHN2913_U_ctl_n422));
   INV_X4 U_ctl_U286 (.ZN(U_ctl_n125), 
	.A(U_ctl_n401));
   NOR3_X2 U_ctl_U285 (.ZN(m_af_data1_in_11_), 
	.A3(U_ctl_n378), 
	.A2(U_ctl_n183), 
	.A1(FE_PHN1079_U_ctl_n400));
   AOI22_X2 U_ctl_U284 (.ZN(U_ctl_n124), 
	.B2(U_ctl_n324), 
	.B1(FE_PHN2913_U_ctl_n422), 
	.A2(U_ctl_n326), 
	.A1(FE_PHN795_U_ctl_n180));
   AOI22_X2 U_ctl_U283 (.ZN(m_df_data_in[31]), 
	.B2(U_ctl_n363), 
	.B1(U_ctl_n222), 
	.A2(U_ctl_n364), 
	.A1(U_ctl_n361));
   AOI22_X2 U_ctl_U282 (.ZN(U_ctl_n410), 
	.B2(U_ctl_n126), 
	.B1(U_ctl_f_col_width[2]), 
	.A2(FE_PHN747_U_ctl_n335), 
	.A1(hwdata[11]));
   OAI21_X2 U_ctl_U281 (.ZN(U_ctl_n133), 
	.B2(U_ctl_n411), 
	.B1(FE_PHN708_U_ctl_n418), 
	.A(U_ctl_n410));
   OAI22_X2 U_ctl_U280 (.ZN(U_ctl_n412), 
	.B2(U_ctl_n326), 
	.B1(U_ctl_fd_miu_col_width_2_), 
	.A2(FE_PHN1106_U_ctl_n133), 
	.A1(FE_PHN2913_U_ctl_n422));
   INV_X4 U_ctl_U279 (.ZN(U_ctl_n129), 
	.A(U_ctl_n412));
   AOI22_X2 U_ctl_U278 (.ZN(m_df_data_in[32]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n362), 
	.A2(U_ctl_n403), 
	.A1(U_ctl_n363));
   AOI22_X2 U_ctl_U277 (.ZN(U_ctl_n413), 
	.B2(U_ctl_n126), 
	.B1(U_ctl_f_col_width[1]), 
	.A2(FE_PHN747_U_ctl_n335), 
	.A1(hwdata[10]));
   OAI21_X2 U_ctl_U276 (.ZN(U_ctl_n134), 
	.B2(U_ctl_n414), 
	.B1(FE_PHN708_U_ctl_n418), 
	.A(U_ctl_n413));
   OAI22_X2 U_ctl_U275 (.ZN(U_ctl_n415), 
	.B2(U_ctl_n326), 
	.B1(U_ctl_fd_miu_col_width_1_), 
	.A2(FE_PHN1107_U_ctl_n134), 
	.A1(FE_PHN2913_U_ctl_n422));
   INV_X4 U_ctl_U274 (.ZN(U_ctl_n130), 
	.A(U_ctl_n415));
   AOI22_X2 U_ctl_U273 (.ZN(U_ctl_n407), 
	.B2(U_ctl_n126), 
	.B1(U_ctl_f_col_width[3]), 
	.A2(FE_PHN747_U_ctl_n335), 
	.A1(hwdata[12]));
   OAI21_X2 U_ctl_U272 (.ZN(U_ctl_n132), 
	.B2(U_ctl_n408), 
	.B1(FE_PHN708_U_ctl_n418), 
	.A(U_ctl_n407));
   OAI22_X2 U_ctl_U271 (.ZN(U_ctl_n409), 
	.B2(U_ctl_n326), 
	.B1(U_ctl_fd_miu_col_width_3_), 
	.A2(FE_PHN975_U_ctl_n132), 
	.A1(FE_PHN2913_U_ctl_n422));
   INV_X4 U_ctl_U270 (.ZN(U_ctl_n128), 
	.A(U_ctl_n409));
   AOI22_X2 U_ctl_U269 (.ZN(U_ctl_n416), 
	.B2(U_ctl_n126), 
	.B1(U_ctl_f_col_width[0]), 
	.A2(FE_PHN747_U_ctl_n335), 
	.A1(hwdata[9]));
   OAI21_X2 U_ctl_U268 (.ZN(U_ctl_n135), 
	.B2(U_ctl_n417), 
	.B1(FE_PHN708_U_ctl_n418), 
	.A(U_ctl_n416));
   OAI22_X2 U_ctl_U267 (.ZN(U_ctl_n419), 
	.B2(U_ctl_n326), 
	.B1(U_ctl_fd_miu_col_width_0_), 
	.A2(FE_PHN1011_U_ctl_n135), 
	.A1(FE_PHN2913_U_ctl_n422));
   INV_X4 U_ctl_U266 (.ZN(U_ctl_n131), 
	.A(U_ctl_n419));
   NAND4_X2 U_ctl_U264 (.ZN(U_ctl_n327), 
	.A4(U_ctl_n326), 
	.A3(1'b1), 
	.A2(U_ctl_n380), 
	.A1(FE_OFN210_hwrite_s));
   NAND2_X2 U_ctl_U263 (.ZN(U_ctl_n405), 
	.A2(U_ctl_f_data_width_0_), 
	.A1(U_ctl_n171));
   OAI211_X2 U_ctl_U262 (.ZN(U_ctl_n127), 
	.C2(U_ctl_n406), 
	.C1(FE_PHN708_U_ctl_n418), 
	.B(U_ctl_n404), 
	.A(U_ctl_n405));
   AOI22_X2 U_ctl_U261 (.ZN(m_df_data_in[28]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n354), 
	.A2(U_ctl_n355), 
	.A1(U_ctl_n363));
   AOI22_X2 U_ctl_U260 (.ZN(m_df_data_in[27]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n352), 
	.A2(U_ctl_n353), 
	.A1(U_ctl_n363));
   AOI22_X2 U_ctl_U259 (.ZN(m_df_data_in[29]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n356), 
	.A2(U_ctl_n357), 
	.A1(U_ctl_n363));
   AOI22_X2 U_ctl_U258 (.ZN(m_df_data_in[30]), 
	.B2(U_ctl_n364), 
	.B1(U_ctl_n359), 
	.A2(U_ctl_n360), 
	.A1(U_ctl_n363));
   NOR2_X2 U_ctl_U257 (.ZN(U_ctl_N236), 
	.A2(U_ctl_n342), 
	.A1(m_af_dummy_req));
   AOI22_X2 U_ctl_U256 (.ZN(U_ctl_n122), 
	.B2(U_ctl_n96), 
	.B1(FE_PHN2913_U_ctl_n422), 
	.A2(U_ctl_n326), 
	.A1(U_ctl_n183));
   AOI22_X2 U_ctl_U255 (.ZN(U_ctl_n123), 
	.B2(FE_PHN2913_U_ctl_n422), 
	.B1(U_ctl_n147), 
	.A2(U_ctl_n326), 
	.A1(FE_PHN888_U_ctl_n150));
   OAI22_X2 U_ctl_U254 (.ZN(U_ctl_n120), 
	.B2(U_ctl_n146), 
	.B1(U_ctl_n326), 
	.A2(1'b1), 
	.A1(hwrite));
   NOR4_X2 U_ctl_U253 (.ZN(U_ctl_n309), 
	.A4(U_ctl_n310), 
	.A3(hiu_burst_size[1]), 
	.A2(hiu_burst_size[5]), 
	.A1(U_ctl_n340));
   AOI211_X2 U_ctl_U252 (.ZN(U_ctl_n313), 
	.C2(U_ctl_n384), 
	.C1(U_ctl_n309), 
	.B(U_ctl_n386), 
	.A(FE_PHN1036_U_ctl_f_hiu_terminate));
   NAND2_X2 U_ctl_U251 (.ZN(U_ctl_n312), 
	.A2(U_ctl_n313), 
	.A1(U_ctl_C64_DATA2_5));
   NOR3_X2 U_ctl_U250 (.ZN(U_ctl_n389), 
	.A3(U_ctl_n384), 
	.A2(U_ctl_n385), 
	.A1(FE_PHN1036_U_ctl_f_hiu_terminate));
   NOR3_X2 U_ctl_U249 (.ZN(U_ctl_n388), 
	.A3(U_ctl_n386), 
	.A2(U_ctl_n144), 
	.A1(U_ctl_fr_prv_1wrap));
   AOI22_X2 U_ctl_U248 (.ZN(U_ctl_n387), 
	.B2(hiu_burst_size[5]), 
	.B1(U_ctl_n388), 
	.A2(U_ctl_n389), 
	.A1(U_ctl_fr_wr_bcnt_5_));
   NAND3_X2 U_ctl_U247 (.ZN(U_ctl_n100), 
	.A3(U_ctl_n311), 
	.A2(U_ctl_n387), 
	.A1(U_ctl_n312));
   OAI22_X2 U_ctl_U246 (.ZN(U_ctl_n420), 
	.B2(U_ctl_n326), 
	.B1(U_ctl_fd_haddr_1_), 
	.A2(haddr[1]), 
	.A1(FE_PHN2913_U_ctl_n422));
   INV_X4 U_ctl_U245 (.ZN(U_ctl_n137), 
	.A(U_ctl_n420));
   AOI211_X2 U_ctl_U242 (.ZN(U_ctl_n296), 
	.C2(U_ctl_n345), 
	.C1(1'b0), 
	.B(1'b0), 
	.A(U_ctl_n301));
   NOR2_X2 U_ctl_U241 (.ZN(U_ctl_n_sel_buf), 
	.A2(U_ctl_n296), 
	.A1(U_ctl_n307));
   AOI22_X2 U_ctl_U240 (.ZN(U_ctl_n141), 
	.B2(FE_PHN2913_U_ctl_n422), 
	.B1(U_ctl_n156), 
	.A2(U_ctl_n326), 
	.A1(1'b1));
   AOI22_X2 U_ctl_U239 (.ZN(U_ctl_n390), 
	.B2(FE_OFN220_hiu_burst_size_0_), 
	.B1(U_ctl_n388), 
	.A2(U_ctl_n389), 
	.A1(FE_PHN999_U_ctl_fr_wr_bcnt_0_));
   NAND3_X2 U_ctl_U238 (.ZN(U_ctl_n105), 
	.A3(U_ctl_n315), 
	.A2(U_ctl_n390), 
	.A1(U_ctl_n316));
   INV_X1 U_ctl_U235 (.ZN(U_ctl_n384), 
	.A(miu_pop_n));
   NOR2_X1 U_ctl_U234 (.ZN(U_ctl_n385), 
	.A2(m_af_new_req), 
	.A1(hiu_rw));
   NAND2_X2 U_ctl_U233 (.ZN(U_ctl_n422), 
	.A2(hready), 
	.A1(1'b1));
   NOR2_X2 U_ctl_U232 (.ZN(U_ctl_DP_OP_140_125_8947_I2), 
	.A2(miu_pop_n), 
	.A1(U_ctl_n309));
   OAI22_X2 U_ctl_U230 (.ZN(U_ctl_n139), 
	.B2(U_ctl_n98), 
	.B1(U_ctl_n326), 
	.A2(U_ctl_n331), 
	.A1(FE_PHN699_U_ctl_n382));
   NAND2_X1 U_ctl_U228 (.ZN(U_ctl_n380), 
	.A2(hsize[0]), 
	.A1(hsize[1]));
   AOI221_X1 U_ctl_U227 (.ZN(U_ctl_n379), 
	.C2(U_ctl_n378), 
	.C1(haddr[0]), 
	.B2(U_ctl_n378), 
	.B1(hsize[0]), 
	.A(hsize[1]));
   INV_X1 U_ctl_U226 (.ZN(U_ctl_n230), 
	.A(hsize[1]));
   NAND3_X2 U_ctl_U224 (.ZN(U_ctl_n187), 
	.A3(U_ctl_n331), 
	.A2(1'b1), 
	.A1(U_ctl_n47));
   AOI22_X1 U_ctl_U223 (.ZN(U_ctl_n140), 
	.B2(U_ctl_n160), 
	.B1(FE_PHN2913_U_ctl_n422), 
	.A2(U_ctl_n383), 
	.A1(1'b1));
   AOI21_X2 U_ctl_U222 (.ZN(U_ctl_n290), 
	.B2(1'b0), 
	.B1(U_ctl_n187), 
	.A(FE_PHN2923_U_ctl_n212));
   NOR2_X1 U_ctl_U217 (.ZN(U_ctl_n398), 
	.A2(hsel_mem), 
	.A1(FE_PHN2917_hsel_reg));
   NAND2_X1 U_ctl_U215 (.ZN(U_ctl_n317), 
	.A2(haddr[4]), 
	.A1(1'b1));
   INV_X4 U_ctl_U207 (.ZN(U_ctl_n63), 
	.A(hsel_mem));
   NAND2_X2 U_ctl_U204 (.ZN(U_ctl_n174), 
	.A2(U_ctl_n50), 
	.A1(1'b1));
   OAI22_X2 U_ctl_U203 (.ZN(U_ctl_n136), 
	.B2(U_ctl_n126), 
	.B1(U_ctl_n326), 
	.A2(m_af_data1_in_0_), 
	.A1(U_ctl_n330));
   OAI22_X2 U_ctl_U202 (.ZN(U_ctl_n138), 
	.B2(U_ctl_n158), 
	.B1(U_ctl_n326), 
	.A2(FE_PHN3141_U_ctl_n421), 
	.A1(m_af_data1_in_0_));
   NAND3_X2 U_ctl_U200 (.ZN(U_ctl_n85), 
	.A3(U_ctl_n208), 
	.A2(1'b1), 
	.A1(m_af_data1_in_0_));
   INV_X2 U_ctl_U197 (.ZN(U_ctl_n235), 
	.A(haddr[6]));
   INV_X2 U_ctl_U196 (.ZN(U_ctl_n346), 
	.A(htrans[1]));
   INV_X2 U_ctl_U195 (.ZN(U_ctl_n378), 
	.A(haddr[1]));
   INV_X2 U_ctl_U194 (.ZN(U_ctl_n366), 
	.A(hwdata[2]));
   INV_X2 U_ctl_U193 (.ZN(m_af_data1_in_2_), 
	.A(hwrite));
   INV_X2 U_ctl_U192 (.ZN(U_ctl_n365), 
	.A(hwdata[1]));
   INV_X2 U_ctl_U191 (.ZN(U_ctl_n371), 
	.A(hwdata[6]));
   INV_X2 U_ctl_U190 (.ZN(U_ctl_n355), 
	.A(hwdata[10]));
   INV_X2 U_ctl_U189 (.ZN(U_ctl_n359), 
	.A(hwdata[28]));
   INV_X2 U_ctl_U188 (.ZN(U_ctl_n368), 
	.A(hwdata[4]));
   INV_X2 U_ctl_U187 (.ZN(U_ctl_n360), 
	.A(hwdata[12]));
   NAND2_X2 U_ctl_U186 (.ZN(m_af_data1_in_0_), 
	.A2(htrans[1]), 
	.A1(FE_PHN5181_hsel_reg));
   INV_X2 U_ctl_U185 (.ZN(U_ctl_n354), 
	.A(hwdata[26]));
   INV_X2 U_ctl_U184 (.ZN(U_ctl_n367), 
	.A(hwdata[3]));
   INV_X2 U_ctl_U183 (.ZN(U_ctl_n357), 
	.A(hwdata[11]));
   INV_X2 U_ctl_U182 (.ZN(U_ctl_n356), 
	.A(hwdata[27]));
   INV_X2 U_ctl_U181 (.ZN(U_ctl_n352), 
	.A(hwdata[25]));
   INV_X2 U_ctl_U180 (.ZN(U_ctl_n353), 
	.A(hwdata[9]));
   INV_X2 U_ctl_U179 (.ZN(U_ctl_n362), 
	.A(hwdata[30]));
   INV_X2 U_ctl_U178 (.ZN(U_ctl_n369), 
	.A(hwdata[5]));
   INV_X2 U_ctl_U177 (.ZN(U_ctl_n370), 
	.A(hwdata[21]));
   INV_X2 U_ctl_U176 (.ZN(U_ctl_n222), 
	.A(hwdata[13]));
   NAND2_X1 U_ctl_U175 (.ZN(U_ctl_n406), 
	.A2(U_ctl_n402), 
	.A1(hwdata[21]));
   INV_X1 U_ctl_U173 (.ZN(U_ctl_n328), 
	.A(U_ctl_n325));
   OR3_X2 U_ctl_U172 (.ZN(U_ctl_n339), 
	.A3(U_ctl_fr_wr_bcnt_5_), 
	.A2(U_ctl_fr_wr_bcnt_4_), 
	.A1(U_ctl_fr_wr_bcnt_2_));
   NAND3_X1 U_ctl_U171 (.ZN(U_ctl_n343), 
	.A3(U_ctl_n142), 
	.A2(U_ctl_f_bh_state_1_), 
	.A1(U_ctl_f_bh_state_0_));
   NOR2_X2 U_ctl_U170 (.ZN(U_ctl_n55), 
	.A2(U_ctl_f_data_width_0_), 
	.A1(U_ctl_fd_wr_width));
   OR3_X2 U_ctl_U169 (.ZN(U_ctl_n293), 
	.A3(U_ctl_f_burst_done2), 
	.A2(FE_PHN2904_U_ctl_f_burst_done), 
	.A1(U_ctl_n144));
   INV_X1 U_ctl_U164 (.ZN(U_ctl_n421), 
	.A(hready));
   NOR2_X1 U_ctl_U161 (.ZN(U_ctl_n169), 
	.A2(big_endian), 
	.A1(U_ctl_n403));
   NOR2_X2 U_ctl_U158 (.ZN(U_ctl_n267), 
	.A2(haddr[4]), 
	.A1(U_ctl_n269));
   INV_X2 U_ctl_U156 (.ZN(U_ctl_n345), 
	.A(U_ctl_n343));
   NOR2_X1 U_ctl_U151 (.ZN(U_ctl_n383), 
	.A2(FE_PHN2913_U_ctl_n422), 
	.A1(1'b0));
   NAND3_X1 U_ctl_U150 (.ZN(U_ctl_n404), 
	.A3(U_ctl_n403), 
	.A2(FE_PHN747_U_ctl_n335), 
	.A1(hwdata[13]));
   INV_X2 U_ctl_U149 (.ZN(U_ctl_n54), 
	.A(FE_PHN747_U_ctl_n335));
   INV_X1 U_ctl_U148 (.ZN(U_ctl_n87), 
	.A(U_ctl_n317));
   NOR2_X2 U_ctl_U146 (.ZN(U_ctl_n331), 
	.A2(1'b0), 
	.A1(U_ctl_n199));
   NOR2_X2 U_ctl_U145 (.ZN(U_ctl_n56), 
	.A2(U_ctl_n54), 
	.A1(hwdata[13]));
   OR4_X2 U_ctl_U143 (.ZN(U_ctl_n330), 
	.A4(U_ctl_n327), 
	.A3(U_ctl_n328), 
	.A2(U_ctl_n329), 
	.A1(U_ctl_n379));
   INV_X2 U_ctl_U142 (.ZN(U_ctl_n250), 
	.A(U_ctl_n331));
   NAND2_X1 U_ctl_U141 (.ZN(U_ctl_n171), 
	.A2(U_ctl_fd_wr_width), 
	.A1(U_ctl_n170));
   NOR2_X2 U_ctl_U140 (.ZN(U_ctl_n58), 
	.A2(U_ctl_n55), 
	.A1(U_ctl_n56));
   OR4_X2 U_ctl_U139 (.ZN(U_ctl_n340), 
	.A4(hiu_burst_size[3]), 
	.A3(FE_OFN217_hiu_burst_size_2_), 
	.A2(FE_OFN214_hiu_burst_size_4_), 
	.A1(FE_OFN220_hiu_burst_size_0_));
   INV_X2 U_ctl_U138 (.ZN(U_ctl_n386), 
	.A(U_ctl_n385));
   NAND2_X2 U_ctl_U137 (.ZN(U_ctl_n150), 
	.A2(U_ctl_n57), 
	.A1(U_ctl_n58));
   INV_X4 U_ctl_U136 (.ZN(U_ctl_n50), 
	.A(FE_PHN795_U_ctl_n180));
   NAND2_X1 U_ctl_U135 (.ZN(U_ctl_n299), 
	.A2(U_ctl_n337), 
	.A1(hwrite));
   INV_X2 U_ctl_U133 (.ZN(U_ctl_n342), 
	.A(hiu_wrap_burst));
   NAND2_X1 U_ctl_U130 (.ZN(U_ctl_n311), 
	.A2(U_ctl_N288), 
	.A1(U_ctl_n314));
   NAND2_X1 U_ctl_U128 (.ZN(U_ctl_n315), 
	.A2(U_ctl_n97), 
	.A1(U_ctl_n314));
   AOI21_X2 U_ctl_U119 (.ZN(U_ctl_n295), 
	.B2(U_ctl_n290), 
	.B1(1'b1), 
	.A(m_df_wr_term));
   NAND2_X1 U_ctl_U116 (.ZN(U_ctl_n316), 
	.A2(U_ctl_n313), 
	.A1(U_ctl_C64_DATA2_0));
   INV_X2 U_ctl_U115 (.ZN(U_ctl_n307), 
	.A(FE_PHN682_U_ctl_n295));
   AND2_X2 U_ctl_U113 (.ZN(U_ctl_N237), 
	.A2(U_ctl_N236), 
	.A1(hiu_terminate));
   OAI21_X2 U_ctl_U108 (.ZN(U_ctl_n92), 
	.B2(U_ctl_n91), 
	.B1(1'b0), 
	.A(1'b1));
   NOR2_X2 U_ctl_U105 (.ZN(U_ctl_n173), 
	.A2(U_ctl_n92), 
	.A1(FE_PHN888_U_ctl_n150));
   NOR2_X2 U_ctl_U104 (.ZN(U_ctl_n88), 
	.A2(U_ctl_n87), 
	.A1(1'b0));
   NAND2_X2 U_ctl_U103 (.ZN(m_af_push1_n), 
	.A2(hready), 
	.A1(U_ctl_n85));
   NOR2_X2 U_ctl_U101 (.ZN(m_rb_start), 
	.A2(hwrite), 
	.A1(FE_PHN673_m_af_push1_n));
   NOR2_X2 U_ctl_U100 (.ZN(U_ctl_n225), 
	.A2(U_ctl_n88), 
	.A1(1'b0));
   NAND2_X2 U_ctl_U96 (.ZN(U_ctl_n194), 
	.A2(U_ctl_fd_miu_col_width_1_), 
	.A1(U_ctl_fd_miu_col_width_3_));
   NAND3_X1 U_ctl_U93 (.ZN(U_ctl_n209), 
	.A3(U_ctl_f_bh_state_0_), 
	.A2(U_ctl_fd_rd_bz), 
	.A1(U_ctl_n305));
   INV_X1 U_ctl_U91 (.ZN(U_ctl_n91), 
	.A(U_ctl_n318));
   OR2_X2 U_ctl_U89 (.ZN(U_ctl_n57), 
	.A2(FE_PHN708_U_ctl_n418), 
	.A1(hwdata[21]));
   INV_X4 U_ctl_U88 (.ZN(U_ctl_n186), 
	.A(U_ctl_n341));
   NAND2_X1 U_ctl_U87 (.ZN(U_ctl_n310), 
	.A2(U_ctl_n97), 
	.A1(U_ctl_n308));
   INV_X1 U_ctl_U79 (.ZN(U_ctl_n301), 
	.A(U_ctl_n306));
   AND2_X4 U_ctl_U74 (.ZN(U_ctl_n47), 
	.A2(U_ctl_n200), 
	.A1(U_ctl_n167));
   NAND2_X1 U_ctl_U73 (.ZN(U_ctl_n104), 
	.A2(U_ctl_n44), 
	.A1(U_ctl_n45));
   NAND2_X1 U_ctl_U72 (.ZN(U_ctl_n45), 
	.A2(U_ctl_N284), 
	.A1(U_ctl_n314));
   AOI222_X1 U_ctl_U71 (.ZN(U_ctl_n44), 
	.C2(U_ctl_n43), 
	.C1(U_ctl_n313), 
	.B2(U_ctl_n388), 
	.B1(hiu_burst_size[1]), 
	.A2(U_ctl_n389), 
	.A1(U_ctl_fr_wr_bcnt_1_));
   XOR2_X1 U_ctl_U70 (.Z(U_ctl_n43), 
	.B(U_ctl_DP_OP_140_125_8947_n9), 
	.A(U_ctl_DP_OP_140_125_8947_n14));
   NOR2_X1 U_ctl_U69 (.ZN(U_ctl_n_bh_state[0]), 
	.A2(U_ctl_n42), 
	.A1(U_ctl_n307));
   AOI21_X1 U_ctl_U68 (.ZN(U_ctl_n42), 
	.B2(1'b0), 
	.B1(U_ctl_f_bh_state_0_), 
	.A(U_ctl_n41));
   OAI22_X1 U_ctl_U67 (.ZN(U_ctl_n41), 
	.B2(U_ctl_n40), 
	.B1(FE_PHN736_m_rb_overflow), 
	.A2(1'b1), 
	.A1(U_ctl_n306));
   NAND3_X1 U_ctl_U66 (.ZN(U_ctl_n40), 
	.A3(U_ctl_n39), 
	.A2(U_ctl_n304), 
	.A1(U_ctl_n305));
   OAI22_X1 U_ctl_U65 (.ZN(U_ctl_n39), 
	.B2(U_ctl_n38), 
	.B1(miu_burst_done), 
	.A2(U_ctl_n95), 
	.A1(U_ctl_n342));
   NOR2_X1 U_ctl_U64 (.ZN(U_ctl_n38), 
	.A2(U_ctl_n341), 
	.A1(U_ctl_f_bh_state_0_));
   OAI211_X1 U_ctl_U61 (.ZN(U_ctl_n117), 
	.C2(U_ctl_n36), 
	.C1(U_ctl_n148), 
	.B(1'b1), 
	.A(1'b1));
   AOI21_X1 U_ctl_U60 (.ZN(U_ctl_n36), 
	.B2(1'b0), 
	.B1(U_ctl_fd_amba_bcnt_1_), 
	.A(U_ctl_n395));
   AOI21_X1 U_ctl_U59 (.ZN(m_af_data1_in_13_), 
	.B2(FE_PHN1079_U_ctl_n400), 
	.B1(U_ctl_n183), 
	.A(U_ctl_n289));
   XOR2_X1 U_ctl_U58 (.Z(U_ctl_N288), 
	.B(U_ctl_n35), 
	.A(U_ctl_fr_wr_bcnt_5_));
   NOR2_X1 U_ctl_U57 (.ZN(U_ctl_n35), 
	.A2(U_ctl_DP_OP_140_125_8947_n22), 
	.A1(U_ctl_fr_wr_bcnt_4_));
   NAND2_X1 U_ctl_U51 (.ZN(U_ctl_n103), 
	.A2(U_ctl_n30), 
	.A1(U_ctl_n28));
   AOI222_X1 U_ctl_U50 (.ZN(U_ctl_n30), 
	.C2(U_ctl_n29), 
	.C1(U_ctl_n313), 
	.B2(U_ctl_n388), 
	.B1(FE_OFN217_hiu_burst_size_2_), 
	.A2(U_ctl_n389), 
	.A1(U_ctl_fr_wr_bcnt_2_));
   XOR2_X1 U_ctl_U49 (.Z(U_ctl_n29), 
	.B(U_ctl_DP_OP_140_125_8947_n13), 
	.A(U_ctl_DP_OP_140_125_8947_n7));
   NAND2_X1 U_ctl_U48 (.ZN(U_ctl_n28), 
	.A2(U_ctl_N285), 
	.A1(U_ctl_n314));
   AOI221_X1 U_ctl_U47 (.ZN(U_ctl_n_bh_state[1]), 
	.C2(1'b1), 
	.C1(1'b0), 
	.B2(1'b1), 
	.B1(FE_PHN700_U_ctl_n297), 
	.A(U_ctl_n307));
   NAND2_X1 U_ctl_U36 (.ZN(U_ctl_n102), 
	.A2(U_ctl_n21), 
	.A1(U_ctl_n19));
   AOI222_X1 U_ctl_U35 (.ZN(U_ctl_n21), 
	.C2(U_ctl_n20), 
	.C1(U_ctl_n313), 
	.B2(U_ctl_n388), 
	.B1(hiu_burst_size[3]), 
	.A2(U_ctl_n389), 
	.A1(U_ctl_fr_wr_bcnt_3_));
   XOR2_X1 U_ctl_U34 (.Z(U_ctl_n20), 
	.B(U_ctl_DP_OP_140_125_8947_n12), 
	.A(U_ctl_DP_OP_140_125_8947_n5));
   NAND2_X1 U_ctl_U33 (.ZN(U_ctl_n19), 
	.A2(U_ctl_N286), 
	.A1(U_ctl_n314));
   NAND3_X1 U_ctl_U29 (.ZN(U_ctl_n166), 
	.A3(U_ctl_n16), 
	.A2(U_ctl_n99), 
	.A1(U_ctl_fd_miu_col_width_3_));
   INV_X1 U_ctl_U28 (.ZN(U_ctl_n16), 
	.A(haddr[8]));
   NAND2_X1 U_ctl_U27 (.ZN(U_ctl_n101), 
	.A2(U_ctl_n15), 
	.A1(U_ctl_n13));
   AOI222_X1 U_ctl_U26 (.ZN(U_ctl_n15), 
	.C2(U_ctl_n14), 
	.C1(U_ctl_n313), 
	.B2(U_ctl_n388), 
	.B1(FE_OFN214_hiu_burst_size_4_), 
	.A2(U_ctl_n389), 
	.A1(U_ctl_fr_wr_bcnt_4_));
   XOR2_X1 U_ctl_U25 (.Z(U_ctl_n14), 
	.B(U_ctl_DP_OP_140_125_8947_n11), 
	.A(U_ctl_DP_OP_140_125_8947_n3));
   NAND2_X1 U_ctl_U24 (.ZN(U_ctl_n13), 
	.A2(U_ctl_N287), 
	.A1(U_ctl_n314));
   NOR2_X2 U_ctl_U23 (.ZN(m_af_data1_in_4_), 
	.A2(1'b0), 
	.A1(U_ctl_n50));
   NOR2_X1 U_ctl_U22 (.ZN(U_ctl_n89), 
	.A2(U_ctl_n183), 
	.A1(U_ctl_n225));
   NOR2_X1 U_ctl_U20 (.ZN(m_df_data_in[0]), 
	.A2(U_ctl_n221), 
	.A1(U_ctl_n11));
   AOI22_X1 U_ctl_U19 (.ZN(U_ctl_n11), 
	.B2(U_ctl_n220), 
	.B1(1'b1), 
	.A2(U_ctl_fd_non_single), 
	.A1(1'b0));
   NOR2_X1 U_ctl_U13 (.ZN(U_ctl_n314), 
	.A2(U_ctl_n6), 
	.A1(miu_pop_n));
   NAND3_X1 U_ctl_U12 (.ZN(U_ctl_n6), 
	.A3(U_ctl_n310), 
	.A2(U_ctl_n386), 
	.A1(U_ctl_n144));
   NAND3_X1 U_ctl_U8 (.ZN(U_ctl_n306), 
	.A3(U_ctl_n305), 
	.A2(FE_PHN736_m_rb_overflow), 
	.A1(U_ctl_n3));
   NAND2_X1 U_ctl_U7 (.ZN(U_ctl_n3), 
	.A2(U_ctl_f_bh_state_0_), 
	.A1(U_ctl_n292));
   DFFR_X2 U_ctl_f_hiu_terminate_reg (.RN(FE_OFN51_HRESETn), 
	.QN(U_ctl_n144), 
	.Q(U_ctl_f_hiu_terminate), 
	.D(hiu_terminate), 
	.CK(hclk));
   DFFR_X2 U_ctl_fr_wr_bcnt_reg_0_ (.RN(FE_OFN51_HRESETn), 
	.QN(U_ctl_n97), 
	.Q(U_ctl_fr_wr_bcnt_0_), 
	.D(FE_PHN744_U_ctl_n105), 
	.CK(HCLK__L5_N17));
   DFFR_X2 U_ctl_fd_miu_col_width_reg_2_ (.RN(FE_OFN55_HRESETn), 
	.QN(U_ctl_n154), 
	.Q(U_ctl_fd_miu_col_width_2_), 
	.D(FE_PHN1509_U_ctl_n129), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_miu_col_width_reg_0_ (.RN(FE_OFN55_HRESETn), 
	.QN(U_ctl_n99), 
	.Q(U_ctl_fd_miu_col_width_0_), 
	.D(FE_PHN1507_U_ctl_n131), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_miu_col_width_reg_1_ (.RN(FE_OFN55_HRESETn), 
	.QN(), 
	.Q(U_ctl_fd_miu_col_width_1_), 
	.D(FE_PHN1511_U_ctl_n130), 
	.CK(HCLK__L5_N27));
   DFFR_X2 U_ctl_fd_miu_data_width_reg_0_ (.RN(FE_OFN55_HRESETn), 
	.QN(U_ctl_n147), 
	.Q(U_ctl_fd_miu_data_width_0_), 
	.D(FE_PHN885_U_ctl_n123), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_amba_bcnt_reg_2_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_ctl_n148), 
	.Q(U_ctl_fd_amba_bcnt_2_), 
	.D(FE_PHN1681_U_ctl_n117), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_ctl_o_two_to_one_reg (.RN(FE_OFN30_HRESETn), 
	.QN(U_ctl_n96), 
	.Q(m_two_to_one), 
	.D(FE_PHN1370_U_ctl_n122), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_wr_width_reg (.RN(FE_OFN55_HRESETn), 
	.QN(U_ctl_n126), 
	.Q(U_ctl_fd_wr_width), 
	.D(FE_PHN1368_U_ctl_n136), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_amba_bcnt_reg_0_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_ctl_n143), 
	.Q(U_ctl_fd_amba_bcnt_0_), 
	.D(FE_PHN1505_U_ctl_n119), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_ctl_fd_non_single_reg (.RN(FE_OFN153_HRESETn), 
	.QN(U_ctl_n160), 
	.Q(U_ctl_fd_non_single), 
	.D(FE_PHN1609_U_ctl_n140), 
	.CK(HCLK__L5_N27));
   DFFR_X2 U_ctl_fd_narrow_trans_reg (.RN(FE_OFN55_HRESETn), 
	.QN(U_ctl_n98), 
	.Q(U_ctl_fd_narrow_trans), 
	.D(FE_PHN1162_U_ctl_n139), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_rd_bz_reg (.RN(FE_OFN153_HRESETn), 
	.QN(U_ctl_n146), 
	.Q(U_ctl_fd_rd_bz), 
	.D(FE_PHN1684_U_ctl_n120), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_incr_reg (.RN(FE_OFN153_HRESETn), 
	.QN(U_ctl_n156), 
	.Q(U_ctl_fd_incr), 
	.D(FE_PHN1904_U_ctl_n141), 
	.CK(HCLK__L5_N27));
   DFFR_X2 U_ctl_fd_amba_bcnt_reg_3_ (.RN(FE_OFN153_HRESETn), 
	.QN(), 
	.Q(U_ctl_fd_amba_bcnt_3_), 
	.D(U_ctl_n116), 
	.CK(HCLK__L5_N27));
   DFFR_X2 U_ctl_fd_double_reg (.RN(FE_OFN30_HRESETn), 
	.QN(U_ctl_n324), 
	.Q(m_double), 
	.D(FE_PHN1232_U_ctl_n124), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_amba_bcnt_reg_1_ (.RN(FE_OFN153_HRESETn), 
	.QN(U_ctl_n145), 
	.Q(U_ctl_fd_amba_bcnt_1_), 
	.D(FE_PHN3152_U_ctl_n118), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_ctl_fd_miu_col_width_reg_3_ (.RN(FE_OFN55_HRESETn), 
	.Q(U_ctl_fd_miu_col_width_3_), 
	.D(FE_PHN1510_U_ctl_n128), 
	.CK(hclk));
   DFFR_X2 U_ctl_fr_prv_1wrap_reg (.RN(FE_OFN51_HRESETn), 
	.Q(U_ctl_fr_prv_1wrap), 
	.D(U_ctl_N236), 
	.CK(HCLK__L5_N35));
   DFFR_X2 U_ctl_f_col_width_reg_2_ (.RN(FE_OFN55_HRESETn), 
	.Q(U_ctl_f_col_width[2]), 
	.D(FE_PHN1106_U_ctl_n133), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_miu_data_width_reg_1_ (.RN(FE_OFN55_HRESETn), 
	.Q(U_ctl_fd_miu_data_width_1_), 
	.D(FE_PHN1233_U_ctl_n125), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_haddr_reg_1_ (.RN(FE_OFN55_HRESETn), 
	.Q(U_ctl_fd_haddr_1_), 
	.D(FE_PHN1611_U_ctl_n137), 
	.CK(HCLK__L5_N27));
   DFFR_X2 U_ctl_f_burst_done2_reg (.RN(FE_OFN51_HRESETn), 
	.Q(U_ctl_f_burst_done2), 
	.D(FE_PHN2904_U_ctl_f_burst_done), 
	.CK(hclk));
   DFFR_X2 U_ctl_fd_reg_access_reg (.RN(FE_OFN55_HRESETn), 
	.QN(U_ctl_n158), 
	.D(FE_PHN1229_U_ctl_n138), 
	.CK(hclk));
   INV_X2 U_ctl_DP_OP_140_125_8947_U31 (.ZN(U_ctl_DP_OP_140_125_8947_n30), 
	.A(U_ctl_DP_OP_140_125_8947_n20));
   XNOR2_X1 U_ctl_DP_OP_140_125_8947_U38 (.ZN(U_ctl_N285), 
	.B(U_ctl_fr_wr_bcnt_2_), 
	.A(U_ctl_DP_OP_140_125_8947_n24));
   XOR2_X1 U_ctl_DP_OP_140_125_8947_U2 (.Z(U_ctl_DP_OP_140_125_8947_n1), 
	.B(U_ctl_DP_OP_140_125_8947_n35), 
	.A(hiu_burst_size[5]));
   XOR2_X1 U_ctl_DP_OP_140_125_8947_U19 (.Z(U_ctl_C64_DATA2_0), 
	.B(U_ctl_DP_OP_140_125_8947_n30), 
	.A(FE_OFN220_hiu_burst_size_0_));
   INV_X2 U_ctl_DP_OP_140_125_8947_U21 (.ZN(U_ctl_DP_OP_140_125_8947_n35), 
	.A(U_ctl_DP_OP_140_125_8947_n15));
   OR2_X2 U_ctl_DP_OP_140_125_8947_U37 (.ZN(U_ctl_DP_OP_140_125_8947_n22), 
	.A2(U_ctl_fr_wr_bcnt_3_), 
	.A1(U_ctl_DP_OP_140_125_8947_n23));
   XNOR2_X1 U_ctl_DP_OP_140_125_8947_U36 (.ZN(U_ctl_N286), 
	.B(U_ctl_fr_wr_bcnt_3_), 
	.A(U_ctl_DP_OP_140_125_8947_n23));
   OR2_X2 U_ctl_DP_OP_140_125_8947_U39 (.ZN(U_ctl_DP_OP_140_125_8947_n23), 
	.A2(U_ctl_fr_wr_bcnt_2_), 
	.A1(U_ctl_DP_OP_140_125_8947_n24));
   OR2_X2 U_ctl_DP_OP_140_125_8947_U41 (.ZN(U_ctl_DP_OP_140_125_8947_n24), 
	.A2(U_ctl_fr_wr_bcnt_1_), 
	.A1(FE_PHN999_U_ctl_fr_wr_bcnt_0_));
   AOI22_X1 U_ctl_DP_OP_140_125_8947_U24 (.ZN(U_ctl_DP_OP_140_125_8947_n16), 
	.B2(U_ctl_fr_wr_bcnt_4_), 
	.B1(miu_pop_n), 
	.A2(U_ctl_DP_OP_140_125_8947_I2), 
	.A1(U_ctl_N287));
   AOI22_X1 U_ctl_DP_OP_140_125_8947_U26 (.ZN(U_ctl_DP_OP_140_125_8947_n17), 
	.B2(U_ctl_fr_wr_bcnt_3_), 
	.B1(miu_pop_n), 
	.A2(U_ctl_DP_OP_140_125_8947_I2), 
	.A1(U_ctl_N286));
   AOI22_X1 U_ctl_DP_OP_140_125_8947_U28 (.ZN(U_ctl_DP_OP_140_125_8947_n18), 
	.B2(U_ctl_fr_wr_bcnt_2_), 
	.B1(miu_pop_n), 
	.A2(U_ctl_DP_OP_140_125_8947_I2), 
	.A1(U_ctl_N285));
   AOI22_X1 U_ctl_DP_OP_140_125_8947_U32 (.ZN(U_ctl_DP_OP_140_125_8947_n20), 
	.B2(FE_PHN999_U_ctl_fr_wr_bcnt_0_), 
	.B1(miu_pop_n), 
	.A2(U_ctl_DP_OP_140_125_8947_I2), 
	.A1(U_ctl_n97));
   AOI22_X1 U_ctl_DP_OP_140_125_8947_U30 (.ZN(U_ctl_DP_OP_140_125_8947_n19), 
	.B2(U_ctl_fr_wr_bcnt_1_), 
	.B1(miu_pop_n), 
	.A2(U_ctl_DP_OP_140_125_8947_I2), 
	.A1(U_ctl_N284));
   AOI22_X1 U_ctl_DP_OP_140_125_8947_U22 (.ZN(U_ctl_DP_OP_140_125_8947_n15), 
	.B2(U_ctl_fr_wr_bcnt_5_), 
	.B1(miu_pop_n), 
	.A2(U_ctl_DP_OP_140_125_8947_I2), 
	.A1(U_ctl_N288));
   INV_X4 U_ctl_DP_OP_140_125_8947_U4 (.ZN(U_ctl_DP_OP_140_125_8947_n10), 
	.A(U_ctl_DP_OP_140_125_8947_n2));
   AOI22_X2 U_ctl_DP_OP_140_125_8947_U5 (.ZN(U_ctl_DP_OP_140_125_8947_n2), 
	.B2(FE_OFN214_hiu_burst_size_4_), 
	.B1(U_ctl_DP_OP_140_125_8947_n34), 
	.A2(U_ctl_DP_OP_140_125_8947_n3), 
	.A1(U_ctl_DP_OP_140_125_8947_n11));
   INV_X4 U_ctl_DP_OP_140_125_8947_U23 (.ZN(U_ctl_DP_OP_140_125_8947_n34), 
	.A(U_ctl_DP_OP_140_125_8947_n16));
   INV_X4 U_ctl_DP_OP_140_125_8947_U8 (.ZN(U_ctl_DP_OP_140_125_8947_n11), 
	.A(U_ctl_DP_OP_140_125_8947_n4));
   AOI22_X2 U_ctl_DP_OP_140_125_8947_U9 (.ZN(U_ctl_DP_OP_140_125_8947_n4), 
	.B2(hiu_burst_size[3]), 
	.B1(U_ctl_DP_OP_140_125_8947_n33), 
	.A2(U_ctl_DP_OP_140_125_8947_n5), 
	.A1(U_ctl_DP_OP_140_125_8947_n12));
   INV_X4 U_ctl_DP_OP_140_125_8947_U25 (.ZN(U_ctl_DP_OP_140_125_8947_n33), 
	.A(U_ctl_DP_OP_140_125_8947_n17));
   INV_X4 U_ctl_DP_OP_140_125_8947_U12 (.ZN(U_ctl_DP_OP_140_125_8947_n12), 
	.A(U_ctl_DP_OP_140_125_8947_n6));
   AOI22_X2 U_ctl_DP_OP_140_125_8947_U13 (.ZN(U_ctl_DP_OP_140_125_8947_n6), 
	.B2(FE_OFN217_hiu_burst_size_2_), 
	.B1(U_ctl_DP_OP_140_125_8947_n32), 
	.A2(U_ctl_DP_OP_140_125_8947_n7), 
	.A1(U_ctl_DP_OP_140_125_8947_n13));
   INV_X4 U_ctl_DP_OP_140_125_8947_U27 (.ZN(U_ctl_DP_OP_140_125_8947_n32), 
	.A(U_ctl_DP_OP_140_125_8947_n18));
   INV_X4 U_ctl_DP_OP_140_125_8947_U16 (.ZN(U_ctl_DP_OP_140_125_8947_n13), 
	.A(U_ctl_DP_OP_140_125_8947_n8));
   AOI22_X2 U_ctl_DP_OP_140_125_8947_U17 (.ZN(U_ctl_DP_OP_140_125_8947_n8), 
	.B2(hiu_burst_size[1]), 
	.B1(U_ctl_DP_OP_140_125_8947_n31), 
	.A2(U_ctl_DP_OP_140_125_8947_n14), 
	.A1(U_ctl_DP_OP_140_125_8947_n9));
   INV_X4 U_ctl_DP_OP_140_125_8947_U29 (.ZN(U_ctl_DP_OP_140_125_8947_n31), 
	.A(U_ctl_DP_OP_140_125_8947_n19));
   XOR2_X2 U_ctl_DP_OP_140_125_8947_U1 (.Z(U_ctl_C64_DATA2_5), 
	.B(U_ctl_DP_OP_140_125_8947_n10), 
	.A(U_ctl_DP_OP_140_125_8947_n1));
   XOR2_X2 U_ctl_DP_OP_140_125_8947_U6 (.Z(U_ctl_DP_OP_140_125_8947_n3), 
	.B(U_ctl_DP_OP_140_125_8947_n34), 
	.A(FE_OFN214_hiu_burst_size_4_));
   XOR2_X2 U_ctl_DP_OP_140_125_8947_U10 (.Z(U_ctl_DP_OP_140_125_8947_n5), 
	.B(U_ctl_DP_OP_140_125_8947_n33), 
	.A(hiu_burst_size[3]));
   XOR2_X2 U_ctl_DP_OP_140_125_8947_U14 (.Z(U_ctl_DP_OP_140_125_8947_n7), 
	.B(U_ctl_DP_OP_140_125_8947_n32), 
	.A(FE_OFN217_hiu_burst_size_2_));
   XOR2_X2 U_ctl_DP_OP_140_125_8947_U18 (.Z(U_ctl_DP_OP_140_125_8947_n9), 
	.B(U_ctl_DP_OP_140_125_8947_n31), 
	.A(hiu_burst_size[1]));
   AND2_X4 U_ctl_DP_OP_140_125_8947_U20 (.ZN(U_ctl_DP_OP_140_125_8947_n14), 
	.A2(FE_OFN220_hiu_burst_size_0_), 
	.A1(U_ctl_DP_OP_140_125_8947_n30));
   XNOR2_X2 U_ctl_DP_OP_140_125_8947_U34 (.ZN(U_ctl_N287), 
	.B(U_ctl_fr_wr_bcnt_4_), 
	.A(U_ctl_DP_OP_140_125_8947_n22));
   XNOR2_X2 U_ctl_DP_OP_140_125_8947_U40 (.ZN(U_ctl_N284), 
	.B(U_ctl_fr_wr_bcnt_1_), 
	.A(FE_PHN999_U_ctl_fr_wr_bcnt_0_));
   DFFR_X1 U_ctl_f_sel_buf_reg (.RN(FE_OFN30_HRESETn), 
	.QN(n48), 
	.Q(m_rb_sel_buf), 
	.D(FE_PHN4632_U_ctl_n_sel_buf), 
	.CK(hclk));
   DFFR_X1 U_ctl_f_bh_state_reg_1_ (.RN(FE_OFN153_HRESETn), 
	.Q(U_ctl_f_bh_state_1_), 
	.D(U_ctl_n_bh_state[1]), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_ctl_fr_prv_1wrap_tm_reg (.RN(FE_OFN153_HRESETn), 
	.Q(U_ctl_fr_prv_1wrap_tm), 
	.D(U_ctl_N237), 
	.CK(hclk));
   DFFR_X1 U_ctl_f_bh_state_reg_2_ (.RN(FE_OFN153_HRESETn), 
	.QN(U_ctl_n142), 
	.Q(U_ctl_f_bh_state_2_), 
	.D(1'b0), 
	.CK(hclk));
   DFFR_X1 U_ctl_f_bh_state_reg_0_ (.RN(FE_OFN153_HRESETn), 
	.QN(U_ctl_n95), 
	.Q(U_ctl_f_bh_state_0_), 
	.D(FE_PHN4640_U_ctl_n_bh_state_0_), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_ctl_fr_wr_bcnt_reg_5_ (.RN(FE_OFN153_HRESETn), 
	.Q(U_ctl_fr_wr_bcnt_5_), 
	.D(FE_PHN1002_U_ctl_n100), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_ctl_fr_wr_bcnt_reg_4_ (.RN(FE_OFN31_HRESETn), 
	.Q(U_ctl_fr_wr_bcnt_4_), 
	.D(FE_PHN3462_U_ctl_n101), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_ctl_fr_wr_bcnt_reg_3_ (.RN(FE_OFN153_HRESETn), 
	.Q(U_ctl_fr_wr_bcnt_3_), 
	.D(FE_PHN3451_U_ctl_n102), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_ctl_fr_wr_bcnt_reg_2_ (.RN(FE_OFN31_HRESETn), 
	.Q(U_ctl_fr_wr_bcnt_2_), 
	.D(FE_PHN3468_U_ctl_n103), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_ctl_fr_wr_bcnt_reg_1_ (.RN(FE_OFN31_HRESETn), 
	.Q(U_ctl_fr_wr_bcnt_1_), 
	.D(FE_PHN1225_U_ctl_n104), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_ctl_f_burst_done_reg (.RN(FE_OFN51_HRESETn), 
	.Q(U_ctl_f_burst_done), 
	.D(FE_PHN714_miu_burst_done), 
	.CK(hclk));
   DFFS_X2 U_ctl_fd_rd_ready_reg (.SN(FE_OFN153_HRESETn), 
	.Q(U_ctl_fd_rd_ready), 
	.D(FE_PHN1604_U_ctl_n106), 
	.CK(hclk));
   DFFS_X2 U_ctl_fd_df_push_n_reg (.SN(FE_OFN30_HRESETn), 
	.QN(m_df_push_n), 
	.D(FE_PHN5239_U_ctl_n299), 
	.CK(hclk));
   DFFS_X2 U_ctl_fd_zero_wait_ok_reg (.SN(FE_OFN55_HRESETn), 
	.QN(U_ctl_n151), 
	.D(FE_PHN4705_U_ctl_N89), 
	.CK(hclk));
   DFFS_X2 U_ctl_f_data_width_reg_0_ (.SN(FE_OFN55_HRESETn), 
	.Q(U_ctl_f_data_width_0_), 
	.D(FE_PHN848_U_ctl_n127), 
	.CK(hclk));
   DFFS_X2 U_ctl_f_col_width_reg_3_ (.SN(FE_OFN30_HRESETn), 
	.Q(U_ctl_f_col_width[3]), 
	.D(FE_PHN975_U_ctl_n132), 
	.CK(hclk));
   DFFS_X2 U_ctl_f_col_width_reg_1_ (.SN(FE_OFN30_HRESETn), 
	.Q(U_ctl_f_col_width[1]), 
	.D(FE_PHN1107_U_ctl_n134), 
	.CK(hclk));
   DFFS_X2 U_ctl_f_col_width_reg_0_ (.SN(FE_OFN55_HRESETn), 
	.Q(U_ctl_f_col_width[0]), 
	.D(FE_PHN1011_U_ctl_n135), 
	.CK(hclk));
   MUX2_X2 U_afifo_U_acore_U191 (.Z(hiu_addr[31]), 
	.S(FE_OFN250_U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_41_), 
	.A(U_afifo_U_acore_f_obuf_41_));
   MUX2_X2 U_afifo_U_acore_U190 (.Z(hiu_addr[30]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_40_), 
	.A(U_afifo_U_acore_f_obuf_40_));
   MUX2_X2 U_afifo_U_acore_U189 (.Z(hiu_addr[29]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_39_), 
	.A(U_afifo_U_acore_f_obuf_39_));
   MUX2_X2 U_afifo_U_acore_U188 (.Z(hiu_addr[28]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_38_), 
	.A(U_afifo_U_acore_f_obuf_38_));
   MUX2_X2 U_afifo_U_acore_U187 (.Z(hiu_addr[27]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_37_), 
	.A(U_afifo_U_acore_f_obuf_37_));
   MUX2_X2 U_afifo_U_acore_U186 (.Z(hiu_addr[26]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_36_), 
	.A(U_afifo_U_acore_f_obuf_36_));
   MUX2_X2 U_afifo_U_acore_U185 (.Z(hiu_addr[25]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_35_), 
	.A(U_afifo_U_acore_f_obuf_35_));
   MUX2_X2 U_afifo_U_acore_U184 (.Z(hiu_addr[24]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_34_), 
	.A(U_afifo_U_acore_f_obuf_34_));
   MUX2_X2 U_afifo_U_acore_U183 (.Z(hiu_addr[23]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_33_), 
	.A(U_afifo_U_acore_f_obuf_33_));
   MUX2_X2 U_afifo_U_acore_U182 (.Z(hiu_addr[22]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_32_), 
	.A(U_afifo_U_acore_f_obuf_32_));
   MUX2_X2 U_afifo_U_acore_U181 (.Z(hiu_addr[21]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_31_), 
	.A(U_afifo_U_acore_f_obuf_31_));
   MUX2_X2 U_afifo_U_acore_U180 (.Z(hiu_addr[20]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_30_), 
	.A(U_afifo_U_acore_f_obuf_30_));
   MUX2_X2 U_afifo_U_acore_U179 (.Z(hiu_addr[8]), 
	.S(U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_18_), 
	.A(U_afifo_U_acore_f_obuf_18_));
   MUX2_X2 U_afifo_U_acore_U178 (.Z(hiu_rw), 
	.S(FE_OFN250_U_afifo_U_acore_n1), 
	.B(U_afifo_U_acore_f_ibuf_2_), 
	.A(U_afifo_U_acore_f_obuf_2_));
   INV_X4 U_afifo_U_acore_U177 (.ZN(U_afifo_U_acore_n45), 
	.A(U_afifo_m_pop_n));
   OAI22_X1 U_afifo_U_acore_U176 (.ZN(U_afifo_U_acore_n_obuf_empty), 
	.B2(U_afifo_U_acore_n170), 
	.B1(U_afifo_m_pop_n), 
	.A2(FE_OFN26_U_afifo_U_acore_n38), 
	.A1(U_afifo_U_acore_n168));
   OAI21_X2 U_afifo_U_acore_U174 (.ZN(hiu_addr[16]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN1852_U_afifo_U_acore_n100), 
	.A(U_afifo_U_acore_n60));
   OAI21_X2 U_afifo_U_acore_U173 (.ZN(hiu_addr[12]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN3384_U_afifo_U_acore_n156), 
	.A(U_afifo_U_acore_n56));
   OAI21_X2 U_afifo_U_acore_U172 (.ZN(hiu_addr[13]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN3409_U_afifo_U_acore_n153), 
	.A(U_afifo_U_acore_n57));
   OAI21_X2 U_afifo_U_acore_U171 (.ZN(hiu_addr[10]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN3262_U_afifo_U_acore_n160), 
	.A(U_afifo_U_acore_n54));
   NOR2_X2 U_afifo_U_acore_U170 (.ZN(U_afifo_U_acore_n49), 
	.A2(U_afifo_U_acore_n44), 
	.A1(U_afifo_U_acore_n45));
   OAI211_X2 U_afifo_U_acore_U169 (.ZN(U_afifo_U_acore_n165), 
	.C2(U_afifo_U_acore_n64), 
	.C1(U_afifo_m_pop_n), 
	.B(FE_PHN815_U_afifo_U_acore_n11), 
	.A(U_afifo_U_acore_n169));
   OAI21_X1 U_afifo_U_acore_U168 (.ZN(U_afifo_U_acore_n65), 
	.B2(FE_PHN815_U_afifo_U_acore_n11), 
	.B1(U_afifo_U_acore_n166), 
	.A(FE_PHN3357_U_afifo_U_acore_f_afull));
   OAI21_X2 U_afifo_U_acore_U167 (.ZN(hiu_addr[15]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN1837_U_afifo_U_acore_n102), 
	.A(U_afifo_U_acore_n59));
   NAND2_X2 U_afifo_U_acore_U166 (.ZN(U_afifo_U_acore_n169), 
	.A2(FE_OFN250_U_afifo_U_acore_n1), 
	.A1(FE_PHN817_U_afifo_U_acore_n2));
   OAI21_X2 U_afifo_U_acore_U165 (.ZN(hiu_addr[9]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN3263_U_afifo_U_acore_n162), 
	.A(U_afifo_U_acore_n53));
   NOR2_X2 U_afifo_U_acore_U164 (.ZN(U_afifo_U_acore_n46), 
	.A2(FE_PHN761_U_afifo_U_acore_f_push_req_n), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   INV_X4 U_afifo_U_acore_U163 (.ZN(U_afifo_U_acore_n43), 
	.A(U_afifo_U_acore_n34));
   NAND2_X2 U_afifo_U_acore_U161 (.ZN(U_afifo_U_acore_n60), 
	.A2(U_afifo_U_acore_f_obuf_26_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   NAND2_X2 U_afifo_U_acore_U160 (.ZN(U_afifo_U_acore_n59), 
	.A2(U_afifo_U_acore_f_obuf_25_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   NAND2_X2 U_afifo_U_acore_U159 (.ZN(U_afifo_U_acore_n61), 
	.A2(U_afifo_U_acore_f_obuf_27_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   OAI21_X2 U_afifo_U_acore_U158 (.ZN(hiu_addr[17]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN1850_U_afifo_U_acore_n98), 
	.A(U_afifo_U_acore_n61));
   NAND2_X2 U_afifo_U_acore_U157 (.ZN(U_afifo_U_acore_n62), 
	.A2(U_afifo_U_acore_f_obuf_28_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   OAI21_X2 U_afifo_U_acore_U156 (.ZN(hiu_addr[18]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN1851_U_afifo_U_acore_n96), 
	.A(U_afifo_U_acore_n62));
   OAI21_X2 U_afifo_U_acore_U155 (.ZN(hiu_addr[19]), 
	.B2(U_afifo_U_acore_n43), 
	.B1(FE_PHN3248_U_afifo_U_acore_n94), 
	.A(U_afifo_U_acore_n63));
   NAND2_X2 U_afifo_U_acore_U154 (.ZN(U_afifo_U_acore_n56), 
	.A2(U_afifo_U_acore_f_obuf_22_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   NAND2_X2 U_afifo_U_acore_U153 (.ZN(U_afifo_U_acore_n57), 
	.A2(U_afifo_U_acore_f_obuf_23_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   NAND2_X2 U_afifo_U_acore_U152 (.ZN(U_afifo_U_acore_n55), 
	.A2(U_afifo_U_acore_f_obuf_21_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   NAND2_X2 U_afifo_U_acore_U151 (.ZN(U_afifo_U_acore_n58), 
	.A2(U_afifo_U_acore_f_obuf_24_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   NOR2_X2 U_afifo_U_acore_U150 (.ZN(U_afifo_m_empty), 
	.A2(U_afifo_U_acore_n169), 
	.A1(FE_PHN815_U_afifo_U_acore_n11));
   INV_X4 U_afifo_U_acore_U149 (.ZN(U_afifo_U_acore_n64), 
	.A(FE_PHN817_U_afifo_U_acore_n2));
   NAND2_X2 U_afifo_U_acore_U148 (.ZN(U_afifo_U_acore_n66), 
	.A2(FE_PHN815_U_afifo_U_acore_n11), 
	.A1(U_afifo_U_acore_n64));
   NAND2_X2 U_afifo_U_acore_U147 (.ZN(U_afifo_m_afull), 
	.A2(U_afifo_U_acore_n12), 
	.A1(U_afifo_U_acore_n66));
   NAND2_X2 U_afifo_U_acore_U146 (.ZN(U_afifo_U_acore_n54), 
	.A2(U_afifo_U_acore_f_obuf_20_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   NAND2_X2 U_afifo_U_acore_U145 (.ZN(U_afifo_U_acore_n53), 
	.A2(U_afifo_U_acore_f_obuf_19_), 
	.A1(FE_OFN197_U_afifo_U_acore_n38));
   NOR2_X2 U_afifo_U_acore_U144 (.ZN(U_afifo_m_aempty), 
	.A2(U_afifo_U_acore_n46), 
	.A1(U_afifo_U_acore_n64));
   AOI22_X2 U_afifo_U_acore_U143 (.ZN(U_afifo_U_acore_n164), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[18]), 
	.A2(U_afifo_U_acore_f_obuf_18_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U142 (.ZN(U_afifo_U_acore_n95), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[28]), 
	.A2(U_afifo_U_acore_f_obuf_28_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U141 (.ZN(U_afifo_U_acore_n97), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[27]), 
	.A2(U_afifo_U_acore_f_obuf_27_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U140 (.ZN(U_afifo_U_acore_n101), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[25]), 
	.A2(U_afifo_U_acore_f_obuf_25_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U139 (.ZN(U_afifo_U_acore_n93), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[29]), 
	.A2(U_afifo_U_acore_f_obuf_29_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U138 (.ZN(U_afifo_U_acore_n99), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[26]), 
	.A2(U_afifo_U_acore_f_obuf_26_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U137 (.ZN(U_afifo_U_acore_n103), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[24]), 
	.A2(U_afifo_U_acore_f_obuf_24_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U136 (.ZN(U_afifo_U_acore_n143), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[23]), 
	.A2(U_afifo_U_acore_f_obuf_23_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U135 (.ZN(U_afifo_U_acore_n155), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[22]), 
	.A2(U_afifo_U_acore_f_obuf_22_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U134 (.ZN(U_afifo_U_acore_n159), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[20]), 
	.A2(U_afifo_U_acore_f_obuf_20_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U133 (.ZN(U_afifo_U_acore_n161), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[19]), 
	.A2(U_afifo_U_acore_f_obuf_19_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U132 (.ZN(U_afifo_U_acore_n157), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[21]), 
	.A2(U_afifo_U_acore_f_obuf_21_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U131 (.ZN(U_afifo_U_acore_n75), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[37]), 
	.A2(U_afifo_U_acore_f_obuf_37_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U130 (.ZN(U_afifo_U_acore_n77), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[36]), 
	.A2(U_afifo_U_acore_f_obuf_36_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U129 (.ZN(U_afifo_U_acore_n73), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[38]), 
	.A2(U_afifo_U_acore_f_obuf_38_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U128 (.ZN(U_afifo_U_acore_n71), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[39]), 
	.A2(U_afifo_U_acore_f_obuf_39_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X2 U_afifo_U_acore_U127 (.ZN(U_afifo_U_acore_n196), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[17]), 
	.A2(U_afifo_U_acore_f_obuf_17_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U126 (.ZN(U_afifo_U_acore_n198), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[16]), 
	.A2(U_afifo_U_acore_f_obuf_16_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U125 (.ZN(U_afifo_U_acore_n200), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[15]), 
	.A2(U_afifo_U_acore_f_obuf_15_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U124 (.ZN(U_afifo_U_acore_n202), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[14]), 
	.A2(U_afifo_U_acore_f_obuf_14_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U123 (.ZN(U_afifo_U_acore_n209), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[0]), 
	.A2(U_afifo_U_acore_f_obuf_0_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U122 (.ZN(U_afifo_U_acore_n204), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[13]), 
	.A2(U_afifo_U_acore_f_obuf_13_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U121 (.ZN(U_afifo_U_acore_n206), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[12]), 
	.A2(U_afifo_U_acore_f_obuf_12_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U120 (.ZN(U_afifo_U_acore_n191), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[43]), 
	.A2(U_afifo_U_acore_f_obuf_43_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U119 (.ZN(U_afifo_U_acore_n208), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[11]), 
	.A2(U_afifo_U_acore_f_obuf_11_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U118 (.ZN(U_afifo_U_acore_n187), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[46]), 
	.A2(U_afifo_U_acore_f_obuf_46_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U117 (.ZN(U_afifo_U_acore_n185), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[47]), 
	.A2(U_afifo_U_acore_f_obuf_47_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U116 (.ZN(U_afifo_U_acore_n193), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[42]), 
	.A2(U_afifo_U_acore_f_obuf_42_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U115 (.ZN(U_afifo_U_acore_n195), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[3]), 
	.A2(U_afifo_U_acore_f_obuf_3_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U114 (.ZN(U_afifo_U_acore_n178), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[5]), 
	.A2(U_afifo_U_acore_f_obuf_5_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U113 (.ZN(U_afifo_U_acore_n189), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[44]), 
	.A2(U_afifo_U_acore_f_obuf_44_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U112 (.ZN(U_afifo_U_acore_n180), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[4]), 
	.A2(U_afifo_U_acore_f_obuf_4_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U111 (.ZN(U_afifo_U_acore_n171), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[9]), 
	.A2(U_afifo_U_acore_f_obuf_9_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U110 (.ZN(U_afifo_U_acore_n188), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[45]), 
	.A2(U_afifo_U_acore_f_obuf_45_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U109 (.ZN(U_afifo_U_acore_n183), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[48]), 
	.A2(U_afifo_U_acore_f_obuf_48_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U108 (.ZN(U_afifo_U_acore_n174), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[7]), 
	.A2(U_afifo_U_acore_f_obuf_7_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U107 (.ZN(U_afifo_U_acore_n182), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[49]), 
	.A2(U_afifo_U_acore_f_obuf_49_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U106 (.ZN(U_afifo_U_acore_n176), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[6]), 
	.A2(U_afifo_U_acore_f_obuf_6_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U105 (.ZN(U_afifo_U_acore_n172), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[8]), 
	.A2(U_afifo_U_acore_f_obuf_8_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U104 (.ZN(U_afifo_U_acore_n67), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[41]), 
	.A2(U_afifo_U_acore_f_obuf_41_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U103 (.ZN(U_afifo_U_acore_n69), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[40]), 
	.A2(U_afifo_U_acore_f_obuf_40_), 
	.A1(U_afifo_U_acore_n39));
   AOI22_X2 U_afifo_U_acore_U102 (.ZN(U_afifo_U_acore_n91), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[2]), 
	.A2(U_afifo_U_acore_f_obuf_2_), 
	.A1(U_afifo_U_acore_n39));
   OAI211_X1 U_afifo_U_acore_U101 (.ZN(U_afifo_U_acore_n_afull), 
	.C2(U_afifo_U_acore_n66), 
	.C1(U_afifo_U_acore_n45), 
	.B(U_afifo_U_acore_m_sf_full), 
	.A(U_afifo_U_acore_n65));
   INV_X8 U_afifo_U_acore_U99 (.ZN(U_afifo_U_acore_n163), 
	.A(U_afifo_U_acore_n166));
   OAI21_X4 U_afifo_U_acore_U96 (.ZN(hiu_burst_size[3]), 
	.B2(U_afifo_U_acore_n7), 
	.B1(U_afifo_U_acore_n1), 
	.A(U_afifo_U_acore_n51));
   NOR2_X2 U_afifo_U_acore_U94 (.ZN(U_afifo_U_acore_n168), 
	.A2(U_afifo_U_acore_n48), 
	.A1(U_afifo_U_acore_n49));
   NAND2_X2 U_afifo_U_acore_U93 (.ZN(U_afifo_U_acore_n211), 
	.A2(FE_PHN817_U_afifo_U_acore_n2), 
	.A1(U_afifo_U_acore_n168));
   INV_X4 U_afifo_U_acore_U92 (.ZN(U_afifo_U_acore_n1), 
	.A(U_afifo_U_acore_n43));
   OAI21_X1 U_afifo_U_acore_U91 (.ZN(U_afifo_m_full), 
	.B2(U_afifo_U_acore_n12), 
	.B1(FE_PHN761_U_afifo_U_acore_f_push_req_n), 
	.A(U_afifo_U_acore_m_sf_full));
   NAND2_X1 U_afifo_U_acore_U90 (.ZN(U_afifo_U_acore_n170), 
	.A2(FE_PHN761_U_afifo_U_acore_f_push_req_n), 
	.A1(FE_PHN817_U_afifo_U_acore_n2));
   OR2_X2 U_afifo_U_acore_U89 (.ZN(U_afifo_U_acore_n51), 
	.A2(FE_OFN26_U_afifo_U_acore_n38), 
	.A1(FE_PHN1560_U_afifo_U_acore_n175));
   NOR2_X1 U_afifo_U_acore_U86 (.ZN(U_afifo_U_acore_n44), 
	.A2(U_afifo_U_acore_n169), 
	.A1(FE_PHN761_U_afifo_U_acore_f_push_req_n));
   NOR2_X1 U_afifo_U_acore_U85 (.ZN(U_afifo_U_acore_n48), 
	.A2(U_afifo_U_acore_n47), 
	.A1(U_afifo_m_pop_n));
   NAND2_X2 U_afifo_U_acore_U84 (.ZN(U_afifo_U_acore_n166), 
	.A2(U_afifo_U_acore_n45), 
	.A1(U_afifo_U_acore_n64));
   INV_X4 U_afifo_U_acore_U83 (.ZN(U_afifo_U_acore_n39), 
	.A(U_afifo_U_acore_n168));
   INV_X4 U_afifo_U_acore_U82 (.ZN(U_afifo_U_acore_n40), 
	.A(U_afifo_U_acore_n168));
   OAI21_X1 U_afifo_U_acore_U80 (.ZN(U_afifo_U_acore_n116), 
	.B2(FE_PHN1558_U_afifo_U_acore_n190), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3367_U_afifo_U_acore_n189));
   OAI21_X1 U_afifo_U_acore_U79 (.ZN(U_afifo_U_acore_n151), 
	.B2(FE_PHN1849_U_afifo_U_acore_n207), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3350_U_afifo_U_acore_n206));
   OAI21_X1 U_afifo_U_acore_U78 (.ZN(U_afifo_U_acore_n147), 
	.B2(FE_PHN3243_U_afifo_U_acore_n199), 
	.B1(U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n198));
   OAI21_X1 U_afifo_U_acore_U77 (.ZN(U_afifo_U_acore_n117), 
	.B2(FE_PHN1563_U_afifo_U_acore_n192), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3344_U_afifo_U_acore_n191));
   OAI21_X1 U_afifo_U_acore_U76 (.ZN(U_afifo_U_acore_n154), 
	.B2(FE_PHN1836_U_afifo_U_acore_n210), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3361_U_afifo_U_acore_n209));
   OAI21_X1 U_afifo_U_acore_U75 (.ZN(U_afifo_U_acore_n110), 
	.B2(FE_PHN1847_U_afifo_U_acore_n181), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3366_U_afifo_U_acore_n180));
   OAI21_X1 U_afifo_U_acore_U74 (.ZN(U_afifo_U_acore_n149), 
	.B2(FE_PHN1839_U_afifo_U_acore_n203), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3348_U_afifo_U_acore_n202));
   OAI21_X1 U_afifo_U_acore_U73 (.ZN(U_afifo_U_acore_n152), 
	.B2(U_afifo_U_acore_n31), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3336_U_afifo_U_acore_n208));
   OAI21_X1 U_afifo_U_acore_U72 (.ZN(U_afifo_U_acore_n109), 
	.B2(FE_PHN1554_U_afifo_U_acore_n179), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3335_U_afifo_U_acore_n178));
   OAI21_X1 U_afifo_U_acore_U71 (.ZN(U_afifo_U_acore_n150), 
	.B2(FE_PHN1561_U_afifo_U_acore_n205), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3331_U_afifo_U_acore_n204));
   OAI21_X1 U_afifo_U_acore_U70 (.ZN(U_afifo_U_acore_n148), 
	.B2(FE_PHN1844_U_afifo_U_acore_n201), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3376_U_afifo_U_acore_n200));
   OAI21_X1 U_afifo_U_acore_U69 (.ZN(U_afifo_U_acore_n115), 
	.B2(U_afifo_U_acore_n30), 
	.B1(U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n188));
   OAI21_X1 U_afifo_U_acore_U68 (.ZN(U_afifo_U_acore_n107), 
	.B2(FE_PHN1560_U_afifo_U_acore_n175), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3359_U_afifo_U_acore_n174));
   OAI21_X1 U_afifo_U_acore_U67 (.ZN(U_afifo_U_acore_n114), 
	.B2(FE_PHN3423_U_afifo_U_acore_n29), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3356_U_afifo_U_acore_n187));
   OAI21_X1 U_afifo_U_acore_U66 (.ZN(U_afifo_U_acore_n111), 
	.B2(U_afifo_U_acore_n28), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3360_U_afifo_U_acore_n182));
   OAI21_X1 U_afifo_U_acore_U65 (.ZN(U_afifo_U_acore_n146), 
	.B2(FE_PHN1835_U_afifo_U_acore_n197), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3342_U_afifo_U_acore_n196));
   OAI21_X1 U_afifo_U_acore_U64 (.ZN(U_afifo_U_acore_n108), 
	.B2(FE_PHN1834_U_afifo_U_acore_n177), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3333_U_afifo_U_acore_n176));
   OAI21_X1 U_afifo_U_acore_U63 (.ZN(U_afifo_U_acore_n121), 
	.B2(FE_PHN3261_U_afifo_U_acore_n33), 
	.B1(U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n195));
   OAI21_X1 U_afifo_U_acore_U62 (.ZN(U_afifo_U_acore_n112), 
	.B2(FE_PHN1841_U_afifo_U_acore_n184), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3369_U_afifo_U_acore_n183));
   OAI21_X1 U_afifo_U_acore_U61 (.ZN(U_afifo_U_acore_n118), 
	.B2(FE_PHN1840_U_afifo_U_acore_n194), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3362_U_afifo_U_acore_n193));
   OAI21_X1 U_afifo_U_acore_U60 (.ZN(U_afifo_U_acore_n120), 
	.B2(FE_PHN1186_U_afifo_U_acore_n70), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3457_U_afifo_U_acore_n69));
   OAI21_X1 U_afifo_U_acore_U59 (.ZN(U_afifo_U_acore_n113), 
	.B2(FE_PHN1564_U_afifo_U_acore_n186), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3340_U_afifo_U_acore_n185));
   OAI21_X1 U_afifo_U_acore_U58 (.ZN(U_afifo_U_acore_n106), 
	.B2(FE_PHN1408_U_afifo_U_acore_n173), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3347_U_afifo_U_acore_n172));
   OAI21_X1 U_afifo_U_acore_U57 (.ZN(U_afifo_U_acore_n105), 
	.B2(U_afifo_U_acore_n32), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3365_U_afifo_U_acore_n171));
   OAI21_X1 U_afifo_U_acore_U56 (.ZN(U_afifo_U_acore_n119), 
	.B2(U_afifo_U_acore_n211), 
	.B1(FE_PHN1192_U_afifo_U_acore_n68), 
	.A(FE_PHN3416_U_afifo_U_acore_n67));
   OAI21_X1 U_afifo_U_acore_U55 (.ZN(U_afifo_U_acore_n132), 
	.B2(FE_PHN1404_U_afifo_U_acore_n92), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3459_U_afifo_U_acore_n91));
   OAI21_X1 U_afifo_U_acore_U54 (.ZN(U_afifo_U_acore_n135), 
	.B2(FE_PHN1850_U_afifo_U_acore_n98), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN4719_U_afifo_U_acore_n97));
   OAI21_X1 U_afifo_U_acore_U53 (.ZN(U_afifo_U_acore_n134), 
	.B2(FE_PHN1851_U_afifo_U_acore_n96), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3323_U_afifo_U_acore_n95));
   OAI21_X1 U_afifo_U_acore_U52 (.ZN(U_afifo_U_acore_n136), 
	.B2(FE_PHN1852_U_afifo_U_acore_n100), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3406_U_afifo_U_acore_n99));
   OAI21_X1 U_afifo_U_acore_U51 (.ZN(U_afifo_U_acore_n133), 
	.B2(FE_PHN3248_U_afifo_U_acore_n94), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n93));
   OAI21_X1 U_afifo_U_acore_U50 (.ZN(U_afifo_U_acore_n137), 
	.B2(FE_PHN1837_U_afifo_U_acore_n102), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3447_U_afifo_U_acore_n101));
   OAI21_X1 U_afifo_U_acore_U49 (.ZN(U_afifo_U_acore_n145), 
	.B2(FE_PHN1189_U_afifo_U_acore_n167), 
	.B1(U_afifo_U_acore_n211), 
	.A(FE_PHN3455_U_afifo_U_acore_n164));
   OAI21_X1 U_afifo_U_acore_U48 (.ZN(U_afifo_U_acore_n138), 
	.B2(FE_PHN3257_U_afifo_U_acore_n104), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n103));
   OAI21_X1 U_afifo_U_acore_U47 (.ZN(U_afifo_U_acore_n144), 
	.B2(FE_PHN3263_U_afifo_U_acore_n162), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n161));
   OAI21_X1 U_afifo_U_acore_U46 (.ZN(U_afifo_U_acore_n142), 
	.B2(FE_PHN3262_U_afifo_U_acore_n160), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n159));
   OAI21_X1 U_afifo_U_acore_U45 (.ZN(U_afifo_U_acore_n139), 
	.B2(FE_PHN3409_U_afifo_U_acore_n153), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3430_U_afifo_U_acore_n143));
   OAI21_X1 U_afifo_U_acore_U44 (.ZN(U_afifo_U_acore_n141), 
	.B2(FE_PHN3412_U_afifo_U_acore_n158), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3460_U_afifo_U_acore_n157));
   OAI21_X1 U_afifo_U_acore_U43 (.ZN(U_afifo_U_acore_n140), 
	.B2(FE_PHN3384_U_afifo_U_acore_n156), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3433_U_afifo_U_acore_n155));
   OAI21_X1 U_afifo_U_acore_U42 (.ZN(U_afifo_U_acore_n131), 
	.B2(FE_PHN1405_U_afifo_U_acore_n90), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3448_U_afifo_U_acore_n89));
   OAI21_X1 U_afifo_U_acore_U41 (.ZN(U_afifo_U_acore_n130), 
	.B2(FE_PHN1193_U_afifo_U_acore_n88), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3444_U_afifo_U_acore_n87));
   OAI21_X1 U_afifo_U_acore_U40 (.ZN(U_afifo_U_acore_n127), 
	.B2(FE_PHN1187_U_afifo_U_acore_n82), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n81));
   OAI21_X1 U_afifo_U_acore_U39 (.ZN(U_afifo_U_acore_n129), 
	.B2(FE_PHN1188_U_afifo_U_acore_n86), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n85));
   OAI21_X1 U_afifo_U_acore_U38 (.ZN(U_afifo_U_acore_n126), 
	.B2(FE_PHN1552_U_afifo_U_acore_n80), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n79));
   OAI21_X1 U_afifo_U_acore_U37 (.ZN(U_afifo_U_acore_n128), 
	.B2(FE_PHN1190_U_afifo_U_acore_n84), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(U_afifo_U_acore_n83));
   NAND2_X1 U_afifo_U_acore_U36 (.ZN(U_afifo_U_acore_n63), 
	.A2(U_afifo_U_acore_f_obuf_29_), 
	.A1(FE_OFN26_U_afifo_U_acore_n38));
   INV_X2 U_afifo_U_acore_U35 (.ZN(U_afifo_U_acore_n47), 
	.A(U_afifo_m_aempty));
   AOI22_X1 U_afifo_U_acore_U34 (.ZN(U_afifo_U_acore_n87), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[31]), 
	.A2(U_afifo_U_acore_f_obuf_31_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X1 U_afifo_U_acore_U33 (.ZN(U_afifo_U_acore_n85), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[32]), 
	.A2(U_afifo_U_acore_f_obuf_32_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X1 U_afifo_U_acore_U32 (.ZN(U_afifo_U_acore_n83), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[33]), 
	.A2(U_afifo_U_acore_f_obuf_33_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X1 U_afifo_U_acore_U31 (.ZN(U_afifo_U_acore_n81), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[34]), 
	.A2(FE_PHN3465_U_afifo_U_acore_f_obuf_34_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X1 U_afifo_U_acore_U30 (.ZN(U_afifo_U_acore_n79), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[35]), 
	.A2(U_afifo_U_acore_f_obuf_35_), 
	.A1(U_afifo_U_acore_n40));
   AOI22_X1 U_afifo_U_acore_U29 (.ZN(U_afifo_U_acore_n89), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_data_out[30]), 
	.A2(U_afifo_U_acore_f_obuf_30_), 
	.A1(U_afifo_U_acore_n40));
   OAI21_X2 U_afifo_U_acore_U28 (.ZN(U_afifo_U_acore_n125), 
	.B2(FE_PHN1191_U_afifo_U_acore_n78), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3401_U_afifo_U_acore_n77));
   OAI21_X2 U_afifo_U_acore_U27 (.ZN(U_afifo_U_acore_n123), 
	.B2(FE_PHN1194_U_afifo_U_acore_n74), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3380_U_afifo_U_acore_n73));
   OAI21_X2 U_afifo_U_acore_U26 (.ZN(U_afifo_U_acore_n124), 
	.B2(FE_PHN1406_U_afifo_U_acore_n76), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3453_U_afifo_U_acore_n75));
   OAI21_X2 U_afifo_U_acore_U25 (.ZN(U_afifo_U_acore_n122), 
	.B2(FE_PHN1197_U_afifo_U_acore_n72), 
	.B1(FE_OFN247_U_afifo_U_acore_n211), 
	.A(FE_PHN3386_U_afifo_U_acore_n71));
   OAI22_X1 U_afifo_U_acore_U24 (.ZN(hiu_addr[7]), 
	.B2(FE_PHN1835_U_afifo_U_acore_n197), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n19), 
	.A1(U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U23 (.ZN(hiu_addr[2]), 
	.B2(FE_PHN1849_U_afifo_U_acore_n207), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n15), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U22 (.ZN(hiu_haddr[0]), 
	.B2(U_afifo_U_acore_n30), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n21), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U21 (.ZN(hiu_addr[6]), 
	.B2(FE_PHN3243_U_afifo_U_acore_n199), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n18), 
	.A1(U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U20 (.ZN(hiu_haddr[1]), 
	.B2(FE_PHN3423_U_afifo_U_acore_n29), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n22), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U19 (.ZN(hiu_addr[5]), 
	.B2(FE_PHN1844_U_afifo_U_acore_n201), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n17), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U18 (.ZN(hiu_addr[1]), 
	.B2(U_afifo_U_acore_n31), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n14), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U17 (.ZN(U_afifo_m_data_out_49), 
	.B2(U_afifo_U_acore_n28), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n10), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U16 (.ZN(hiu_hsize[1]), 
	.B2(FE_PHN1563_U_afifo_U_acore_n192), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n26), 
	.A1(U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U15 (.ZN(hiu_hsize[2]), 
	.B2(FE_PHN1558_U_afifo_U_acore_n190), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n27), 
	.A1(U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U14 (.ZN(U_afifo_m_data_out_3), 
	.B2(FE_PHN3261_U_afifo_U_acore_n33), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n25), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U13 (.ZN(U_afifo_m_data_out_0_), 
	.B2(FE_PHN1836_U_afifo_U_acore_n210), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n3), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U12 (.ZN(hiu_hsize[0]), 
	.B2(FE_PHN1840_U_afifo_U_acore_n194), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n20), 
	.A1(U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U11 (.ZN(hiu_addr[4]), 
	.B2(FE_PHN1839_U_afifo_U_acore_n203), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n9), 
	.A1(U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U10 (.ZN(hiu_addr[3]), 
	.B2(FE_PHN1561_U_afifo_U_acore_n205), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n16), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X2 U_afifo_U_acore_U9 (.ZN(hiu_burst_size[1]), 
	.B2(FE_PHN1554_U_afifo_U_acore_n179), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n5), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X2 U_afifo_U_acore_U8 (.ZN(hiu_burst_size[2]), 
	.B2(FE_PHN1834_U_afifo_U_acore_n177), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n6), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U7 (.ZN(hiu_haddr[2]), 
	.B2(FE_PHN1564_U_afifo_U_acore_n186), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n23), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X2 U_afifo_U_acore_U6 (.ZN(hiu_burst_size[4]), 
	.B2(FE_PHN1408_U_afifo_U_acore_n173), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n13), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI22_X1 U_afifo_U_acore_U5 (.ZN(hiu_haddr[3]), 
	.B2(FE_PHN1841_U_afifo_U_acore_n184), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n24), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   OAI21_X2 U_afifo_U_acore_U4 (.ZN(hiu_addr[14]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN3257_U_afifo_U_acore_n104), 
	.A(U_afifo_U_acore_n58));
   OAI21_X2 U_afifo_U_acore_U3 (.ZN(hiu_addr[11]), 
	.B2(FE_OFN197_U_afifo_U_acore_n38), 
	.B1(FE_PHN3412_U_afifo_U_acore_n158), 
	.A(U_afifo_U_acore_n55));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_5_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_n179), 
	.D(FE_PHN1239_U_afifo_m_data_in_5_), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_6_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_n177), 
	.D(U_afifo_m_data_in[6]), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_7_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_n175), 
	.D(FE_PHN1907_U_afifo_m_data_in_7_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_8_ (.RN(FE_OFN191_HRESETn), 
	.QN(U_afifo_U_acore_n173), 
	.D(U_afifo_m_data_in[8]), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_44_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n190), 
	.D(U_afifo_m_data_in[44]), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_0_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_n210), 
	.D(U_afifo_m_data_in[0]), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_43_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n192), 
	.D(FE_PHN1686_U_afifo_m_data_in_43_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_18_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n167), 
	.Q(U_afifo_U_acore_f_ibuf_18_), 
	.D(U_afifo_m_data_in[18]), 
	.CK(HCLK__L5_N37));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_15_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n201), 
	.D(FE_PHN1622_U_afifo_m_data_in_15_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_14_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n203), 
	.D(FE_PHN1618_U_afifo_m_data_in_14_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_47_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_n186), 
	.D(U_afifo_m_data_in[47]), 
	.CK(HCLK__L5_N34));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_48_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_n184), 
	.D(FE_PHN1616_U_afifo_m_data_in_48_), 
	.CK(HCLK__L5_N34));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_2_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_n92), 
	.Q(U_afifo_U_acore_f_ibuf_2_), 
	.D(FE_PHN1687_U_afifo_m_data_in_2_), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_19_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n162), 
	.D(FE_PHN1786_U_afifo_m_data_in_19_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_20_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_n160), 
	.D(FE_PHN1769_U_afifo_m_data_in_20_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_21_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_n158), 
	.D(FE_PHN1749_U_afifo_m_data_in_21_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_22_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_n156), 
	.D(U_afifo_m_data_in[22]), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_23_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n153), 
	.D(FE_PHN1685_U_afifo_m_data_in_23_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_24_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n104), 
	.D(FE_PHN1688_U_afifo_m_data_in_24_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_25_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_n102), 
	.D(U_afifo_m_data_in[25]), 
	.CK(HCLK__L5_N37));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_26_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_n100), 
	.D(U_afifo_m_data_in[26]), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_27_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_n98), 
	.D(FE_PHN1818_U_afifo_m_data_in_27_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_28_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_n96), 
	.D(FE_PHN1789_U_afifo_m_data_in_28_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_29_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n94), 
	.D(FE_PHN1515_U_afifo_m_data_in_29_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_30_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_n90), 
	.Q(U_afifo_U_acore_f_ibuf_30_), 
	.D(FE_PHN1750_U_afifo_m_data_in_30_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_31_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_n88), 
	.Q(U_afifo_U_acore_f_ibuf_31_), 
	.D(FE_PHN1763_U_afifo_m_data_in_31_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_32_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_n86), 
	.Q(U_afifo_U_acore_f_ibuf_32_), 
	.D(FE_PHN1178_U_afifo_m_data_in_32_), 
	.CK(HCLK__L5_N37));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_33_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_n84), 
	.Q(U_afifo_U_acore_f_ibuf_33_), 
	.D(FE_PHN1783_U_afifo_m_data_in_33_), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_34_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_n82), 
	.Q(U_afifo_U_acore_f_ibuf_34_), 
	.D(U_afifo_m_data_in[34]), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_35_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n80), 
	.Q(U_afifo_U_acore_f_ibuf_35_), 
	.D(U_afifo_m_data_in[35]), 
	.CK(HCLK__L5_N39));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_36_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_n78), 
	.Q(U_afifo_U_acore_f_ibuf_36_), 
	.D(U_afifo_m_data_in[36]), 
	.CK(HCLK__L5_N37));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_37_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n76), 
	.Q(U_afifo_U_acore_f_ibuf_37_), 
	.D(U_afifo_m_data_in[37]), 
	.CK(HCLK__L5_N37));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_38_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n74), 
	.Q(U_afifo_U_acore_f_ibuf_38_), 
	.D(FE_PHN1513_U_afifo_m_data_in_38_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_39_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_n72), 
	.Q(U_afifo_U_acore_f_ibuf_39_), 
	.D(U_afifo_m_data_in[39]), 
	.CK(HCLK__L5_N33));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_40_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n70), 
	.Q(U_afifo_U_acore_f_ibuf_40_), 
	.D(U_afifo_m_data_in[40]), 
	.CK(HCLK__L5_N37));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_41_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_n68), 
	.Q(U_afifo_U_acore_f_ibuf_41_), 
	.D(U_afifo_m_data_in[41]), 
	.CK(HCLK__L5_N33));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_42_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_n194), 
	.D(FE_PHN1373_U_afifo_m_data_in_42_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_17_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n197), 
	.D(FE_PHN1621_U_afifo_m_data_in_17_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_13_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_n205), 
	.D(U_afifo_m_data_in[13]), 
	.CK(HCLK__L5_N34));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_16_ (.RN(FE_OFN169_HRESETn), 
	.QN(U_afifo_U_acore_n199), 
	.D(FE_PHN1620_U_afifo_m_data_in_16_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_12_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n207), 
	.D(FE_PHN1374_U_afifo_m_data_in_12_), 
	.CK(HCLK__L5_N38));
   DFFR_X2 U_afifo_U_acore_f_ibuf_reg_4_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_U_acore_n181), 
	.D(FE_PHN1238_U_afifo_m_data_in_4_), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_f_afull_reg (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_n12), 
	.Q(U_afifo_U_acore_f_afull), 
	.D(FE_PHN962_U_afifo_U_acore_n_afull), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_9_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_n8), 
	.Q(U_afifo_U_acore_f_obuf_9_), 
	.D(FE_PHN1312_U_afifo_U_acore_n105), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_8_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_n13), 
	.Q(U_afifo_U_acore_f_obuf_8_), 
	.D(FE_PHN1278_U_afifo_U_acore_n106), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_7_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n7), 
	.Q(U_afifo_U_acore_f_obuf_7_), 
	.D(FE_PHN1280_U_afifo_U_acore_n107), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_6_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_afifo_U_acore_n6), 
	.Q(U_afifo_U_acore_f_obuf_6_), 
	.D(FE_PHN1286_U_afifo_U_acore_n108), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_5_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_n5), 
	.Q(U_afifo_U_acore_f_obuf_5_), 
	.D(FE_PHN1289_U_afifo_U_acore_n109), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_4_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_n4), 
	.Q(U_afifo_U_acore_f_obuf_4_), 
	.D(FE_PHN1307_U_afifo_U_acore_n110), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_49_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_U_acore_n10), 
	.Q(U_afifo_U_acore_f_obuf_49_), 
	.D(FE_PHN1298_U_afifo_U_acore_n111), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_48_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_n24), 
	.Q(U_afifo_U_acore_f_obuf_48_), 
	.D(FE_PHN1293_U_afifo_U_acore_n112), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_47_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_afifo_U_acore_n23), 
	.Q(U_afifo_U_acore_f_obuf_47_), 
	.D(FE_PHN1277_U_afifo_U_acore_n113), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_46_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_U_acore_n22), 
	.Q(U_afifo_U_acore_f_obuf_46_), 
	.D(FE_PHN1297_U_afifo_U_acore_n114), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_45_ (.RN(FE_OFN171_HRESETn), 
	.QN(U_afifo_U_acore_n21), 
	.Q(U_afifo_U_acore_f_obuf_45_), 
	.D(FE_PHN1304_U_afifo_U_acore_n115), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_44_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n27), 
	.Q(U_afifo_U_acore_f_obuf_44_), 
	.D(FE_PHN1272_U_afifo_U_acore_n116), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_43_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n26), 
	.Q(U_afifo_U_acore_f_obuf_43_), 
	.D(FE_PHN1285_U_afifo_U_acore_n117), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_42_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n20), 
	.Q(U_afifo_U_acore_f_obuf_42_), 
	.D(FE_PHN1302_U_afifo_U_acore_n118), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_41_ (.RN(FE_OFN35_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_41_), 
	.D(FE_PHN1257_U_afifo_U_acore_n119), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_40_ (.RN(FE_OFN47_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_40_), 
	.D(FE_PHN1266_U_afifo_U_acore_n120), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_3_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_n25), 
	.Q(U_afifo_U_acore_f_obuf_3_), 
	.D(FE_PHN1309_U_afifo_U_acore_n121), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_39_ (.RN(FE_OFN149_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_39_), 
	.D(FE_PHN1259_U_afifo_U_acore_n122), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_38_ (.RN(FE_OFN32_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_38_), 
	.D(FE_PHN1260_U_afifo_U_acore_n123), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_37_ (.RN(FE_OFN58_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_37_), 
	.D(FE_PHN1263_U_afifo_U_acore_n124), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_36_ (.RN(FE_OFN58_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_36_), 
	.D(FE_PHN1258_U_afifo_U_acore_n125), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_35_ (.RN(FE_OFN47_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_35_), 
	.D(FE_PHN1274_U_afifo_U_acore_n126), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_34_ (.RN(FE_OFN29_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_34_), 
	.D(FE_PHN1267_U_afifo_U_acore_n127), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_33_ (.RN(FE_OFN58_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_33_), 
	.D(FE_PHN1273_U_afifo_U_acore_n128), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_32_ (.RN(FE_OFN58_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_32_), 
	.D(FE_PHN1261_U_afifo_U_acore_n129), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_31_ (.RN(FE_OFN58_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_31_), 
	.D(FE_PHN1281_U_afifo_U_acore_n130), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_30_ (.RN(FE_OFN58_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_30_), 
	.D(FE_PHN1270_U_afifo_U_acore_n131), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_2_ (.RN(FE_OFN31_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_2_), 
	.D(FE_PHN1264_U_afifo_U_acore_n132), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_29_ (.RN(FE_OFN47_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_29_), 
	.D(FE_PHN3180_U_afifo_U_acore_n133), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_28_ (.RN(FE_OFN58_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_28_), 
	.D(FE_PHN1319_U_afifo_U_acore_n134), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_27_ (.RN(FE_OFN58_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_27_), 
	.D(FE_PHN1316_U_afifo_U_acore_n135), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_26_ (.RN(FE_OFN58_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_26_), 
	.D(FE_PHN1317_U_afifo_U_acore_n136), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_25_ (.RN(FE_OFN149_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_25_), 
	.D(FE_PHN1308_U_afifo_U_acore_n137), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_24_ (.RN(FE_OFN35_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_24_), 
	.D(FE_PHN1325_U_afifo_U_acore_n138), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_23_ (.RN(FE_OFN149_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_23_), 
	.D(FE_PHN1324_U_afifo_U_acore_n139), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_22_ (.RN(FE_OFN149_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_22_), 
	.D(FE_PHN1318_U_afifo_U_acore_n140), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_21_ (.RN(FE_OFN149_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_21_), 
	.D(FE_PHN1332_U_afifo_U_acore_n141), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_20_ (.RN(FE_OFN149_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_20_), 
	.D(FE_PHN1330_U_afifo_U_acore_n142), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_19_ (.RN(FE_OFN149_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_19_), 
	.D(FE_PHN1327_U_afifo_U_acore_n144), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_18_ (.RN(FE_OFN35_HRESETn), 
	.Q(U_afifo_U_acore_f_obuf_18_), 
	.D(FE_PHN1265_U_afifo_U_acore_n145), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_17_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_n19), 
	.Q(U_afifo_U_acore_f_obuf_17_), 
	.D(FE_PHN1284_U_afifo_U_acore_n146), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_16_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_n18), 
	.Q(U_afifo_U_acore_f_obuf_16_), 
	.D(FE_PHN1301_U_afifo_U_acore_n147), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_15_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_n17), 
	.Q(U_afifo_U_acore_f_obuf_15_), 
	.D(FE_PHN1313_U_afifo_U_acore_n148), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_14_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n9), 
	.Q(U_afifo_U_acore_f_obuf_14_), 
	.D(FE_PHN1290_U_afifo_U_acore_n149), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_13_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_n16), 
	.Q(U_afifo_U_acore_f_obuf_13_), 
	.D(FE_PHN1276_U_afifo_U_acore_n150), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_12_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_n15), 
	.Q(U_afifo_U_acore_f_obuf_12_), 
	.D(FE_PHN1305_U_afifo_U_acore_n151), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_11_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_n14), 
	.Q(U_afifo_U_acore_f_obuf_11_), 
	.D(FE_PHN1296_U_afifo_U_acore_n152), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_f_obuf_reg_0_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_afifo_U_acore_n3), 
	.Q(U_afifo_U_acore_f_obuf_0_), 
	.D(FE_PHN1282_U_afifo_U_acore_n154), 
	.CK(HCLK__L5_N36));
   DFFS_X2 U_afifo_U_acore_f_obuf_empty_reg (.SN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_n38), 
	.Q(U_afifo_U_acore_n34), 
	.D(FE_PHN3426_U_afifo_U_acore_n_obuf_empty), 
	.CK(HCLK__L5_N38));
   DFFS_X2 U_afifo_U_acore_f_push_req_n_reg (.SN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_n11), 
	.Q(U_afifo_U_acore_f_push_req_n), 
	.D(U_afifo_n55), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_afifo_U_acore_f_ibuf_reg_3_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_U_acore_n33), 
	.D(1'b0), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_f_ibuf_reg_9_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_n32), 
	.D(1'b0), 
	.CK(HCLK__L5_N27));
   DFFR_X1 U_afifo_U_acore_f_ibuf_reg_11_ (.RN(FE_OFN168_HRESETn), 
	.QN(U_afifo_U_acore_n31), 
	.D(U_afifo_m_data_in[11]), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_f_ibuf_reg_45_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_n30), 
	.D(U_afifo_m_data_in[45]), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_f_ibuf_reg_46_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_U_acore_n29), 
	.D(U_afifo_m_data_in[46]), 
	.CK(HCLK__L5_N27));
   DFFR_X1 U_afifo_U_acore_f_ibuf_reg_49_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_n28), 
	.D(FE_PHN1680_U_afifo_m_data_in_49_), 
	.CK(HCLK__L5_N36));
   AOI22_X1 U_dfifo_U_dcore_U224 (.ZN(U_dfifo_U_dcore_n129), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(U_dfifo_m_data_out_0_), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(FE_PHN3246_U_dfifo_U_dcore_f_buf_data_0_));
   AOI22_X1 U_dfifo_U_dcore_U223 (.ZN(U_dfifo_U_dcore_n124), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(U_dfifo_m_data_out_1_), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(FE_PHN1417_U_dfifo_U_dcore_f_buf_data_1_));
   AOI22_X1 U_dfifo_U_dcore_U222 (.ZN(U_dfifo_U_dcore_n122), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(hiu_data[31]), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(U_dfifo_U_dcore_f_buf_data_33_));
   AOI22_X1 U_dfifo_U_dcore_U221 (.ZN(U_dfifo_U_dcore_n120), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(hiu_data[30]), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(U_dfifo_U_dcore_f_buf_data_32_));
   AOI22_X1 U_dfifo_U_dcore_U220 (.ZN(U_dfifo_U_dcore_n118), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(hiu_data[29]), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(FE_PHN3037_U_dfifo_U_dcore_f_buf_data_31_));
   AOI22_X1 U_dfifo_U_dcore_U219 (.ZN(U_dfifo_U_dcore_n116), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(hiu_data[28]), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(FE_PHN3040_U_dfifo_U_dcore_f_buf_data_30_));
   AOI22_X1 U_dfifo_U_dcore_U218 (.ZN(U_dfifo_U_dcore_n114), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(hiu_data[27]), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(U_dfifo_U_dcore_f_buf_data_29_));
   AOI22_X1 U_dfifo_U_dcore_U217 (.ZN(U_dfifo_U_dcore_n112), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(hiu_data[26]), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(FE_PHN3035_U_dfifo_U_dcore_f_buf_data_28_));
   AOI22_X1 U_dfifo_U_dcore_U216 (.ZN(U_dfifo_U_dcore_n110), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(hiu_data[25]), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(U_dfifo_U_dcore_f_buf_data_27_));
   AOI22_X1 U_dfifo_U_dcore_U215 (.ZN(U_dfifo_U_dcore_n108), 
	.B2(U_dfifo_U_dcore_n125), 
	.B1(hiu_data[24]), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(U_dfifo_U_dcore_f_buf_data_26_));
   NAND2_X2 U_dfifo_U_dcore_U213 (.ZN(U_dfifo_U_dcore_n106), 
	.A2(U_dfifo_U_dcore_n125), 
	.A1(U_dfifo_U_dcore_n28));
   NOR2_X4 U_dfifo_U_dcore_U212 (.ZN(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_U_dcore_n209), 
	.A1(U_dfifo_m_empty));
   AND2_X4 U_dfifo_U_dcore_U211 (.ZN(U_dfifo_U_dcore_n2), 
	.A2(U_dfifo_U_dcore_n27), 
	.A1(m_df_push_n));
   NOR4_X4 U_dfifo_U_dcore_U210 (.ZN(U_dfifo_U_dcore_n126), 
	.A4(U_dfifo_U_dcore_n25), 
	.A3(U_dfifo_U_dcore_n26), 
	.A2(U_dfifo_m_aempty), 
	.A1(U_dfifo_m_empty));
   INV_X4 U_dfifo_U_dcore_U209 (.ZN(U_dfifo_U_dcore_n25), 
	.A(U_dfifo_U_dcore_m_sf_empty));
   NOR2_X2 U_dfifo_U_dcore_U208 (.ZN(U_dfifo_m_aempty), 
	.A2(U_dfifo_U_dcore_n25), 
	.A1(U_dfifo_U_dcore_f_buf_has_data));
   AOI21_X2 U_dfifo_U_dcore_U207 (.ZN(U_dfifo_U_dcore_n125), 
	.B2(m_df_push_n), 
	.B1(U_dfifo_m_empty), 
	.A(U_dfifo_n5));
   NAND2_X1 U_dfifo_U_dcore_U206 (.ZN(U_dfifo_U_dcore_n55), 
	.A2(m_two_to_one), 
	.A1(U_dfifo_m_empty));
   NAND2_X2 U_dfifo_U_dcore_U205 (.ZN(U_dfifo_U_dcore_n88), 
	.A2(U_dfifo_U_dcore_n55), 
	.A1(U_dfifo_U_dcore_n125));
   AOI21_X2 U_dfifo_U_dcore_U204 (.ZN(U_dfifo_U_dcore_n59), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[25]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A(U_dfifo_U_dcore_n57));
   AOI21_X2 U_dfifo_U_dcore_U203 (.ZN(U_dfifo_U_dcore_n27), 
	.B2(U_dfifo_m_aempty), 
	.B1(U_dfifo_n5), 
	.A(U_dfifo_m_empty));
   NOR2_X4 U_dfifo_U_dcore_U202 (.ZN(U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_n27), 
	.A1(U_dfifo_U_dcore_n125));
   OAI211_X2 U_dfifo_U_dcore_U201 (.ZN(U_dfifo_U_dcore_n142), 
	.C2(U_dfifo_U_dcore_n88), 
	.C1(FE_PHN3618_U_dfifo_U_dcore_n14), 
	.B(U_dfifo_U_dcore_n58), 
	.A(U_dfifo_U_dcore_n59));
   AOI21_X2 U_dfifo_U_dcore_U200 (.ZN(U_dfifo_U_dcore_n87), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[18]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A(U_dfifo_U_dcore_n85));
   OAI211_X2 U_dfifo_U_dcore_U199 (.ZN(U_dfifo_U_dcore_n149), 
	.C2(U_dfifo_U_dcore_n88), 
	.C1(FE_PHN3632_U_dfifo_U_dcore_n13), 
	.B(U_dfifo_U_dcore_n86), 
	.A(U_dfifo_U_dcore_n87));
   NOR2_X2 U_dfifo_U_dcore_U198 (.ZN(U_dfifo_U_dcore_n103), 
	.A2(U_dfifo_n5), 
	.A1(U_dfifo_m_empty));
   OAI211_X2 U_dfifo_U_dcore_U197 (.ZN(U_dfifo_U_dcore_n150), 
	.C2(U_dfifo_U_dcore_n5), 
	.C1(U_dfifo_U_dcore_n106), 
	.B(U_dfifo_U_dcore_n89), 
	.A(U_dfifo_U_dcore_n90));
   OAI211_X2 U_dfifo_U_dcore_U196 (.ZN(U_dfifo_U_dcore_n157), 
	.C2(U_dfifo_U_dcore_n11), 
	.C1(U_dfifo_U_dcore_n106), 
	.B(U_dfifo_U_dcore_n104), 
	.A(U_dfifo_U_dcore_n105));
   NAND2_X2 U_dfifo_U_dcore_U195 (.ZN(U_dfifo_U_dcore_n21), 
	.A2(U_dfifo_U_dcore_f_buf_has_data), 
	.A1(U_dfifo_U_dcore_m_sf_afull));
   AOI22_X2 U_dfifo_U_dcore_U194 (.ZN(U_dfifo_U_dcore_n53), 
	.B2(m_df_data_in[9]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3114_U_dfifo_U_dcore_f_buf_data_9_), 
	.A1(U_dfifo_U_dcore_n126));
   NAND4_X2 U_dfifo_U_dcore_U193 (.ZN(U_dfifo_U_dcore_n141), 
	.A4(U_dfifo_U_dcore_n56), 
	.A3(U_dfifo_U_dcore_n52), 
	.A2(U_dfifo_U_dcore_n53), 
	.A1(U_dfifo_U_dcore_n54));
   AOI22_X2 U_dfifo_U_dcore_U192 (.ZN(U_dfifo_U_dcore_n30), 
	.B2(FE_OFN255_U_dfifo_U_dcore_n3), 
	.B1(m_df_data_in[2]), 
	.A2(U_dfifo_U_dcore_n126), 
	.A1(FE_PHN3039_U_dfifo_U_dcore_f_buf_data_2_));
   NAND4_X2 U_dfifo_U_dcore_U191 (.ZN(U_dfifo_U_dcore_n134), 
	.A4(U_dfifo_U_dcore_n84), 
	.A3(U_dfifo_U_dcore_n29), 
	.A2(U_dfifo_U_dcore_n30), 
	.A1(U_dfifo_U_dcore_n31));
   AOI21_X2 U_dfifo_U_dcore_U190 (.ZN(U_dfifo_U_dcore_n63), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[24]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A(U_dfifo_U_dcore_n61));
   OAI211_X2 U_dfifo_U_dcore_U189 (.ZN(U_dfifo_U_dcore_n143), 
	.C2(U_dfifo_U_dcore_n88), 
	.C1(U_dfifo_U_dcore_n15), 
	.B(U_dfifo_U_dcore_n62), 
	.A(U_dfifo_U_dcore_n63));
   OAI211_X2 U_dfifo_U_dcore_U188 (.ZN(U_dfifo_U_dcore_n154), 
	.C2(U_dfifo_U_dcore_n8), 
	.C1(U_dfifo_U_dcore_n106), 
	.B(U_dfifo_U_dcore_n97), 
	.A(U_dfifo_U_dcore_n98));
   OAI211_X2 U_dfifo_U_dcore_U187 (.ZN(U_dfifo_U_dcore_n151), 
	.C2(U_dfifo_U_dcore_n6), 
	.C1(U_dfifo_U_dcore_n106), 
	.B(U_dfifo_U_dcore_n91), 
	.A(U_dfifo_U_dcore_n92));
   OAI211_X2 U_dfifo_U_dcore_U186 (.ZN(U_dfifo_U_dcore_n153), 
	.C2(U_dfifo_U_dcore_n7), 
	.C1(U_dfifo_U_dcore_n106), 
	.B(U_dfifo_U_dcore_n95), 
	.A(U_dfifo_U_dcore_n96));
   OAI211_X2 U_dfifo_U_dcore_U185 (.ZN(U_dfifo_U_dcore_n152), 
	.C2(U_dfifo_U_dcore_n12), 
	.C1(U_dfifo_U_dcore_n106), 
	.B(U_dfifo_U_dcore_n93), 
	.A(U_dfifo_U_dcore_n94));
   AOI22_X2 U_dfifo_U_dcore_U184 (.ZN(U_dfifo_U_dcore_n121), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[33]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_df_data_in[33]), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U183 (.ZN(U_dfifo_U_dcore_n165), 
	.A2(U_dfifo_U_dcore_n121), 
	.A1(U_dfifo_U_dcore_n122));
   AOI22_X2 U_dfifo_U_dcore_U182 (.ZN(U_dfifo_U_dcore_n107), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[26]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_df_data_in[26]), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U181 (.ZN(U_dfifo_U_dcore_n158), 
	.A2(U_dfifo_U_dcore_n107), 
	.A1(U_dfifo_U_dcore_n108));
   AOI21_X2 U_dfifo_U_dcore_U180 (.ZN(U_dfifo_U_dcore_n67), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[23]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A(U_dfifo_U_dcore_n65));
   OAI211_X2 U_dfifo_U_dcore_U179 (.ZN(U_dfifo_U_dcore_n144), 
	.C2(U_dfifo_U_dcore_n88), 
	.C1(U_dfifo_U_dcore_n16), 
	.B(U_dfifo_U_dcore_n66), 
	.A(U_dfifo_U_dcore_n67));
   OAI211_X2 U_dfifo_U_dcore_U178 (.ZN(U_dfifo_U_dcore_n156), 
	.C2(U_dfifo_U_dcore_n10), 
	.C1(U_dfifo_U_dcore_n106), 
	.B(U_dfifo_U_dcore_n101), 
	.A(U_dfifo_U_dcore_n102));
   OAI211_X2 U_dfifo_U_dcore_U177 (.ZN(U_dfifo_U_dcore_n155), 
	.C2(U_dfifo_U_dcore_n9), 
	.C1(U_dfifo_U_dcore_n106), 
	.B(U_dfifo_U_dcore_n99), 
	.A(U_dfifo_U_dcore_n100));
   OAI22_X2 U_dfifo_U_dcore_U176 (.ZN(U_dfifo_U_dcore_n234), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_33_), 
	.A2(m_df_data_in[33]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U175 (.ZN(U_dfifo_U_dcore_n201), 
	.A(U_dfifo_U_dcore_n234));
   OAI22_X2 U_dfifo_U_dcore_U174 (.ZN(U_dfifo_U_dcore_n227), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_26_), 
	.A2(m_df_data_in[26]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U173 (.ZN(U_dfifo_U_dcore_n194), 
	.A(U_dfifo_U_dcore_n227));
   OAI22_X2 U_dfifo_U_dcore_U172 (.ZN(U_dfifo_U_dcore_n219), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_18_), 
	.A2(m_df_data_in[18]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U171 (.ZN(U_dfifo_U_dcore_n186), 
	.A(U_dfifo_U_dcore_n219));
   OAI22_X2 U_dfifo_U_dcore_U170 (.ZN(U_dfifo_U_dcore_n226), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_25_), 
	.A2(m_df_data_in[25]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U169 (.ZN(U_dfifo_U_dcore_n193), 
	.A(U_dfifo_U_dcore_n226));
   AOI21_X2 U_dfifo_U_dcore_U168 (.ZN(U_dfifo_U_dcore_n79), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[20]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A(U_dfifo_U_dcore_n77));
   OAI211_X2 U_dfifo_U_dcore_U167 (.ZN(U_dfifo_U_dcore_n147), 
	.C2(U_dfifo_U_dcore_n88), 
	.C1(U_dfifo_U_dcore_n19), 
	.B(U_dfifo_U_dcore_n78), 
	.A(U_dfifo_U_dcore_n79));
   AOI21_X2 U_dfifo_U_dcore_U166 (.ZN(U_dfifo_U_dcore_n83), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[19]), 
	.B1(FE_OFN252_U_dfifo_U_dcore_n127), 
	.A(U_dfifo_U_dcore_n81));
   OAI211_X2 U_dfifo_U_dcore_U165 (.ZN(U_dfifo_U_dcore_n148), 
	.C2(U_dfifo_U_dcore_n88), 
	.C1(U_dfifo_U_dcore_n20), 
	.B(U_dfifo_U_dcore_n82), 
	.A(U_dfifo_U_dcore_n83));
   AOI21_X2 U_dfifo_U_dcore_U164 (.ZN(U_dfifo_U_dcore_n71), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[22]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A(U_dfifo_U_dcore_n69));
   OAI211_X2 U_dfifo_U_dcore_U163 (.ZN(U_dfifo_U_dcore_n145), 
	.C2(U_dfifo_U_dcore_n88), 
	.C1(U_dfifo_U_dcore_n17), 
	.B(U_dfifo_U_dcore_n70), 
	.A(U_dfifo_U_dcore_n71));
   AOI21_X2 U_dfifo_U_dcore_U162 (.ZN(U_dfifo_U_dcore_n75), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[21]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A(U_dfifo_U_dcore_n73));
   OAI211_X2 U_dfifo_U_dcore_U161 (.ZN(U_dfifo_U_dcore_n146), 
	.C2(U_dfifo_U_dcore_n88), 
	.C1(U_dfifo_U_dcore_n18), 
	.B(U_dfifo_U_dcore_n74), 
	.A(U_dfifo_U_dcore_n75));
   NAND4_X2 U_dfifo_U_dcore_U160 (.ZN(U_dfifo_U_dcore_n140), 
	.A4(U_dfifo_U_dcore_n60), 
	.A3(U_dfifo_U_dcore_n47), 
	.A2(U_dfifo_U_dcore_n48), 
	.A1(U_dfifo_U_dcore_n49));
   OAI221_X2 U_dfifo_U_dcore_U159 (.ZN(U_dfifo_U_dcore_n208), 
	.C2(U_dfifo_U_dcore_n25), 
	.C1(U_dfifo_U_dcore_n26), 
	.B2(U_dfifo_U_dcore_n24), 
	.B1(U_dfifo_n5), 
	.A(U_dfifo_U_dcore_f_buf_has_data));
   NAND4_X2 U_dfifo_U_dcore_U158 (.ZN(U_dfifo_U_dcore_n137), 
	.A4(U_dfifo_U_dcore_n72), 
	.A3(U_dfifo_U_dcore_n38), 
	.A2(U_dfifo_U_dcore_n39), 
	.A1(U_dfifo_U_dcore_n40));
   NAND4_X2 U_dfifo_U_dcore_U157 (.ZN(U_dfifo_U_dcore_n136), 
	.A4(U_dfifo_U_dcore_n76), 
	.A3(U_dfifo_U_dcore_n35), 
	.A2(U_dfifo_U_dcore_n36), 
	.A1(U_dfifo_U_dcore_n37));
   NAND4_X2 U_dfifo_U_dcore_U156 (.ZN(U_dfifo_U_dcore_n139), 
	.A4(U_dfifo_U_dcore_n64), 
	.A3(U_dfifo_U_dcore_n44), 
	.A2(U_dfifo_U_dcore_n45), 
	.A1(U_dfifo_U_dcore_n46));
   NAND4_X2 U_dfifo_U_dcore_U155 (.ZN(U_dfifo_U_dcore_n138), 
	.A4(U_dfifo_U_dcore_n68), 
	.A3(U_dfifo_U_dcore_n41), 
	.A2(U_dfifo_U_dcore_n42), 
	.A1(U_dfifo_U_dcore_n43));
   NAND4_X2 U_dfifo_U_dcore_U154 (.ZN(U_dfifo_U_dcore_n135), 
	.A4(U_dfifo_U_dcore_n80), 
	.A3(U_dfifo_U_dcore_n32), 
	.A2(U_dfifo_U_dcore_n33), 
	.A1(U_dfifo_U_dcore_n34));
   OAI22_X2 U_dfifo_U_dcore_U153 (.ZN(U_dfifo_U_dcore_n132), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3039_U_dfifo_U_dcore_f_buf_data_2_), 
	.A2(m_df_data_in[2]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U152 (.ZN(U_dfifo_U_dcore_n170), 
	.A(U_dfifo_U_dcore_n132));
   OAI22_X2 U_dfifo_U_dcore_U151 (.ZN(U_dfifo_U_dcore_n218), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3117_U_dfifo_U_dcore_f_buf_data_17_), 
	.A2(m_df_data_in[17]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U150 (.ZN(U_dfifo_U_dcore_n185), 
	.A(U_dfifo_U_dcore_n218));
   OAI22_X2 U_dfifo_U_dcore_U149 (.ZN(U_dfifo_U_dcore_n210), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3114_U_dfifo_U_dcore_f_buf_data_9_), 
	.A2(m_df_data_in[9]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U148 (.ZN(U_dfifo_U_dcore_n177), 
	.A(U_dfifo_U_dcore_n210));
   OAI22_X2 U_dfifo_U_dcore_U147 (.ZN(U_dfifo_U_dcore_n211), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_10_), 
	.A2(m_df_data_in[10]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U146 (.ZN(U_dfifo_U_dcore_n178), 
	.A(U_dfifo_U_dcore_n211));
   AOI22_X2 U_dfifo_U_dcore_U145 (.ZN(U_dfifo_U_dcore_n117), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[31]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_df_data_in[31]), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U144 (.ZN(U_dfifo_U_dcore_n163), 
	.A2(U_dfifo_U_dcore_n117), 
	.A1(U_dfifo_U_dcore_n118));
   AOI22_X2 U_dfifo_U_dcore_U143 (.ZN(U_dfifo_U_dcore_n119), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[32]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_df_data_in[32]), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U142 (.ZN(U_dfifo_U_dcore_n164), 
	.A2(U_dfifo_U_dcore_n119), 
	.A1(U_dfifo_U_dcore_n120));
   AOI22_X2 U_dfifo_U_dcore_U141 (.ZN(U_dfifo_U_dcore_n128), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[0]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_df_data_in[0]), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U140 (.ZN(U_dfifo_U_dcore_n167), 
	.A2(U_dfifo_U_dcore_n128), 
	.A1(U_dfifo_U_dcore_n129));
   OAI22_X2 U_dfifo_U_dcore_U139 (.ZN(U_dfifo_U_dcore_n225), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_24_), 
	.A2(m_df_data_in[24]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U138 (.ZN(U_dfifo_U_dcore_n192), 
	.A(U_dfifo_U_dcore_n225));
   OAI22_X2 U_dfifo_U_dcore_U137 (.ZN(U_dfifo_U_dcore_n232), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3037_U_dfifo_U_dcore_f_buf_data_31_), 
	.A2(m_df_data_in[31]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U136 (.ZN(U_dfifo_U_dcore_n199), 
	.A(U_dfifo_U_dcore_n232));
   OAI22_X2 U_dfifo_U_dcore_U135 (.ZN(U_dfifo_U_dcore_n233), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_32_), 
	.A2(m_df_data_in[32]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U134 (.ZN(U_dfifo_U_dcore_n200), 
	.A(U_dfifo_U_dcore_n233));
   AOI22_X2 U_dfifo_U_dcore_U133 (.ZN(U_dfifo_U_dcore_n111), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[28]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_df_data_in[28]), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U132 (.ZN(U_dfifo_U_dcore_n160), 
	.A2(U_dfifo_U_dcore_n111), 
	.A1(U_dfifo_U_dcore_n112));
   AOI22_X2 U_dfifo_U_dcore_U131 (.ZN(U_dfifo_U_dcore_n109), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[27]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_df_data_in[27]), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U130 (.ZN(U_dfifo_U_dcore_n159), 
	.A2(U_dfifo_U_dcore_n109), 
	.A1(U_dfifo_U_dcore_n110));
   AOI22_X2 U_dfifo_U_dcore_U129 (.ZN(U_dfifo_U_dcore_n113), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[29]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_df_data_in[29]), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U128 (.ZN(U_dfifo_U_dcore_n161), 
	.A2(U_dfifo_U_dcore_n113), 
	.A1(U_dfifo_U_dcore_n114));
   AOI22_X2 U_dfifo_U_dcore_U127 (.ZN(U_dfifo_U_dcore_n115), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[30]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_df_data_in[30]), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U126 (.ZN(U_dfifo_U_dcore_n162), 
	.A2(U_dfifo_U_dcore_n115), 
	.A1(U_dfifo_U_dcore_n116));
   OAI22_X2 U_dfifo_U_dcore_U125 (.ZN(U_dfifo_U_dcore_n216), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3118_U_dfifo_U_dcore_f_buf_data_15_), 
	.A2(m_df_data_in[15]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U124 (.ZN(U_dfifo_U_dcore_n183), 
	.A(U_dfifo_U_dcore_n216));
   OAI22_X2 U_dfifo_U_dcore_U123 (.ZN(U_dfifo_U_dcore_n217), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_16_), 
	.A2(m_df_data_in[16]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U122 (.ZN(U_dfifo_U_dcore_n184), 
	.A(U_dfifo_U_dcore_n217));
   OAI22_X2 U_dfifo_U_dcore_U121 (.ZN(U_dfifo_U_dcore_n207), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_8_), 
	.A2(m_df_data_in[8]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U120 (.ZN(U_dfifo_U_dcore_n176), 
	.A(U_dfifo_U_dcore_n207));
   OAI22_X2 U_dfifo_U_dcore_U119 (.ZN(U_dfifo_U_dcore_n212), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_11_), 
	.A2(m_df_data_in[11]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U118 (.ZN(U_dfifo_U_dcore_n179), 
	.A(U_dfifo_U_dcore_n212));
   OAI22_X2 U_dfifo_U_dcore_U117 (.ZN(U_dfifo_U_dcore_n214), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_13_), 
	.A2(m_df_data_in[13]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U116 (.ZN(U_dfifo_U_dcore_n181), 
	.A(U_dfifo_U_dcore_n214));
   OAI22_X2 U_dfifo_U_dcore_U115 (.ZN(U_dfifo_U_dcore_n213), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_12_), 
	.A2(m_df_data_in[12]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U114 (.ZN(U_dfifo_U_dcore_n180), 
	.A(U_dfifo_U_dcore_n213));
   OAI22_X2 U_dfifo_U_dcore_U113 (.ZN(U_dfifo_U_dcore_n215), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_14_), 
	.A2(m_df_data_in[14]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U112 (.ZN(U_dfifo_U_dcore_n182), 
	.A(U_dfifo_U_dcore_n215));
   OAI22_X2 U_dfifo_U_dcore_U111 (.ZN(U_dfifo_U_dcore_n224), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_23_), 
	.A2(m_df_data_in[23]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U110 (.ZN(U_dfifo_U_dcore_n191), 
	.A(U_dfifo_U_dcore_n224));
   OAI22_X2 U_dfifo_U_dcore_U109 (.ZN(U_dfifo_U_dcore_n220), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3122_U_dfifo_U_dcore_f_buf_data_19_), 
	.A2(m_df_data_in[19]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U108 (.ZN(U_dfifo_U_dcore_n187), 
	.A(U_dfifo_U_dcore_n220));
   OAI22_X2 U_dfifo_U_dcore_U107 (.ZN(U_dfifo_U_dcore_n221), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_20_), 
	.A2(m_df_data_in[20]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U106 (.ZN(U_dfifo_U_dcore_n188), 
	.A(U_dfifo_U_dcore_n221));
   OAI22_X2 U_dfifo_U_dcore_U105 (.ZN(U_dfifo_U_dcore_n222), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_21_), 
	.A2(m_df_data_in[21]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U104 (.ZN(U_dfifo_U_dcore_n189), 
	.A(U_dfifo_U_dcore_n222));
   OAI22_X2 U_dfifo_U_dcore_U103 (.ZN(U_dfifo_U_dcore_n223), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3116_U_dfifo_U_dcore_f_buf_data_22_), 
	.A2(m_df_data_in[22]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U102 (.ZN(U_dfifo_U_dcore_n190), 
	.A(U_dfifo_U_dcore_n223));
   OAI22_X2 U_dfifo_U_dcore_U101 (.ZN(U_dfifo_U_dcore_n130), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3246_U_dfifo_U_dcore_f_buf_data_0_), 
	.A2(m_df_data_in[0]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U100 (.ZN(U_dfifo_U_dcore_n168), 
	.A(U_dfifo_U_dcore_n130));
   OAI22_X2 U_dfifo_U_dcore_U99 (.ZN(U_dfifo_U_dcore_n206), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3121_U_dfifo_U_dcore_f_buf_data_7_), 
	.A2(m_df_data_in[7]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U98 (.ZN(U_dfifo_U_dcore_n175), 
	.A(U_dfifo_U_dcore_n206));
   OAI22_X2 U_dfifo_U_dcore_U97 (.ZN(U_dfifo_U_dcore_n205), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3124_U_dfifo_U_dcore_f_buf_data_6_), 
	.A2(m_df_data_in[6]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U96 (.ZN(U_dfifo_U_dcore_n174), 
	.A(U_dfifo_U_dcore_n205));
   OAI22_X2 U_dfifo_U_dcore_U95 (.ZN(U_dfifo_U_dcore_n133), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3120_U_dfifo_U_dcore_f_buf_data_3_), 
	.A2(m_df_data_in[3]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U94 (.ZN(U_dfifo_U_dcore_n171), 
	.A(U_dfifo_U_dcore_n133));
   OAI22_X2 U_dfifo_U_dcore_U93 (.ZN(U_dfifo_U_dcore_n202), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3036_U_dfifo_U_dcore_f_buf_data_4_), 
	.A2(m_df_data_in[4]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U92 (.ZN(U_dfifo_U_dcore_n172), 
	.A(U_dfifo_U_dcore_n202));
   OAI22_X2 U_dfifo_U_dcore_U91 (.ZN(U_dfifo_U_dcore_n204), 
	.B2(FE_OFN256_U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3038_U_dfifo_U_dcore_f_buf_data_5_), 
	.A2(m_df_data_in[5]), 
	.A1(U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U90 (.ZN(U_dfifo_U_dcore_n173), 
	.A(U_dfifo_U_dcore_n204));
   OAI22_X2 U_dfifo_U_dcore_U89 (.ZN(U_dfifo_U_dcore_n228), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_27_), 
	.A2(m_df_data_in[27]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U88 (.ZN(U_dfifo_U_dcore_n195), 
	.A(U_dfifo_U_dcore_n228));
   OAI22_X2 U_dfifo_U_dcore_U87 (.ZN(U_dfifo_U_dcore_n230), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(U_dfifo_U_dcore_f_buf_data_29_), 
	.A2(m_df_data_in[29]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U86 (.ZN(U_dfifo_U_dcore_n197), 
	.A(U_dfifo_U_dcore_n230));
   OAI22_X2 U_dfifo_U_dcore_U85 (.ZN(U_dfifo_U_dcore_n229), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3035_U_dfifo_U_dcore_f_buf_data_28_), 
	.A2(m_df_data_in[28]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U84 (.ZN(U_dfifo_U_dcore_n196), 
	.A(U_dfifo_U_dcore_n229));
   OAI22_X2 U_dfifo_U_dcore_U83 (.ZN(U_dfifo_U_dcore_n231), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(FE_PHN3040_U_dfifo_U_dcore_f_buf_data_30_), 
	.A2(m_df_data_in[30]), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U82 (.ZN(U_dfifo_U_dcore_n198), 
	.A(U_dfifo_U_dcore_n231));
   NAND2_X2 U_dfifo_U_dcore_U81 (.ZN(U_dfifo_U_dcore_n166), 
	.A2(U_dfifo_U_dcore_n123), 
	.A1(U_dfifo_U_dcore_n124));
   OAI22_X2 U_dfifo_U_dcore_U80 (.ZN(U_dfifo_U_dcore_n131), 
	.B2(U_dfifo_U_dcore_n2), 
	.B1(FE_PHN1417_U_dfifo_U_dcore_f_buf_data_1_), 
	.A2(m_double), 
	.A1(FE_OFN258_U_dfifo_U_dcore_n1));
   INV_X4 U_dfifo_U_dcore_U79 (.ZN(U_dfifo_U_dcore_n169), 
	.A(U_dfifo_U_dcore_n131));
   OAI21_X1 U_dfifo_U_dcore_U78 (.ZN(U_dfifo_U_dcore_n203), 
	.B2(U_dfifo_U_dcore_n23), 
	.B1(U_dfifo_n5), 
	.A(FE_OFN258_U_dfifo_U_dcore_n1));
   AOI22_X2 U_dfifo_U_dcore_U77 (.ZN(U_dfifo_U_dcore_n48), 
	.B2(m_df_data_in[8]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_8_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U76 (.ZN(U_dfifo_U_dcore_n39), 
	.B2(m_df_data_in[5]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3038_U_dfifo_U_dcore_f_buf_data_5_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U75 (.ZN(U_dfifo_U_dcore_n36), 
	.B2(m_df_data_in[4]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3036_U_dfifo_U_dcore_f_buf_data_4_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U74 (.ZN(U_dfifo_U_dcore_n45), 
	.B2(m_df_data_in[7]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3121_U_dfifo_U_dcore_f_buf_data_7_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U73 (.ZN(U_dfifo_U_dcore_n42), 
	.B2(m_df_data_in[6]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3124_U_dfifo_U_dcore_f_buf_data_6_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U72 (.ZN(U_dfifo_U_dcore_n33), 
	.B2(m_df_data_in[3]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3120_U_dfifo_U_dcore_f_buf_data_3_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U71 (.ZN(U_dfifo_U_dcore_n89), 
	.B2(m_df_data_in[10]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_10_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U70 (.ZN(U_dfifo_U_dcore_n104), 
	.B2(m_df_data_in[17]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3117_U_dfifo_U_dcore_f_buf_data_17_), 
	.A1(U_dfifo_U_dcore_n126));
   NOR3_X1 U_dfifo_U_dcore_U69 (.ZN(U_dfifo_U_dcore_n51), 
	.A3(U_dfifo_U_dcore_n55), 
	.A2(m_df_push_n), 
	.A1(U_dfifo_n5));
   AOI22_X2 U_dfifo_U_dcore_U68 (.ZN(U_dfifo_U_dcore_n58), 
	.B2(m_df_data_in[25]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_25_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U67 (.ZN(U_dfifo_U_dcore_n86), 
	.B2(m_df_data_in[18]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_18_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U66 (.ZN(U_dfifo_U_dcore_n62), 
	.B2(m_df_data_in[24]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_24_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U65 (.ZN(U_dfifo_U_dcore_n97), 
	.B2(m_df_data_in[14]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_14_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U64 (.ZN(U_dfifo_U_dcore_n91), 
	.B2(m_df_data_in[11]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_11_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U63 (.ZN(U_dfifo_U_dcore_n95), 
	.B2(m_df_data_in[13]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_13_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U62 (.ZN(U_dfifo_U_dcore_n93), 
	.B2(m_df_data_in[12]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_12_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U61 (.ZN(U_dfifo_U_dcore_n66), 
	.B2(m_df_data_in[23]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_23_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U60 (.ZN(U_dfifo_U_dcore_n101), 
	.B2(m_df_data_in[16]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_16_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U59 (.ZN(U_dfifo_U_dcore_n99), 
	.B2(m_df_data_in[15]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3118_U_dfifo_U_dcore_f_buf_data_15_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U58 (.ZN(U_dfifo_U_dcore_n78), 
	.B2(m_df_data_in[20]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_20_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U57 (.ZN(U_dfifo_U_dcore_n82), 
	.B2(m_df_data_in[19]), 
	.B1(FE_OFN255_U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3122_U_dfifo_U_dcore_f_buf_data_19_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U56 (.ZN(U_dfifo_U_dcore_n70), 
	.B2(m_df_data_in[22]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(FE_PHN3116_U_dfifo_U_dcore_f_buf_data_22_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U55 (.ZN(U_dfifo_U_dcore_n74), 
	.B2(m_df_data_in[21]), 
	.B1(U_dfifo_U_dcore_n3), 
	.A2(U_dfifo_U_dcore_f_buf_data_21_), 
	.A1(U_dfifo_U_dcore_n126));
   AOI22_X2 U_dfifo_U_dcore_U54 (.ZN(U_dfifo_U_dcore_n123), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[1]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(m_double), 
	.A1(U_dfifo_U_dcore_n3));
   NAND2_X2 U_dfifo_U_dcore_U53 (.ZN(U_dfifo_U_dcore_n209), 
	.A2(U_dfifo_U_dcore_n25), 
	.A1(U_dfifo_n5));
   NOR2_X1 U_dfifo_U_dcore_U52 (.ZN(U_dfifo_U_dcore_n50), 
	.A2(U_dfifo_U_dcore_n106), 
	.A1(m_two_to_one));
   NAND2_X1 U_dfifo_U_dcore_U51 (.ZN(U_dfifo_U_dcore_n22), 
	.A2(U_dfifo_U_dcore_n4), 
	.A1(FE_PHN1423_U_dfifo_U_dcore_m_sf_full));
   INV_X2 U_dfifo_U_dcore_U50 (.ZN(U_dfifo_U_dcore_n24), 
	.A(FE_PHN1423_U_dfifo_U_dcore_m_sf_full));
   INV_X2 U_dfifo_U_dcore_U49 (.ZN(U_dfifo_U_dcore_n26), 
	.A(U_dfifo_n5));
   NAND2_X1 U_dfifo_U_dcore_U48 (.ZN(U_dfifo_U_dcore_n76), 
	.A2(FE_OFN225_hiu_data_26_), 
	.A1(U_dfifo_U_dcore_n51));
   NOR2_X1 U_dfifo_U_dcore_U47 (.ZN(U_dfifo_U_dcore_n_empty), 
	.A2(U_dfifo_U_dcore_n27), 
	.A1(m_df_push_n));
   NAND2_X1 U_dfifo_U_dcore_U46 (.ZN(U_dfifo_U_dcore_n56), 
	.A2(hiu_data[31]), 
	.A1(U_dfifo_U_dcore_n51));
   NAND2_X1 U_dfifo_U_dcore_U45 (.ZN(U_dfifo_U_dcore_n80), 
	.A2(hiu_data[25]), 
	.A1(U_dfifo_U_dcore_n51));
   NAND2_X1 U_dfifo_U_dcore_U44 (.ZN(U_dfifo_U_dcore_n60), 
	.A2(hiu_data[30]), 
	.A1(U_dfifo_U_dcore_n51));
   NAND2_X1 U_dfifo_U_dcore_U43 (.ZN(U_dfifo_U_dcore_n64), 
	.A2(hiu_data[29]), 
	.A1(U_dfifo_U_dcore_n51));
   NAND2_X1 U_dfifo_U_dcore_U42 (.ZN(U_dfifo_U_dcore_n72), 
	.A2(hiu_data[27]), 
	.A1(U_dfifo_U_dcore_n51));
   NAND2_X1 U_dfifo_U_dcore_U41 (.ZN(U_dfifo_U_dcore_n68), 
	.A2(hiu_data[28]), 
	.A1(U_dfifo_U_dcore_n51));
   NAND2_X1 U_dfifo_U_dcore_U40 (.ZN(U_dfifo_U_dcore_n84), 
	.A2(U_dfifo_U_dcore_n51), 
	.A1(hiu_data[24]));
   INV_X2 U_dfifo_U_dcore_U39 (.ZN(U_dfifo_U_dcore_n57), 
	.A(U_dfifo_U_dcore_n56));
   AOI22_X1 U_dfifo_U_dcore_U38 (.ZN(U_dfifo_U_dcore_n34), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[3]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[1]), 
	.A1(U_dfifo_U_dcore_n103));
   INV_X2 U_dfifo_U_dcore_U37 (.ZN(U_dfifo_U_dcore_n73), 
	.A(U_dfifo_U_dcore_n72));
   AOI22_X1 U_dfifo_U_dcore_U36 (.ZN(U_dfifo_U_dcore_n31), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[2]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[0]), 
	.A1(U_dfifo_U_dcore_n103));
   INV_X2 U_dfifo_U_dcore_U35 (.ZN(U_dfifo_U_dcore_n69), 
	.A(U_dfifo_U_dcore_n68));
   AOI22_X1 U_dfifo_U_dcore_U34 (.ZN(U_dfifo_U_dcore_n92), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[11]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[9]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U33 (.ZN(U_dfifo_U_dcore_n54), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[9]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[7]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U32 (.ZN(U_dfifo_U_dcore_n94), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[12]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[10]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U31 (.ZN(U_dfifo_U_dcore_n90), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[10]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[8]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U30 (.ZN(U_dfifo_U_dcore_n49), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[8]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[6]), 
	.A1(U_dfifo_U_dcore_n103));
   INV_X2 U_dfifo_U_dcore_U29 (.ZN(U_dfifo_U_dcore_n85), 
	.A(U_dfifo_U_dcore_n84));
   AOI22_X1 U_dfifo_U_dcore_U28 (.ZN(U_dfifo_U_dcore_n96), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[13]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[11]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U27 (.ZN(U_dfifo_U_dcore_n46), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[7]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[5]), 
	.A1(U_dfifo_U_dcore_n103));
   INV_X2 U_dfifo_U_dcore_U26 (.ZN(U_dfifo_U_dcore_n61), 
	.A(U_dfifo_U_dcore_n60));
   INV_X2 U_dfifo_U_dcore_U25 (.ZN(U_dfifo_U_dcore_n81), 
	.A(U_dfifo_U_dcore_n80));
   AOI22_X1 U_dfifo_U_dcore_U24 (.ZN(U_dfifo_U_dcore_n98), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[14]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[12]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U23 (.ZN(U_dfifo_U_dcore_n37), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[4]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[2]), 
	.A1(U_dfifo_U_dcore_n103));
   INV_X2 U_dfifo_U_dcore_U22 (.ZN(U_dfifo_U_dcore_n77), 
	.A(U_dfifo_U_dcore_n76));
   AOI22_X1 U_dfifo_U_dcore_U21 (.ZN(U_dfifo_U_dcore_n43), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[6]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[4]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U20 (.ZN(U_dfifo_U_dcore_n105), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[17]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[15]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U19 (.ZN(U_dfifo_U_dcore_n100), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[15]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[13]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U18 (.ZN(U_dfifo_U_dcore_n102), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[16]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[14]), 
	.A1(U_dfifo_U_dcore_n103));
   AOI22_X1 U_dfifo_U_dcore_U17 (.ZN(U_dfifo_U_dcore_n40), 
	.B2(U_dfifo_U_dcore_m_sf_data_out[5]), 
	.B1(U_dfifo_U_dcore_n127), 
	.A2(U_dfifo_m_btm_data[3]), 
	.A1(U_dfifo_U_dcore_n103));
   INV_X2 U_dfifo_U_dcore_U16 (.ZN(U_dfifo_U_dcore_n65), 
	.A(U_dfifo_U_dcore_n64));
   NAND2_X1 U_dfifo_U_dcore_U15 (.ZN(U_dfifo_U_dcore_n44), 
	.A2(hiu_data[21]), 
	.A1(U_dfifo_U_dcore_n50));
   NAND2_X1 U_dfifo_U_dcore_U14 (.ZN(U_dfifo_U_dcore_n32), 
	.A2(hiu_data[17]), 
	.A1(U_dfifo_U_dcore_n50));
   NAND2_X1 U_dfifo_U_dcore_U13 (.ZN(U_dfifo_U_dcore_n41), 
	.A2(hiu_data[20]), 
	.A1(U_dfifo_U_dcore_n50));
   NAND2_X1 U_dfifo_U_dcore_U12 (.ZN(U_dfifo_U_dcore_n38), 
	.A2(hiu_data[19]), 
	.A1(U_dfifo_U_dcore_n50));
   NAND2_X1 U_dfifo_U_dcore_U11 (.ZN(U_dfifo_U_dcore_n52), 
	.A2(hiu_data[23]), 
	.A1(U_dfifo_U_dcore_n50));
   NAND2_X1 U_dfifo_U_dcore_U10 (.ZN(U_dfifo_U_dcore_n29), 
	.A2(U_dfifo_U_dcore_n50), 
	.A1(hiu_data[16]));
   NAND2_X1 U_dfifo_U_dcore_U9 (.ZN(U_dfifo_U_dcore_n47), 
	.A2(hiu_data[22]), 
	.A1(U_dfifo_U_dcore_n50));
   NAND2_X1 U_dfifo_U_dcore_U8 (.ZN(U_dfifo_U_dcore_n35), 
	.A2(hiu_data[18]), 
	.A1(U_dfifo_U_dcore_n50));
   INV_X2 U_dfifo_U_dcore_U7 (.ZN(U_dfifo_U_dcore_n28), 
	.A(U_dfifo_U_dcore_n103));
   INV_X4 U_dfifo_U_dcore_U6 (.ZN(U_dfifo_U_dcore_n1), 
	.A(U_dfifo_U_dcore_n2));
   NAND2_X1 U_dfifo_U_dcore_U5 (.ZN(U_dfifo_m_afull), 
	.A2(U_dfifo_U_dcore_n22), 
	.A1(U_dfifo_U_dcore_n21));
   INV_X4 U_dfifo_U_dcore_U4 (.ZN(U_dfifo_m_full), 
	.A(U_dfifo_U_dcore_n23));
   NAND2_X2 U_dfifo_U_dcore_U3 (.ZN(U_dfifo_U_dcore_n23), 
	.A2(U_dfifo_U_dcore_f_buf_has_data), 
	.A1(FE_PHN1423_U_dfifo_U_dcore_m_sf_full));
   DFFR_X2 U_dfifo_U_dcore_f_data_out_reg_18_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_dfifo_U_dcore_n13), 
	.Q(hiu_data[16]), 
	.D(FE_PHN1181_U_dfifo_U_dcore_n149), 
	.CK(HCLK__L5_N18));
   DFFR_X2 U_dfifo_U_dcore_f_data_out_reg_25_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_dfifo_U_dcore_n14), 
	.Q(hiu_data[23]), 
	.D(FE_PHN1179_U_dfifo_U_dcore_n142), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_2_ (.RN(FE_OFN53_HRESETn), 
	.Q(U_dfifo_m_btm_data[0]), 
	.D(FE_PHN1018_U_dfifo_U_dcore_n134), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_3_ (.RN(FE_OFN53_HRESETn), 
	.Q(U_dfifo_m_btm_data[1]), 
	.D(FE_PHN857_U_dfifo_U_dcore_n135), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_4_ (.RN(FE_OFN53_HRESETn), 
	.Q(U_dfifo_m_btm_data[2]), 
	.D(FE_PHN785_U_dfifo_U_dcore_n136), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_5_ (.RN(FE_OFN28_HRESETn), 
	.Q(U_dfifo_m_btm_data[3]), 
	.D(FE_PHN1022_U_dfifo_U_dcore_n137), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_6_ (.RN(FE_OFN28_HRESETn), 
	.Q(U_dfifo_m_btm_data[4]), 
	.D(FE_PHN1021_U_dfifo_U_dcore_n138), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_7_ (.RN(FE_OFN53_HRESETn), 
	.Q(U_dfifo_m_btm_data[5]), 
	.D(FE_PHN784_U_dfifo_U_dcore_n139), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_8_ (.RN(FE_OFN53_HRESETn), 
	.Q(U_dfifo_m_btm_data[6]), 
	.D(FE_PHN858_U_dfifo_U_dcore_n140), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_9_ (.RN(FE_OFN53_HRESETn), 
	.Q(U_dfifo_m_btm_data[7]), 
	.D(FE_PHN1019_U_dfifo_U_dcore_n141), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_24_ (.RN(FE_OFN28_HRESETn), 
	.QN(U_dfifo_U_dcore_n15), 
	.Q(hiu_data[22]), 
	.D(FE_PHN1182_U_dfifo_U_dcore_n143), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_23_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_dfifo_U_dcore_n16), 
	.Q(hiu_data[21]), 
	.D(FE_PHN861_U_dfifo_U_dcore_n144), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_22_ (.RN(FE_OFN160_HRESETn), 
	.QN(U_dfifo_U_dcore_n17), 
	.Q(hiu_data[20]), 
	.D(FE_PHN1630_U_dfifo_U_dcore_n145), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_21_ (.RN(FE_OFN196_HRESETn), 
	.QN(U_dfifo_U_dcore_n18), 
	.Q(hiu_data[19]), 
	.D(FE_PHN1180_U_dfifo_U_dcore_n146), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_20_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_dfifo_U_dcore_n19), 
	.Q(hiu_data[18]), 
	.D(FE_PHN956_U_dfifo_U_dcore_n147), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_19_ (.RN(FE_OFN28_HRESETn), 
	.QN(U_dfifo_U_dcore_n20), 
	.Q(hiu_data[17]), 
	.D(FE_PHN860_U_dfifo_U_dcore_n148), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_10_ (.RN(FE_OFN196_HRESETn), 
	.Q(U_dfifo_m_btm_data[8]), 
	.D(FE_PHN954_U_dfifo_U_dcore_n150), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_11_ (.RN(FE_OFN160_HRESETn), 
	.Q(U_dfifo_m_btm_data[9]), 
	.D(FE_PHN812_U_dfifo_U_dcore_n151), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_12_ (.RN(FE_OFN196_HRESETn), 
	.Q(U_dfifo_m_btm_data[10]), 
	.D(FE_PHN909_U_dfifo_U_dcore_n152), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_13_ (.RN(FE_OFN196_HRESETn), 
	.Q(U_dfifo_m_btm_data[11]), 
	.D(FE_PHN910_U_dfifo_U_dcore_n153), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_14_ (.RN(FE_OFN196_HRESETn), 
	.Q(U_dfifo_m_btm_data[12]), 
	.D(FE_PHN1084_U_dfifo_U_dcore_n154), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_15_ (.RN(FE_OFN196_HRESETn), 
	.Q(U_dfifo_m_btm_data[13]), 
	.D(FE_PHN810_U_dfifo_U_dcore_n155), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_16_ (.RN(FE_OFN196_HRESETn), 
	.Q(U_dfifo_m_btm_data[14]), 
	.D(FE_PHN811_U_dfifo_U_dcore_n156), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_17_ (.RN(FE_OFN53_HRESETn), 
	.Q(U_dfifo_m_btm_data[15]), 
	.D(FE_PHN809_U_dfifo_U_dcore_n157), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_26_ (.RN(FE_OFN196_HRESETn), 
	.QN(U_dfifo_U_dcore_n5), 
	.Q(hiu_data[24]), 
	.D(FE_PHN920_U_dfifo_U_dcore_n158), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_27_ (.RN(FE_OFN196_HRESETn), 
	.QN(U_dfifo_U_dcore_n6), 
	.Q(hiu_data[25]), 
	.D(FE_PHN913_U_dfifo_U_dcore_n159), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_28_ (.RN(FE_OFN196_HRESETn), 
	.QN(U_dfifo_U_dcore_n12), 
	.Q(hiu_data[26]), 
	.D(FE_PHN911_U_dfifo_U_dcore_n160), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_29_ (.RN(FE_OFN196_HRESETn), 
	.QN(U_dfifo_U_dcore_n7), 
	.Q(hiu_data[27]), 
	.D(FE_PHN915_U_dfifo_U_dcore_n161), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_30_ (.RN(FE_OFN196_HRESETn), 
	.QN(U_dfifo_U_dcore_n8), 
	.Q(hiu_data[28]), 
	.D(FE_PHN912_U_dfifo_U_dcore_n162), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_31_ (.RN(FE_OFN196_HRESETn), 
	.QN(U_dfifo_U_dcore_n9), 
	.Q(hiu_data[29]), 
	.D(FE_PHN908_U_dfifo_U_dcore_n163), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_32_ (.RN(FE_OFN196_HRESETn), 
	.QN(U_dfifo_U_dcore_n10), 
	.Q(hiu_data[30]), 
	.D(FE_PHN914_U_dfifo_U_dcore_n164), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_33_ (.RN(FE_OFN196_HRESETn), 
	.QN(U_dfifo_U_dcore_n11), 
	.Q(hiu_data[31]), 
	.D(FE_PHN919_U_dfifo_U_dcore_n165), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_1_ (.RN(FE_OFN156_HRESETn), 
	.Q(U_dfifo_m_data_out_1_), 
	.D(FE_PHN903_U_dfifo_U_dcore_n166), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_0_ (.RN(FE_OFN43_HRESETn), 
	.Q(U_dfifo_m_data_out_0_), 
	.D(FE_PHN923_U_dfifo_U_dcore_n167), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_has_data_reg (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_n4), 
	.Q(U_dfifo_U_dcore_f_buf_has_data), 
	.D(FE_PHN3125_U_dfifo_U_dcore_n203), 
	.CK(HCLK__L5_N5));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_0_ (.RN(FE_OFN43_HRESETn), 
	.QN(n60), 
	.Q(U_dfifo_U_dcore_f_buf_data_0_), 
	.D(FE_PHN1579_U_dfifo_U_dcore_n168), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_1_ (.RN(FE_OFN156_HRESETn), 
	.QN(n59), 
	.Q(U_dfifo_U_dcore_f_buf_data_1_), 
	.D(FE_PHN1650_U_dfifo_U_dcore_n169), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_2_ (.RN(FE_OFN53_HRESETn), 
	.QN(n52), 
	.Q(U_dfifo_U_dcore_f_buf_data_2_), 
	.D(FE_PHN1246_U_dfifo_U_dcore_n170), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_3_ (.RN(FE_OFN28_HRESETn), 
	.QN(n58), 
	.Q(U_dfifo_U_dcore_f_buf_data_3_), 
	.D(FE_PHN1439_U_dfifo_U_dcore_n171), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_4_ (.RN(FE_OFN53_HRESETn), 
	.QN(n57), 
	.Q(U_dfifo_U_dcore_f_buf_data_4_), 
	.D(FE_PHN1442_U_dfifo_U_dcore_n172), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_5_ (.RN(FE_OFN53_HRESETn), 
	.QN(n56), 
	.Q(U_dfifo_U_dcore_f_buf_data_5_), 
	.D(FE_PHN1446_U_dfifo_U_dcore_n173), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_6_ (.RN(FE_OFN53_HRESETn), 
	.QN(n55), 
	.Q(U_dfifo_U_dcore_f_buf_data_6_), 
	.D(FE_PHN1440_U_dfifo_U_dcore_n174), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_7_ (.RN(FE_OFN53_HRESETn), 
	.QN(n54), 
	.Q(U_dfifo_U_dcore_f_buf_data_7_), 
	.D(FE_PHN1437_U_dfifo_U_dcore_n175), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_8_ (.RN(FE_OFN53_HRESETn), 
	.QN(n53), 
	.Q(U_dfifo_U_dcore_f_buf_data_8_), 
	.D(FE_PHN1438_U_dfifo_U_dcore_n176), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_9_ (.RN(FE_OFN53_HRESETn), 
	.QN(n67), 
	.Q(U_dfifo_U_dcore_f_buf_data_9_), 
	.D(FE_PHN1245_U_dfifo_U_dcore_n177), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_10_ (.RN(FE_OFN69_HRESETn), 
	.QN(n66), 
	.Q(U_dfifo_U_dcore_f_buf_data_10_), 
	.D(FE_PHN890_U_dfifo_U_dcore_n178), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_11_ (.RN(FE_OFN196_HRESETn), 
	.QN(n65), 
	.Q(U_dfifo_U_dcore_f_buf_data_11_), 
	.D(FE_PHN1436_U_dfifo_U_dcore_n179), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_12_ (.RN(FE_OFN196_HRESETn), 
	.QN(n64), 
	.Q(U_dfifo_U_dcore_f_buf_data_12_), 
	.D(FE_PHN1125_U_dfifo_U_dcore_n180), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_13_ (.RN(FE_OFN53_HRESETn), 
	.QN(n63), 
	.Q(U_dfifo_U_dcore_f_buf_data_13_), 
	.D(FE_PHN1441_U_dfifo_U_dcore_n181), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_14_ (.RN(FE_OFN69_HRESETn), 
	.QN(n62), 
	.Q(U_dfifo_U_dcore_f_buf_data_14_), 
	.D(FE_PHN1443_U_dfifo_U_dcore_n182), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_15_ (.RN(FE_OFN196_HRESETn), 
	.QN(n61), 
	.Q(U_dfifo_U_dcore_f_buf_data_15_), 
	.D(FE_PHN1434_U_dfifo_U_dcore_n183), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_16_ (.RN(FE_OFN196_HRESETn), 
	.QN(n83), 
	.Q(U_dfifo_U_dcore_f_buf_data_16_), 
	.D(FE_PHN1435_U_dfifo_U_dcore_n184), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_17_ (.RN(FE_OFN53_HRESETn), 
	.QN(n82), 
	.Q(U_dfifo_U_dcore_f_buf_data_17_), 
	.D(FE_PHN1244_U_dfifo_U_dcore_n185), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_18_ (.RN(FE_OFN69_HRESETn), 
	.QN(n81), 
	.Q(U_dfifo_U_dcore_f_buf_data_18_), 
	.D(FE_PHN1562_U_dfifo_U_dcore_n186), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_19_ (.RN(FE_OFN28_HRESETn), 
	.QN(n80), 
	.Q(U_dfifo_U_dcore_f_buf_data_19_), 
	.D(FE_PHN1466_U_dfifo_U_dcore_n187), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_20_ (.RN(FE_OFN157_HRESETn), 
	.QN(n79), 
	.Q(U_dfifo_U_dcore_f_buf_data_20_), 
	.D(FE_PHN1467_U_dfifo_U_dcore_n188), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_21_ (.RN(FE_OFN196_HRESETn), 
	.QN(n78), 
	.Q(U_dfifo_U_dcore_f_buf_data_21_), 
	.D(FE_PHN1459_U_dfifo_U_dcore_n189), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_22_ (.RN(FE_OFN196_HRESETn), 
	.QN(n77), 
	.Q(U_dfifo_U_dcore_f_buf_data_22_), 
	.D(FE_PHN1458_U_dfifo_U_dcore_n190), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_23_ (.RN(FE_OFN53_HRESETn), 
	.QN(n76), 
	.Q(U_dfifo_U_dcore_f_buf_data_23_), 
	.D(FE_PHN1464_U_dfifo_U_dcore_n191), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_24_ (.RN(FE_OFN53_HRESETn), 
	.QN(n75), 
	.Q(U_dfifo_U_dcore_f_buf_data_24_), 
	.D(FE_PHN1465_U_dfifo_U_dcore_n192), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_25_ (.RN(FE_OFN43_HRESETn), 
	.QN(n74), 
	.Q(U_dfifo_U_dcore_f_buf_data_25_), 
	.D(FE_PHN1550_U_dfifo_U_dcore_n193), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_26_ (.RN(FE_OFN43_HRESETn), 
	.QN(n85), 
	.Q(U_dfifo_U_dcore_f_buf_data_26_), 
	.D(FE_PHN1547_U_dfifo_U_dcore_n194), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_27_ (.RN(FE_OFN43_HRESETn), 
	.QN(n84), 
	.Q(U_dfifo_U_dcore_f_buf_data_27_), 
	.D(FE_PHN1452_U_dfifo_U_dcore_n195), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_28_ (.RN(FE_OFN43_HRESETn), 
	.QN(n73), 
	.Q(U_dfifo_U_dcore_f_buf_data_28_), 
	.D(FE_PHN1453_U_dfifo_U_dcore_n196), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_29_ (.RN(FE_OFN43_HRESETn), 
	.QN(n72), 
	.Q(U_dfifo_U_dcore_f_buf_data_29_), 
	.D(FE_PHN1454_U_dfifo_U_dcore_n197), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_30_ (.RN(FE_OFN43_HRESETn), 
	.QN(n71), 
	.Q(U_dfifo_U_dcore_f_buf_data_30_), 
	.D(FE_PHN1451_U_dfifo_U_dcore_n198), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_31_ (.RN(FE_OFN62_HRESETn), 
	.QN(n70), 
	.Q(U_dfifo_U_dcore_f_buf_data_31_), 
	.D(FE_PHN1248_U_dfifo_U_dcore_n199), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_32_ (.RN(FE_OFN43_HRESETn), 
	.QN(n68), 
	.Q(U_dfifo_U_dcore_f_buf_data_32_), 
	.D(FE_PHN1250_U_dfifo_U_dcore_n200), 
	.CK(HCLK__L5_N5));
   DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_33_ (.RN(FE_OFN43_HRESETn), 
	.QN(n69), 
	.Q(U_dfifo_U_dcore_f_buf_data_33_), 
	.D(FE_PHN1544_U_dfifo_U_dcore_n201), 
	.CK(HCLK__L5_N14));
   DFFS_X2 U_dfifo_U_dcore_f_empty_reg (.SN(FE_OFN54_HRESETn), 
	.Q(U_dfifo_m_empty), 
	.D(FE_PHN4384_U_dfifo_U_dcore_n_empty), 
	.CK(HCLK__L5_N6));
   AOI22_X1 U_afifo_U_acore_U_sub_fifo_U276 (.ZN(U_afifo_U_acore_U_sub_fifo_n372), 
	.B2(U_afifo_U_acore_n166), 
	.B1(FE_PHN2979_U_afifo_U_acore_U_sub_fifo_count_0_), 
	.A2(U_afifo_U_acore_U_sub_fifo_n371), 
	.A1(FE_PHN867_U_afifo_U_acore_U_sub_fifo_count_1_));
   NOR2_X1 U_afifo_U_acore_U_sub_fifo_U275 (.ZN(U_afifo_U_acore_U_sub_fifo_n371), 
	.A2(U_afifo_U_acore_n166), 
	.A1(FE_PHN2979_U_afifo_U_acore_U_sub_fifo_count_0_));
   OAI21_X1 U_afifo_U_acore_U_sub_fifo_U274 (.ZN(U_afifo_U_acore_U_sub_fifo_n324), 
	.B2(FE_PHN1049_U_afifo_U_acore_U_sub_fifo_n11), 
	.B1(U_afifo_U_acore_U_sub_fifo_n370), 
	.A(U_afifo_U_acore_U_sub_fifo_n1));
   OAI21_X1 U_afifo_U_acore_U_sub_fifo_U273 (.ZN(U_afifo_U_acore_U_sub_fifo_n323), 
	.B2(FE_PHN993_U_afifo_U_acore_U_sub_fifo_n149), 
	.B1(U_afifo_U_acore_U_sub_fifo_n370), 
	.A(U_afifo_U_acore_U_sub_fifo_n369));
   OAI21_X1 U_afifo_U_acore_U_sub_fifo_U272 (.ZN(U_afifo_U_acore_U_sub_fifo_n165), 
	.B2(U_afifo_U_acore_U_sub_fifo_n167), 
	.B1(U_afifo_U_acore_n166), 
	.A(FE_PHN867_U_afifo_U_acore_U_sub_fifo_count_1_));
   NAND2_X1 U_afifo_U_acore_U_sub_fifo_U271 (.ZN(U_afifo_U_acore_U_sub_fifo_n166), 
	.A2(U_afifo_U_acore_n166), 
	.A1(FE_PHN2979_U_afifo_U_acore_U_sub_fifo_count_0_));
   NAND3_X2 U_afifo_U_acore_U_sub_fifo_U270 (.ZN(U_afifo_U_acore_U_sub_fifo_n169), 
	.A3(U_afifo_U_acore_U_sub_fifo_n370), 
	.A2(U_afifo_U_acore_U_sub_fifo_in_ptr_1_), 
	.A1(FE_PHN993_U_afifo_U_acore_U_sub_fifo_n149));
   NAND3_X2 U_afifo_U_acore_U_sub_fifo_U269 (.ZN(U_afifo_U_acore_U_sub_fifo_n369), 
	.A3(U_afifo_U_acore_U_sub_fifo_n370), 
	.A2(FE_PHN993_U_afifo_U_acore_U_sub_fifo_n149), 
	.A1(FE_PHN1049_U_afifo_U_acore_U_sub_fifo_n11));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U267 (.ZN(U_afifo_U_acore_m_sf_data_out[18]), 
	.C2(FE_OFN263_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n7), 
	.B2(U_afifo_U_acore_U_sub_fifo_n57), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n132), 
	.A1(U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U266 (.ZN(U_afifo_U_acore_m_sf_data_out[28]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n28), 
	.B2(U_afifo_U_acore_U_sub_fifo_n77), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1822_U_afifo_U_acore_U_sub_fifo_n122), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U265 (.ZN(U_afifo_U_acore_m_sf_data_out[27]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n29), 
	.B2(U_afifo_U_acore_U_sub_fifo_n78), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1812_U_afifo_U_acore_U_sub_fifo_n123), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U264 (.ZN(U_afifo_U_acore_m_sf_data_out[25]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n6), 
	.B2(U_afifo_U_acore_U_sub_fifo_n56), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1827_U_afifo_U_acore_U_sub_fifo_n125), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U263 (.ZN(U_afifo_U_acore_m_sf_data_out[29]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n27), 
	.B2(U_afifo_U_acore_U_sub_fifo_n76), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1810_U_afifo_U_acore_U_sub_fifo_n121), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U262 (.ZN(U_afifo_U_acore_m_sf_data_out[26]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n30), 
	.B2(U_afifo_U_acore_U_sub_fifo_n79), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1792_U_afifo_U_acore_U_sub_fifo_n124), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   INV_X4 U_afifo_U_acore_U_sub_fifo_U261 (.ZN(U_afifo_U_acore_U_sub_fifo_n150), 
	.A(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   INV_X4 U_afifo_U_acore_U_sub_fifo_U260 (.ZN(U_afifo_U_acore_U_sub_fifo_n151), 
	.A(U_afifo_U_acore_U_sub_fifo_n150));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U259 (.ZN(U_afifo_U_acore_m_sf_data_out[24]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n31), 
	.B2(U_afifo_U_acore_U_sub_fifo_n80), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1843_U_afifo_U_acore_U_sub_fifo_n126), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U258 (.ZN(U_afifo_U_acore_m_sf_data_out[23]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n32), 
	.B2(U_afifo_U_acore_U_sub_fifo_n81), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1805_U_afifo_U_acore_U_sub_fifo_n127), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U257 (.ZN(U_afifo_U_acore_m_sf_data_out[22]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n33), 
	.B2(U_afifo_U_acore_U_sub_fifo_n82), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1806_U_afifo_U_acore_U_sub_fifo_n128), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U256 (.ZN(U_afifo_U_acore_m_sf_data_out[20]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n35), 
	.B2(U_afifo_U_acore_U_sub_fifo_n84), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1828_U_afifo_U_acore_U_sub_fifo_n130), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U255 (.ZN(U_afifo_U_acore_m_sf_data_out[19]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n36), 
	.B2(U_afifo_U_acore_U_sub_fifo_n85), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1797_U_afifo_U_acore_U_sub_fifo_n131), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U254 (.ZN(U_afifo_U_acore_m_sf_data_out[21]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n34), 
	.B2(U_afifo_U_acore_U_sub_fifo_n83), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1832_U_afifo_U_acore_U_sub_fifo_n129), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U253 (.ZN(U_afifo_U_acore_m_sf_data_out[34]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n23), 
	.B2(U_afifo_U_acore_U_sub_fifo_n72), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n116), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U252 (.ZN(U_afifo_U_acore_m_sf_data_out[37]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n4), 
	.B2(U_afifo_U_acore_U_sub_fifo_n54), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n113), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U251 (.ZN(U_afifo_U_acore_m_sf_data_out[36]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n21), 
	.B2(U_afifo_U_acore_U_sub_fifo_n70), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n114), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U250 (.ZN(U_afifo_U_acore_m_sf_data_out[30]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n26), 
	.B2(U_afifo_U_acore_U_sub_fifo_n75), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1796_U_afifo_U_acore_U_sub_fifo_n120), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U249 (.ZN(U_afifo_U_acore_m_sf_data_out[38]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n20), 
	.B2(U_afifo_U_acore_U_sub_fifo_n69), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n112), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U248 (.ZN(U_afifo_U_acore_m_sf_data_out[33]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n24), 
	.B2(U_afifo_U_acore_U_sub_fifo_n73), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n117), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U247 (.ZN(U_afifo_U_acore_m_sf_data_out[35]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n22), 
	.B2(U_afifo_U_acore_U_sub_fifo_n71), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1831_U_afifo_U_acore_U_sub_fifo_n115), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U246 (.ZN(U_afifo_U_acore_m_sf_data_out[39]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n19), 
	.B2(U_afifo_U_acore_U_sub_fifo_n68), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n111), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U245 (.ZN(U_afifo_U_acore_m_sf_data_out[31]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n25), 
	.B2(U_afifo_U_acore_U_sub_fifo_n74), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n119), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U244 (.ZN(U_afifo_U_acore_m_sf_data_out[32]), 
	.C2(FE_OFN262_U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n5), 
	.B2(U_afifo_U_acore_U_sub_fifo_n55), 
	.B1(FE_OFN261_U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n118), 
	.A1(FE_OFN202_U_afifo_U_acore_U_sub_fifo_n162));
   INV_X4 U_afifo_U_acore_U_sub_fifo_U242 (.ZN(U_afifo_U_acore_U_sub_fifo_n167), 
	.A(U_afifo_U_acore_n165));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U241 (.ZN(U_afifo_U_acore_U_sub_fifo_n231), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n17), 
	.A2(FE_PHN1192_U_afifo_U_acore_n68), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U239 (.ZN(U_afifo_U_acore_U_sub_fifo_n261), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n42), 
	.A2(U_afifo_U_acore_n31), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U238 (.ZN(U_afifo_U_acore_U_sub_fifo_n233), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n19), 
	.A2(FE_PHN1197_U_afifo_U_acore_n72), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U237 (.ZN(U_afifo_U_acore_U_sub_fifo_n242), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n26), 
	.A2(FE_PHN1405_U_afifo_U_acore_n90), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U236 (.ZN(U_afifo_U_acore_U_sub_fifo_n239), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n24), 
	.A2(FE_PHN1190_U_afifo_U_acore_n84), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U235 (.ZN(U_afifo_U_acore_U_sub_fifo_n236), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n21), 
	.A2(FE_PHN1191_U_afifo_U_acore_n78), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U234 (.ZN(U_afifo_U_acore_U_sub_fifo_n254), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n7), 
	.A2(FE_PHN1189_U_afifo_U_acore_n167), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U233 (.ZN(U_afifo_U_acore_U_sub_fifo_n232), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n18), 
	.A2(FE_PHN1186_U_afifo_U_acore_n70), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U232 (.ZN(U_afifo_U_acore_U_sub_fifo_n234), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n20), 
	.A2(FE_PHN1194_U_afifo_U_acore_n74), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U231 (.ZN(U_afifo_U_acore_U_sub_fifo_n238), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n23), 
	.A2(FE_PHN1187_U_afifo_U_acore_n82), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U230 (.ZN(U_afifo_U_acore_U_sub_fifo_n241), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n25), 
	.A2(FE_PHN1193_U_afifo_U_acore_n88), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U229 (.ZN(U_afifo_U_acore_U_sub_fifo_n240), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n5), 
	.A2(FE_PHN1188_U_afifo_U_acore_n86), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U228 (.ZN(U_afifo_U_acore_U_sub_fifo_n237), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n22), 
	.A2(FE_PHN1552_U_afifo_U_acore_n80), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U226 (.ZN(U_afifo_U_acore_U_sub_fifo_n227), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n14), 
	.A2(U_afifo_U_acore_n30), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U224 (.ZN(U_afifo_U_acore_U_sub_fifo_n263), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n43), 
	.A2(U_afifo_U_acore_n32), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U222 (.ZN(U_afifo_U_acore_U_sub_fifo_n226), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n13), 
	.A2(FE_PHN3423_U_afifo_U_acore_n29), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U221 (.ZN(U_afifo_U_acore_U_sub_fifo_n235), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n4), 
	.A2(FE_PHN1406_U_afifo_U_acore_n76), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U219 (.ZN(U_afifo_U_acore_U_sub_fifo_n253), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n36), 
	.A2(FE_PHN3263_U_afifo_U_acore_n162), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U217 (.ZN(U_afifo_U_acore_U_sub_fifo_n256), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n38), 
	.A2(FE_PHN3243_U_afifo_U_acore_n199), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U215 (.ZN(U_afifo_U_acore_U_sub_fifo_n250), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n33), 
	.A2(FE_PHN3384_U_afifo_U_acore_n156), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U213 (.ZN(U_afifo_U_acore_U_sub_fifo_n230), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n16), 
	.A2(FE_PHN1840_U_afifo_U_acore_n194), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U211 (.ZN(U_afifo_U_acore_U_sub_fifo_n258), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n40), 
	.A2(FE_PHN1839_U_afifo_U_acore_n203), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U209 (.ZN(U_afifo_U_acore_U_sub_fifo_n249), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n32), 
	.A2(FE_PHN3409_U_afifo_U_acore_n153), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U207 (.ZN(U_afifo_U_acore_U_sub_fifo_n251), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n34), 
	.A2(FE_PHN3412_U_afifo_U_acore_n158), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U205 (.ZN(U_afifo_U_acore_U_sub_fifo_n243), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n27), 
	.A2(FE_PHN3248_U_afifo_U_acore_n94), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U203 (.ZN(U_afifo_U_acore_U_sub_fifo_n246), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n30), 
	.A2(FE_PHN1852_U_afifo_U_acore_n100), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U201 (.ZN(U_afifo_U_acore_U_sub_fifo_n225), 
	.B2(U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n61), 
	.A2(FE_PHN1564_U_afifo_U_acore_n186), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U199 (.ZN(U_afifo_U_acore_U_sub_fifo_n252), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n35), 
	.A2(FE_PHN3262_U_afifo_U_acore_n160), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U197 (.ZN(U_afifo_U_acore_U_sub_fifo_n259), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n8), 
	.A2(FE_PHN1561_U_afifo_U_acore_n205), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U195 (.ZN(U_afifo_U_acore_U_sub_fifo_n244), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n28), 
	.A2(FE_PHN1851_U_afifo_U_acore_n96), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U193 (.ZN(U_afifo_U_acore_U_sub_fifo_n247), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n6), 
	.A2(FE_PHN1837_U_afifo_U_acore_n102), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U191 (.ZN(U_afifo_U_acore_U_sub_fifo_n260), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n41), 
	.A2(FE_PHN1849_U_afifo_U_acore_n207), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U189 (.ZN(U_afifo_U_acore_U_sub_fifo_n248), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n31), 
	.A2(FE_PHN3257_U_afifo_U_acore_n104), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U187 (.ZN(U_afifo_U_acore_U_sub_fifo_n257), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n39), 
	.A2(FE_PHN1844_U_afifo_U_acore_n201), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U185 (.ZN(U_afifo_U_acore_U_sub_fifo_n264), 
	.B2(U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n44), 
	.A2(FE_PHN1408_U_afifo_U_acore_n173), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U183 (.ZN(U_afifo_U_acore_U_sub_fifo_n229), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n15), 
	.A2(FE_PHN1563_U_afifo_U_acore_n192), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U181 (.ZN(U_afifo_U_acore_U_sub_fifo_n255), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n37), 
	.A2(FE_PHN1835_U_afifo_U_acore_n197), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U179 (.ZN(U_afifo_U_acore_U_sub_fifo_n245), 
	.B2(FE_OFN203_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n29), 
	.A2(FE_PHN1850_U_afifo_U_acore_n98), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U177 (.ZN(U_afifo_U_acore_U_sub_fifo_n265), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n45), 
	.A2(FE_PHN1560_U_afifo_U_acore_n175), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U175 (.ZN(U_afifo_U_acore_U_sub_fifo_n228), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n3), 
	.A2(FE_PHN1558_U_afifo_U_acore_n190), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U173 (.ZN(U_afifo_U_acore_U_sub_fifo_n267), 
	.B2(U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n9), 
	.A2(FE_PHN1554_U_afifo_U_acore_n179), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U171 (.ZN(U_afifo_U_acore_U_sub_fifo_n266), 
	.B2(U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n46), 
	.A2(FE_PHN1834_U_afifo_U_acore_n177), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U169 (.ZN(U_afifo_U_acore_U_sub_fifo_n269), 
	.B2(U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n48), 
	.A2(FE_PHN3261_U_afifo_U_acore_n33), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U168 (.ZN(U_afifo_U_acore_U_sub_fifo_n270), 
	.B2(U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n49), 
	.A2(FE_PHN1404_U_afifo_U_acore_n92), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U166 (.ZN(U_afifo_U_acore_U_sub_fifo_n268), 
	.B2(U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n47), 
	.A2(FE_PHN1847_U_afifo_U_acore_n181), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U164 (.ZN(U_afifo_U_acore_U_sub_fifo_n272), 
	.B2(U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n50), 
	.A2(FE_PHN1836_U_afifo_U_acore_n210), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U163 (.ZN(U_afifo_U_acore_m_sf_data_out[17]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n37), 
	.B2(U_afifo_U_acore_U_sub_fifo_n86), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1833_U_afifo_U_acore_U_sub_fifo_n133), 
	.A1(U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U162 (.ZN(U_afifo_U_acore_m_sf_data_out[16]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n38), 
	.B2(U_afifo_U_acore_U_sub_fifo_n87), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1826_U_afifo_U_acore_U_sub_fifo_n134), 
	.A1(U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U161 (.ZN(U_afifo_U_acore_m_sf_data_out[15]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n39), 
	.B2(U_afifo_U_acore_U_sub_fifo_n88), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1799_U_afifo_U_acore_U_sub_fifo_n135), 
	.A1(U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U160 (.ZN(U_afifo_U_acore_m_sf_data_out[14]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n40), 
	.B2(U_afifo_U_acore_U_sub_fifo_n89), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1821_U_afifo_U_acore_U_sub_fifo_n136), 
	.A1(U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U159 (.ZN(U_afifo_U_acore_m_sf_data_out[0]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n50), 
	.B2(U_afifo_U_acore_U_sub_fifo_n99), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1830_U_afifo_U_acore_U_sub_fifo_n148), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U158 (.ZN(U_afifo_U_acore_m_sf_data_out[13]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n8), 
	.B2(U_afifo_U_acore_U_sub_fifo_n58), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n137), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U157 (.ZN(U_afifo_U_acore_m_sf_data_out[12]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n41), 
	.B2(U_afifo_U_acore_U_sub_fifo_n90), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1814_U_afifo_U_acore_U_sub_fifo_n138), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U156 (.ZN(U_afifo_U_acore_m_sf_data_out[43]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n15), 
	.B2(U_afifo_U_acore_U_sub_fifo_n64), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n107), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U155 (.ZN(U_afifo_U_acore_m_sf_data_out[11]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n42), 
	.B2(U_afifo_U_acore_U_sub_fifo_n91), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1820_U_afifo_U_acore_U_sub_fifo_n139), 
	.A1(U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U154 (.ZN(U_afifo_U_acore_m_sf_data_out[46]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n13), 
	.B2(U_afifo_U_acore_U_sub_fifo_n62), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1793_U_afifo_U_acore_U_sub_fifo_n104), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U153 (.ZN(U_afifo_U_acore_m_sf_data_out[47]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n61), 
	.B2(U_afifo_U_acore_U_sub_fifo_n52), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n103), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U152 (.ZN(U_afifo_U_acore_m_sf_data_out[42]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n16), 
	.B2(U_afifo_U_acore_U_sub_fifo_n65), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1801_U_afifo_U_acore_U_sub_fifo_n108), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U151 (.ZN(U_afifo_U_acore_m_sf_data_out[3]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n48), 
	.B2(U_afifo_U_acore_U_sub_fifo_n97), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1804_U_afifo_U_acore_U_sub_fifo_n146), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U150 (.ZN(U_afifo_U_acore_m_sf_data_out[5]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n9), 
	.B2(U_afifo_U_acore_U_sub_fifo_n59), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n144), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U149 (.ZN(U_afifo_U_acore_m_sf_data_out[44]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n3), 
	.B2(U_afifo_U_acore_U_sub_fifo_n53), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1825_U_afifo_U_acore_U_sub_fifo_n106), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U148 (.ZN(U_afifo_U_acore_m_sf_data_out[4]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n47), 
	.B2(U_afifo_U_acore_U_sub_fifo_n96), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1800_U_afifo_U_acore_U_sub_fifo_n145), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U147 (.ZN(U_afifo_U_acore_m_sf_data_out[9]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n43), 
	.B2(U_afifo_U_acore_U_sub_fifo_n92), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1808_U_afifo_U_acore_U_sub_fifo_n140), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U146 (.ZN(U_afifo_U_acore_m_sf_data_out[45]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n14), 
	.B2(U_afifo_U_acore_U_sub_fifo_n63), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n105), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U145 (.ZN(U_afifo_U_acore_m_sf_data_out[48]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n60), 
	.B2(U_afifo_U_acore_U_sub_fifo_n51), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1816_U_afifo_U_acore_U_sub_fifo_n102), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U144 (.ZN(U_afifo_U_acore_m_sf_data_out[7]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n45), 
	.B2(U_afifo_U_acore_U_sub_fifo_n94), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n142), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U143 (.ZN(U_afifo_U_acore_m_sf_data_out[49]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n12), 
	.B2(U_afifo_U_acore_U_sub_fifo_n101), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n2), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U142 (.ZN(U_afifo_U_acore_m_sf_data_out[6]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n46), 
	.B2(U_afifo_U_acore_U_sub_fifo_n95), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(FE_PHN1815_U_afifo_U_acore_U_sub_fifo_n143), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U141 (.ZN(U_afifo_U_acore_m_sf_data_out[8]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n44), 
	.B2(U_afifo_U_acore_U_sub_fifo_n93), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n141), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U139 (.ZN(U_afifo_U_acore_U_sub_fifo_n223), 
	.B2(U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n12), 
	.A2(U_afifo_U_acore_n28), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U137 (.ZN(U_afifo_U_acore_U_sub_fifo_n224), 
	.B2(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1), 
	.B1(U_afifo_U_acore_U_sub_fifo_n60), 
	.A2(FE_PHN1841_U_afifo_U_acore_n184), 
	.A1(U_afifo_U_acore_U_sub_fifo_n153));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U136 (.ZN(U_afifo_U_acore_m_sf_data_out[41]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n17), 
	.B2(U_afifo_U_acore_U_sub_fifo_n66), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n109), 
	.A1(U_afifo_U_acore_U_sub_fifo_n162));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U135 (.ZN(U_afifo_U_acore_m_sf_data_out[40]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n18), 
	.B2(U_afifo_U_acore_U_sub_fifo_n67), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n110), 
	.A1(U_afifo_U_acore_U_sub_fifo_n151));
   OAI222_X2 U_afifo_U_acore_U_sub_fifo_U134 (.ZN(U_afifo_U_acore_m_sf_data_out[2]), 
	.C2(U_afifo_U_acore_U_sub_fifo_n161), 
	.C1(U_afifo_U_acore_U_sub_fifo_n49), 
	.B2(U_afifo_U_acore_U_sub_fifo_n98), 
	.B1(U_afifo_U_acore_U_sub_fifo_n163), 
	.A2(U_afifo_U_acore_U_sub_fifo_n147), 
	.A1(FE_OFN7_U_afifo_U_acore_U_sub_fifo_n162));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U133 (.ZN(U_afifo_U_acore_U_sub_fifo_n187), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n71), 
	.A2(FE_PHN1552_U_afifo_U_acore_n80), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U132 (.ZN(U_afifo_U_acore_U_sub_fifo_n192), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n75), 
	.A2(FE_PHN1405_U_afifo_U_acore_n90), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U131 (.ZN(U_afifo_U_acore_U_sub_fifo_n183), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n68), 
	.A2(FE_PHN1197_U_afifo_U_acore_n72), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U130 (.ZN(U_afifo_U_acore_U_sub_fifo_n190), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n55), 
	.A2(FE_PHN1188_U_afifo_U_acore_n86), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U129 (.ZN(U_afifo_U_acore_U_sub_fifo_n188), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n72), 
	.A2(FE_PHN1187_U_afifo_U_acore_n82), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U128 (.ZN(U_afifo_U_acore_U_sub_fifo_n181), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n66), 
	.A2(FE_PHN1192_U_afifo_U_acore_n68), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U127 (.ZN(U_afifo_U_acore_U_sub_fifo_n186), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n70), 
	.A2(FE_PHN1191_U_afifo_U_acore_n78), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U126 (.ZN(U_afifo_U_acore_U_sub_fifo_n185), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n54), 
	.A2(FE_PHN1406_U_afifo_U_acore_n76), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U125 (.ZN(U_afifo_U_acore_U_sub_fifo_n184), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n69), 
	.A2(FE_PHN1194_U_afifo_U_acore_n74), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U124 (.ZN(U_afifo_U_acore_U_sub_fifo_n182), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n67), 
	.A2(FE_PHN1186_U_afifo_U_acore_n70), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U123 (.ZN(U_afifo_U_acore_U_sub_fifo_n191), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n74), 
	.A2(FE_PHN1193_U_afifo_U_acore_n88), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U122 (.ZN(U_afifo_U_acore_U_sub_fifo_n173), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n101), 
	.A2(U_afifo_U_acore_n28), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U121 (.ZN(U_afifo_U_acore_U_sub_fifo_n201), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n83), 
	.A2(FE_PHN3412_U_afifo_U_acore_n158), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U120 (.ZN(U_afifo_U_acore_U_sub_fifo_n180), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n65), 
	.A2(FE_PHN1840_U_afifo_U_acore_n194), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U119 (.ZN(U_afifo_U_acore_U_sub_fifo_n209), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n58), 
	.A2(FE_PHN1561_U_afifo_U_acore_n205), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U118 (.ZN(U_afifo_U_acore_U_sub_fifo_n179), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n64), 
	.A2(FE_PHN1563_U_afifo_U_acore_n192), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U117 (.ZN(U_afifo_U_acore_U_sub_fifo_n178), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n53), 
	.A2(FE_PHN1558_U_afifo_U_acore_n190), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U116 (.ZN(U_afifo_U_acore_U_sub_fifo_n200), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n82), 
	.A2(FE_PHN3384_U_afifo_U_acore_n156), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U115 (.ZN(U_afifo_U_acore_U_sub_fifo_n177), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n63), 
	.A2(U_afifo_U_acore_n30), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U114 (.ZN(U_afifo_U_acore_U_sub_fifo_n176), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n62), 
	.A2(FE_PHN3423_U_afifo_U_acore_n29), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U113 (.ZN(U_afifo_U_acore_U_sub_fifo_n175), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n52), 
	.A2(FE_PHN1564_U_afifo_U_acore_n186), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U112 (.ZN(U_afifo_U_acore_U_sub_fifo_n174), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n51), 
	.A2(FE_PHN1841_U_afifo_U_acore_n184), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U111 (.ZN(U_afifo_U_acore_U_sub_fifo_n193), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n76), 
	.A2(FE_PHN3248_U_afifo_U_acore_n94), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U110 (.ZN(U_afifo_U_acore_U_sub_fifo_n194), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n77), 
	.A2(FE_PHN1851_U_afifo_U_acore_n96), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U109 (.ZN(U_afifo_U_acore_U_sub_fifo_n211), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n91), 
	.A2(U_afifo_U_acore_n31), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U108 (.ZN(U_afifo_U_acore_U_sub_fifo_n198), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n80), 
	.A2(FE_PHN3257_U_afifo_U_acore_n104), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U107 (.ZN(U_afifo_U_acore_U_sub_fifo_n195), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n78), 
	.A2(FE_PHN1850_U_afifo_U_acore_n98), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U106 (.ZN(U_afifo_U_acore_U_sub_fifo_n219), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n97), 
	.A2(FE_PHN3261_U_afifo_U_acore_n33), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U105 (.ZN(U_afifo_U_acore_U_sub_fifo_n199), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n81), 
	.A2(FE_PHN3409_U_afifo_U_acore_n153), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U104 (.ZN(U_afifo_U_acore_U_sub_fifo_n196), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n79), 
	.A2(FE_PHN1852_U_afifo_U_acore_n100), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U103 (.ZN(U_afifo_U_acore_U_sub_fifo_n208), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n89), 
	.A2(FE_PHN1839_U_afifo_U_acore_n203), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U102 (.ZN(U_afifo_U_acore_U_sub_fifo_n217), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n59), 
	.A2(FE_PHN1554_U_afifo_U_acore_n179), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U101 (.ZN(U_afifo_U_acore_U_sub_fifo_n210), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n90), 
	.A2(FE_PHN1849_U_afifo_U_acore_n207), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U100 (.ZN(U_afifo_U_acore_U_sub_fifo_n202), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n84), 
	.A2(FE_PHN3262_U_afifo_U_acore_n160), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U99 (.ZN(U_afifo_U_acore_U_sub_fifo_n203), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n85), 
	.A2(FE_PHN3263_U_afifo_U_acore_n162), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U98 (.ZN(U_afifo_U_acore_U_sub_fifo_n216), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n95), 
	.A2(FE_PHN1834_U_afifo_U_acore_n177), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U97 (.ZN(U_afifo_U_acore_U_sub_fifo_n204), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n57), 
	.A2(FE_PHN1189_U_afifo_U_acore_n167), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U96 (.ZN(U_afifo_U_acore_U_sub_fifo_n205), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n86), 
	.A2(FE_PHN1835_U_afifo_U_acore_n197), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U95 (.ZN(U_afifo_U_acore_U_sub_fifo_n215), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n94), 
	.A2(FE_PHN1560_U_afifo_U_acore_n175), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U94 (.ZN(U_afifo_U_acore_U_sub_fifo_n206), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n87), 
	.A2(FE_PHN3243_U_afifo_U_acore_n199), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U93 (.ZN(U_afifo_U_acore_U_sub_fifo_n214), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n93), 
	.A2(FE_PHN1408_U_afifo_U_acore_n173), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U92 (.ZN(U_afifo_U_acore_U_sub_fifo_n207), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n88), 
	.A2(FE_PHN1844_U_afifo_U_acore_n201), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U91 (.ZN(U_afifo_U_acore_U_sub_fifo_n213), 
	.B2(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n92), 
	.A2(U_afifo_U_acore_n32), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U90 (.ZN(U_afifo_U_acore_U_sub_fifo_n220), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n98), 
	.A2(FE_PHN1404_U_afifo_U_acore_n92), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U89 (.ZN(U_afifo_U_acore_U_sub_fifo_n189), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n73), 
	.A2(FE_PHN1190_U_afifo_U_acore_n84), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U88 (.ZN(U_afifo_U_acore_U_sub_fifo_n222), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n99), 
	.A2(FE_PHN1836_U_afifo_U_acore_n210), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U87 (.ZN(U_afifo_U_acore_U_sub_fifo_n218), 
	.B2(U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n96), 
	.A2(FE_PHN1847_U_afifo_U_acore_n181), 
	.A1(U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U86 (.ZN(U_afifo_U_acore_U_sub_fifo_n197), 
	.B2(FE_OFN207_U_afifo_U_acore_U_sub_fifo_n169), 
	.B1(U_afifo_U_acore_U_sub_fifo_n56), 
	.A2(FE_PHN1837_U_afifo_U_acore_n102), 
	.A1(FE_OFN260_U_afifo_U_acore_U_sub_fifo_n212));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U85 (.ZN(U_afifo_U_acore_U_sub_fifo_n319), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1804_U_afifo_U_acore_U_sub_fifo_n146), 
	.A2(FE_PHN3261_U_afifo_U_acore_n33), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U84 (.ZN(U_afifo_U_acore_U_sub_fifo_n281), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n109), 
	.A2(FE_PHN1192_U_afifo_U_acore_n68), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U83 (.ZN(U_afifo_U_acore_U_sub_fifo_n322), 
	.B2(U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1830_U_afifo_U_acore_U_sub_fifo_n148), 
	.A2(FE_PHN1836_U_afifo_U_acore_n210), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U82 (.ZN(U_afifo_U_acore_U_sub_fifo_n279), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n107), 
	.A2(FE_PHN1563_U_afifo_U_acore_n192), 
	.A1(FE_OFN264_U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U81 (.ZN(U_afifo_U_acore_U_sub_fifo_n317), 
	.B2(U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n144), 
	.A2(FE_PHN1554_U_afifo_U_acore_n179), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U80 (.ZN(U_afifo_U_acore_U_sub_fifo_n276), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1793_U_afifo_U_acore_U_sub_fifo_n104), 
	.A2(FE_PHN3423_U_afifo_U_acore_n29), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U79 (.ZN(U_afifo_U_acore_U_sub_fifo_n275), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n103), 
	.A2(FE_PHN1564_U_afifo_U_acore_n186), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U78 (.ZN(U_afifo_U_acore_U_sub_fifo_n318), 
	.B2(U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1800_U_afifo_U_acore_U_sub_fifo_n145), 
	.A2(FE_PHN1847_U_afifo_U_acore_n181), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U77 (.ZN(U_afifo_U_acore_U_sub_fifo_n278), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1825_U_afifo_U_acore_U_sub_fifo_n106), 
	.A2(FE_PHN1558_U_afifo_U_acore_n190), 
	.A1(FE_OFN264_U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U76 (.ZN(U_afifo_U_acore_U_sub_fifo_n285), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n113), 
	.A2(FE_PHN1406_U_afifo_U_acore_n76), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U75 (.ZN(U_afifo_U_acore_U_sub_fifo_n280), 
	.B2(U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1801_U_afifo_U_acore_U_sub_fifo_n108), 
	.A2(FE_PHN1840_U_afifo_U_acore_n194), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U74 (.ZN(U_afifo_U_acore_U_sub_fifo_n320), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n147), 
	.A2(FE_PHN1404_U_afifo_U_acore_n92), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U73 (.ZN(U_afifo_U_acore_U_sub_fifo_n286), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n114), 
	.A2(FE_PHN1191_U_afifo_U_acore_n78), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U72 (.ZN(U_afifo_U_acore_U_sub_fifo_n283), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n111), 
	.A2(FE_PHN1197_U_afifo_U_acore_n72), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U71 (.ZN(U_afifo_U_acore_U_sub_fifo_n284), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n112), 
	.A2(FE_PHN1194_U_afifo_U_acore_n74), 
	.A1(FE_OFN264_U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U70 (.ZN(U_afifo_U_acore_U_sub_fifo_n316), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1815_U_afifo_U_acore_U_sub_fifo_n143), 
	.A2(FE_PHN1834_U_afifo_U_acore_n177), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U69 (.ZN(U_afifo_U_acore_U_sub_fifo_n282), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n110), 
	.A2(FE_PHN1186_U_afifo_U_acore_n70), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U68 (.ZN(U_afifo_U_acore_U_sub_fifo_n273), 
	.B2(U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n2), 
	.A2(U_afifo_U_acore_n28), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U67 (.ZN(U_afifo_U_acore_U_sub_fifo_n289), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n117), 
	.A2(FE_PHN1190_U_afifo_U_acore_n84), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U66 (.ZN(U_afifo_U_acore_U_sub_fifo_n296), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1792_U_afifo_U_acore_U_sub_fifo_n124), 
	.A2(FE_PHN1852_U_afifo_U_acore_n100), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U65 (.ZN(U_afifo_U_acore_U_sub_fifo_n309), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n137), 
	.A2(FE_PHN1561_U_afifo_U_acore_n205), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U64 (.ZN(U_afifo_U_acore_U_sub_fifo_n290), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n118), 
	.A2(FE_PHN1188_U_afifo_U_acore_n86), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U63 (.ZN(U_afifo_U_acore_U_sub_fifo_n301), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1832_U_afifo_U_acore_U_sub_fifo_n129), 
	.A2(FE_PHN3412_U_afifo_U_acore_n158), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U62 (.ZN(U_afifo_U_acore_U_sub_fifo_n303), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1797_U_afifo_U_acore_U_sub_fifo_n131), 
	.A2(FE_PHN3263_U_afifo_U_acore_n162), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U61 (.ZN(U_afifo_U_acore_U_sub_fifo_n293), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1810_U_afifo_U_acore_U_sub_fifo_n121), 
	.A2(FE_PHN3248_U_afifo_U_acore_n94), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U60 (.ZN(U_afifo_U_acore_U_sub_fifo_n292), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1796_U_afifo_U_acore_U_sub_fifo_n120), 
	.A2(FE_PHN1405_U_afifo_U_acore_n90), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U59 (.ZN(U_afifo_U_acore_U_sub_fifo_n298), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1843_U_afifo_U_acore_U_sub_fifo_n126), 
	.A2(FE_PHN3257_U_afifo_U_acore_n104), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U58 (.ZN(U_afifo_U_acore_U_sub_fifo_n307), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1799_U_afifo_U_acore_U_sub_fifo_n135), 
	.A2(FE_PHN1844_U_afifo_U_acore_n201), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U57 (.ZN(U_afifo_U_acore_U_sub_fifo_n291), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n119), 
	.A2(FE_PHN1193_U_afifo_U_acore_n88), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U56 (.ZN(U_afifo_U_acore_U_sub_fifo_n314), 
	.B2(U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n141), 
	.A2(FE_PHN1408_U_afifo_U_acore_n173), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U55 (.ZN(U_afifo_U_acore_U_sub_fifo_n308), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1821_U_afifo_U_acore_U_sub_fifo_n136), 
	.A2(FE_PHN1839_U_afifo_U_acore_n203), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U54 (.ZN(U_afifo_U_acore_U_sub_fifo_n300), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1806_U_afifo_U_acore_U_sub_fifo_n128), 
	.A2(FE_PHN3384_U_afifo_U_acore_n156), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U53 (.ZN(U_afifo_U_acore_U_sub_fifo_n287), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1831_U_afifo_U_acore_U_sub_fifo_n115), 
	.A2(FE_PHN1552_U_afifo_U_acore_n80), 
	.A1(FE_OFN264_U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U52 (.ZN(U_afifo_U_acore_U_sub_fifo_n305), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1833_U_afifo_U_acore_U_sub_fifo_n133), 
	.A2(FE_PHN1835_U_afifo_U_acore_n197), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U51 (.ZN(U_afifo_U_acore_U_sub_fifo_n304), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n132), 
	.A2(FE_PHN1189_U_afifo_U_acore_n167), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U50 (.ZN(U_afifo_U_acore_U_sub_fifo_n288), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n116), 
	.A2(FE_PHN1187_U_afifo_U_acore_n82), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U49 (.ZN(U_afifo_U_acore_U_sub_fifo_n297), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1827_U_afifo_U_acore_U_sub_fifo_n125), 
	.A2(FE_PHN1837_U_afifo_U_acore_n102), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U48 (.ZN(U_afifo_U_acore_U_sub_fifo_n299), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1805_U_afifo_U_acore_U_sub_fifo_n127), 
	.A2(FE_PHN3409_U_afifo_U_acore_n153), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U47 (.ZN(U_afifo_U_acore_U_sub_fifo_n315), 
	.B2(U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n142), 
	.A2(FE_PHN1560_U_afifo_U_acore_n175), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U46 (.ZN(U_afifo_U_acore_U_sub_fifo_n274), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1816_U_afifo_U_acore_U_sub_fifo_n102), 
	.A2(FE_PHN1841_U_afifo_U_acore_n184), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U45 (.ZN(U_afifo_U_acore_U_sub_fifo_n294), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1822_U_afifo_U_acore_U_sub_fifo_n122), 
	.A2(FE_PHN1851_U_afifo_U_acore_n96), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U44 (.ZN(U_afifo_U_acore_U_sub_fifo_n311), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1820_U_afifo_U_acore_U_sub_fifo_n139), 
	.A2(U_afifo_U_acore_n31), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U43 (.ZN(U_afifo_U_acore_U_sub_fifo_n313), 
	.B2(U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1808_U_afifo_U_acore_U_sub_fifo_n140), 
	.A2(U_afifo_U_acore_n32), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U42 (.ZN(U_afifo_U_acore_U_sub_fifo_n302), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1828_U_afifo_U_acore_U_sub_fifo_n130), 
	.A2(FE_PHN3262_U_afifo_U_acore_n160), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U41 (.ZN(U_afifo_U_acore_U_sub_fifo_n310), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1814_U_afifo_U_acore_U_sub_fifo_n138), 
	.A2(FE_PHN1849_U_afifo_U_acore_n207), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U40 (.ZN(U_afifo_U_acore_U_sub_fifo_n295), 
	.B2(FE_OFN206_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1812_U_afifo_U_acore_U_sub_fifo_n123), 
	.A2(FE_PHN1850_U_afifo_U_acore_n98), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U39 (.ZN(U_afifo_U_acore_U_sub_fifo_n277), 
	.B2(U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(U_afifo_U_acore_U_sub_fifo_n105), 
	.A2(U_afifo_U_acore_n30), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   AOI22_X2 U_afifo_U_acore_U_sub_fifo_U38 (.ZN(U_afifo_U_acore_U_sub_fifo_n306), 
	.B2(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369), 
	.B1(FE_PHN1826_U_afifo_U_acore_U_sub_fifo_n134), 
	.A2(FE_PHN3243_U_afifo_U_acore_n199), 
	.A1(U_afifo_U_acore_U_sub_fifo_n152));
   NOR2_X2 U_afifo_U_acore_U_sub_fifo_U37 (.ZN(U_afifo_U_acore_U_sub_fifo_n160), 
	.A2(FE_PHN817_U_afifo_U_acore_n2), 
	.A1(U_afifo_U_acore_n166));
   OAI21_X2 U_afifo_U_acore_U_sub_fifo_U36 (.ZN(U_afifo_U_acore_U_sub_fifo_n171), 
	.B2(U_afifo_U_acore_U_sub_fifo_n163), 
	.B1(U_afifo_U_acore_U_sub_fifo_n160), 
	.A(U_afifo_U_acore_U_sub_fifo_n159));
   NAND2_X2 U_afifo_U_acore_U_sub_fifo_U35 (.ZN(U_afifo_U_acore_U_sub_fifo_n158), 
	.A2(U_afifo_U_acore_U_sub_fifo_n150), 
	.A1(U_afifo_U_acore_U_sub_fifo_n160));
   OAI21_X2 U_afifo_U_acore_U_sub_fifo_U34 (.ZN(U_afifo_U_acore_U_sub_fifo_n170), 
	.B2(U_afifo_U_acore_U_sub_fifo_n161), 
	.B1(U_afifo_U_acore_U_sub_fifo_n160), 
	.A(U_afifo_U_acore_U_sub_fifo_n158));
   OAI211_X1 U_afifo_U_acore_U_sub_fifo_U32 (.ZN(U_afifo_U_acore_U_sub_fifo_n172), 
	.C2(U_afifo_U_acore_U_sub_fifo_n166), 
	.C1(U_afifo_U_acore_n165), 
	.B(U_afifo_U_acore_m_sf_full), 
	.A(U_afifo_U_acore_U_sub_fifo_n165));
   INV_X8 U_afifo_U_acore_U_sub_fifo_U30 (.ZN(U_afifo_U_acore_U_sub_fifo_n153), 
	.A(FE_OFN6_U_afifo_U_acore_U_sub_fifo_n1));
   INV_X8 U_afifo_U_acore_U_sub_fifo_U28 (.ZN(U_afifo_U_acore_U_sub_fifo_n161), 
	.A(FE_PHN1592_U_afifo_U_acore_U_sub_fifo_out_ptr_0_));
   INV_X8 U_afifo_U_acore_U_sub_fifo_U27 (.ZN(U_afifo_U_acore_U_sub_fifo_n163), 
	.A(U_afifo_U_acore_U_sub_fifo_out_ptr_1_));
   INV_X8 U_afifo_U_acore_U_sub_fifo_U26 (.ZN(U_afifo_U_acore_U_sub_fifo_n212), 
	.A(FE_OFN4_U_afifo_U_acore_U_sub_fifo_n169));
   NAND2_X2 U_afifo_U_acore_U_sub_fifo_U25 (.ZN(U_afifo_U_acore_U_sub_fifo_n162), 
	.A2(U_afifo_U_acore_U_sub_fifo_n163), 
	.A1(U_afifo_U_acore_U_sub_fifo_n161));
   AND2_X4 U_afifo_U_acore_U_sub_fifo_U24 (.ZN(U_afifo_U_acore_n2), 
	.A2(U_afifo_U_acore_U_sub_fifo_n10), 
	.A1(U_afifo_U_acore_U_sub_fifo_n100));
   NAND2_X2 U_afifo_U_acore_U_sub_fifo_U23 (.ZN(U_afifo_U_acore_m_sf_full), 
	.A2(FE_PHN2979_U_afifo_U_acore_U_sub_fifo_count_0_), 
	.A1(FE_PHN867_U_afifo_U_acore_U_sub_fifo_count_1_));
   OAI21_X2 U_afifo_U_acore_U_sub_fifo_U22 (.ZN(U_afifo_U_acore_U_sub_fifo_n373), 
	.B2(U_afifo_U_acore_n163), 
	.B1(U_afifo_U_acore_m_sf_full), 
	.A(U_afifo_U_acore_U_sub_fifo_n167));
   NAND3_X1 U_afifo_U_acore_U_sub_fifo_U21 (.ZN(U_afifo_U_acore_U_sub_fifo_n159), 
	.A3(FE_PHN1592_U_afifo_U_acore_U_sub_fifo_out_ptr_0_), 
	.A2(U_afifo_U_acore_U_sub_fifo_n163), 
	.A1(U_afifo_U_acore_U_sub_fifo_n160));
   INV_X4 U_afifo_U_acore_U_sub_fifo_U20 (.ZN(U_afifo_U_acore_U_sub_fifo_n370), 
	.A(U_afifo_U_acore_U_sub_fifo_n373));
   XOR2_X1 U_afifo_U_acore_U_sub_fifo_U19 (.Z(U_afifo_U_acore_U_sub_fifo_n325), 
	.B(U_afifo_U_acore_U_sub_fifo_n372), 
	.A(U_afifo_U_acore_U_sub_fifo_n373));
   INV_X8 U_afifo_U_acore_U_sub_fifo_U4 (.ZN(U_afifo_U_acore_U_sub_fifo_n152), 
	.A(FE_OFN259_U_afifo_U_acore_U_sub_fifo_n369));
   OR3_X4 U_afifo_U_acore_U_sub_fifo_U3 (.ZN(U_afifo_U_acore_U_sub_fifo_n1), 
	.A3(FE_PHN993_U_afifo_U_acore_U_sub_fifo_n149), 
	.A2(U_afifo_U_acore_U_sub_fifo_n373), 
	.A1(U_afifo_U_acore_U_sub_fifo_in_ptr_1_));
   DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__0_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n50), 
	.D(FE_PHN1962_U_afifo_U_acore_U_sub_fifo_n272), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__2_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n49), 
	.D(FE_PHN1948_U_afifo_U_acore_U_sub_fifo_n270), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__3_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n48), 
	.D(FE_PHN1950_U_afifo_U_acore_U_sub_fifo_n269), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__4_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n47), 
	.D(FE_PHN1784_U_afifo_U_acore_U_sub_fifo_n268), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__5_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n9), 
	.D(FE_PHN1966_U_afifo_U_acore_U_sub_fifo_n267), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__6_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n46), 
	.D(FE_PHN1959_U_afifo_U_acore_U_sub_fifo_n266), 
	.CK(HCLK__L5_N36));
   DFFR_X2 U_afifo_U_acore_U_sub_fifo_in_ptr_reg_0_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n149), 
	.D(FE_PHN1635_U_afifo_U_acore_U_sub_fifo_n323), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_out_ptr_reg_0_ (.RN(FE_OFN57_HRESETn), 
	.Q(U_afifo_U_acore_U_sub_fifo_out_ptr_0_), 
	.D(U_afifo_U_acore_U_sub_fifo_n170), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_out_ptr_reg_1_ (.RN(FE_OFN47_HRESETn), 
	.Q(U_afifo_U_acore_U_sub_fifo_out_ptr_1_), 
	.D(FE_PHN1223_U_afifo_U_acore_U_sub_fifo_n171), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_count_reg_1_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n100), 
	.Q(U_afifo_U_acore_U_sub_fifo_count_1_), 
	.D(FE_PHN868_U_afifo_U_acore_U_sub_fifo_n172), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__49_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n101), 
	.D(FE_PHN2295_U_afifo_U_acore_U_sub_fifo_n173), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__48_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n51), 
	.D(FE_PHN2015_U_afifo_U_acore_U_sub_fifo_n174), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__47_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n52), 
	.D(FE_PHN2017_U_afifo_U_acore_U_sub_fifo_n175), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__46_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n62), 
	.D(FE_PHN2019_U_afifo_U_acore_U_sub_fifo_n176), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__45_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n63), 
	.D(FE_PHN2278_U_afifo_U_acore_U_sub_fifo_n177), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__44_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n53), 
	.D(FE_PHN2008_U_afifo_U_acore_U_sub_fifo_n178), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__43_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n64), 
	.D(FE_PHN2264_U_afifo_U_acore_U_sub_fifo_n179), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__42_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n65), 
	.D(FE_PHN2292_U_afifo_U_acore_U_sub_fifo_n180), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__41_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n66), 
	.D(FE_PHN2234_U_afifo_U_acore_U_sub_fifo_n181), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__40_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n67), 
	.D(FE_PHN2231_U_afifo_U_acore_U_sub_fifo_n182), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__39_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n68), 
	.D(FE_PHN2262_U_afifo_U_acore_U_sub_fifo_n183), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__38_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n69), 
	.D(FE_PHN1987_U_afifo_U_acore_U_sub_fifo_n184), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__37_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n54), 
	.D(FE_PHN2242_U_afifo_U_acore_U_sub_fifo_n185), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__36_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n70), 
	.D(FE_PHN2253_U_afifo_U_acore_U_sub_fifo_n186), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__35_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n71), 
	.D(FE_PHN1988_U_afifo_U_acore_U_sub_fifo_n187), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__34_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n72), 
	.D(FE_PHN1975_U_afifo_U_acore_U_sub_fifo_n188), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__33_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n73), 
	.D(FE_PHN2248_U_afifo_U_acore_U_sub_fifo_n189), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__32_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n55), 
	.D(FE_PHN2227_U_afifo_U_acore_U_sub_fifo_n190), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__31_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n74), 
	.D(FE_PHN2263_U_afifo_U_acore_U_sub_fifo_n191), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__30_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n75), 
	.D(FE_PHN2236_U_afifo_U_acore_U_sub_fifo_n192), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__29_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n76), 
	.D(FE_PHN2009_U_afifo_U_acore_U_sub_fifo_n193), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__28_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n77), 
	.D(FE_PHN2287_U_afifo_U_acore_U_sub_fifo_n194), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__27_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n78), 
	.D(FE_PHN2001_U_afifo_U_acore_U_sub_fifo_n195), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__26_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n79), 
	.D(FE_PHN2018_U_afifo_U_acore_U_sub_fifo_n196), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__25_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n56), 
	.D(FE_PHN2359_U_afifo_U_acore_U_sub_fifo_n197), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__24_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n80), 
	.D(FE_PHN2258_U_afifo_U_acore_U_sub_fifo_n198), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__23_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n81), 
	.D(FE_PHN2251_U_afifo_U_acore_U_sub_fifo_n199), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__22_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n82), 
	.D(FE_PHN2275_U_afifo_U_acore_U_sub_fifo_n200), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__21_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n83), 
	.D(FE_PHN2006_U_afifo_U_acore_U_sub_fifo_n201), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__20_ (.RN(FE_OFN150_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n84), 
	.D(FE_PHN2007_U_afifo_U_acore_U_sub_fifo_n202), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__19_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n85), 
	.D(FE_PHN2266_U_afifo_U_acore_U_sub_fifo_n203), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__18_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n57), 
	.D(FE_PHN2247_U_afifo_U_acore_U_sub_fifo_n204), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__17_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n86), 
	.D(FE_PHN2343_U_afifo_U_acore_U_sub_fifo_n205), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__16_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n87), 
	.D(FE_PHN1994_U_afifo_U_acore_U_sub_fifo_n206), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__15_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n88), 
	.D(FE_PHN2012_U_afifo_U_acore_U_sub_fifo_n207), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__14_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n89), 
	.D(FE_PHN2351_U_afifo_U_acore_U_sub_fifo_n208), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__13_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n58), 
	.D(FE_PHN1553_U_afifo_U_acore_U_sub_fifo_n209), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__12_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n90), 
	.D(FE_PHN2290_U_afifo_U_acore_U_sub_fifo_n210), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__11_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n91), 
	.D(FE_PHN2279_U_afifo_U_acore_U_sub_fifo_n211), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__9_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n92), 
	.D(FE_PHN2281_U_afifo_U_acore_U_sub_fifo_n213), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__8_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n93), 
	.D(FE_PHN1811_U_afifo_U_acore_U_sub_fifo_n214), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__7_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n94), 
	.D(FE_PHN2272_U_afifo_U_acore_U_sub_fifo_n215), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__6_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n95), 
	.D(FE_PHN1813_U_afifo_U_acore_U_sub_fifo_n216), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__5_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n59), 
	.D(FE_PHN1996_U_afifo_U_acore_U_sub_fifo_n217), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__4_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n96), 
	.D(FE_PHN2020_U_afifo_U_acore_U_sub_fifo_n218), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__3_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n97), 
	.D(FE_PHN1819_U_afifo_U_acore_U_sub_fifo_n219), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__2_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n98), 
	.D(FE_PHN1974_U_afifo_U_acore_U_sub_fifo_n220), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__0_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n99), 
	.D(FE_PHN1794_U_afifo_U_acore_U_sub_fifo_n222), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__49_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n12), 
	.D(FE_PHN2024_U_afifo_U_acore_U_sub_fifo_n223), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__48_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n60), 
	.D(FE_PHN2282_U_afifo_U_acore_U_sub_fifo_n224), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__47_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n61), 
	.D(FE_PHN1993_U_afifo_U_acore_U_sub_fifo_n225), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__46_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n13), 
	.D(FE_PHN2277_U_afifo_U_acore_U_sub_fifo_n226), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__45_ (.RN(FE_OFN169_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n14), 
	.D(FE_PHN2260_U_afifo_U_acore_U_sub_fifo_n227), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__44_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n3), 
	.D(FE_PHN2255_U_afifo_U_acore_U_sub_fifo_n228), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__43_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n15), 
	.D(FE_PHN1999_U_afifo_U_acore_U_sub_fifo_n229), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__42_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n16), 
	.D(FE_PHN2013_U_afifo_U_acore_U_sub_fifo_n230), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__41_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n17), 
	.D(FE_PHN2237_U_afifo_U_acore_U_sub_fifo_n231), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__40_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n18), 
	.D(FE_PHN2230_U_afifo_U_acore_U_sub_fifo_n232), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__39_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n19), 
	.D(FE_PHN1989_U_afifo_U_acore_U_sub_fifo_n233), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__38_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n20), 
	.D(FE_PHN2250_U_afifo_U_acore_U_sub_fifo_n234), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__37_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n4), 
	.D(FE_PHN2239_U_afifo_U_acore_U_sub_fifo_n235), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__36_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n21), 
	.D(FE_PHN1980_U_afifo_U_acore_U_sub_fifo_n236), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__35_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n22), 
	.D(FE_PHN2256_U_afifo_U_acore_U_sub_fifo_n237), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__34_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n23), 
	.D(FE_PHN1973_U_afifo_U_acore_U_sub_fifo_n238), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__33_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n24), 
	.D(FE_PHN1979_U_afifo_U_acore_U_sub_fifo_n239), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__32_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n5), 
	.D(FE_PHN1976_U_afifo_U_acore_U_sub_fifo_n240), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__31_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n25), 
	.D(FE_PHN2243_U_afifo_U_acore_U_sub_fifo_n241), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__30_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n26), 
	.D(FE_PHN1982_U_afifo_U_acore_U_sub_fifo_n242), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__29_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n27), 
	.D(FE_PHN2274_U_afifo_U_acore_U_sub_fifo_n243), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__28_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n28), 
	.D(FE_PHN2005_U_afifo_U_acore_U_sub_fifo_n244), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__27_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n29), 
	.D(FE_PHN2273_U_afifo_U_acore_U_sub_fifo_n245), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__26_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n30), 
	.D(FE_PHN2252_U_afifo_U_acore_U_sub_fifo_n246), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__25_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n6), 
	.D(FE_PHN2010_U_afifo_U_acore_U_sub_fifo_n247), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__24_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n31), 
	.D(FE_PHN2362_U_afifo_U_acore_U_sub_fifo_n248), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__23_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n32), 
	.D(FE_PHN2267_U_afifo_U_acore_U_sub_fifo_n249), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__22_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n33), 
	.D(FE_PHN2021_U_afifo_U_acore_U_sub_fifo_n250), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__21_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n34), 
	.D(FE_PHN1995_U_afifo_U_acore_U_sub_fifo_n251), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__20_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n35), 
	.D(FE_PHN2269_U_afifo_U_acore_U_sub_fifo_n252), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__19_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n36), 
	.D(FE_PHN2276_U_afifo_U_acore_U_sub_fifo_n253), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__18_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n7), 
	.D(FE_PHN2246_U_afifo_U_acore_U_sub_fifo_n254), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__17_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n37), 
	.D(FE_PHN1986_U_afifo_U_acore_U_sub_fifo_n255), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__16_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n38), 
	.D(FE_PHN2268_U_afifo_U_acore_U_sub_fifo_n256), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__15_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n39), 
	.D(FE_PHN2321_U_afifo_U_acore_U_sub_fifo_n257), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__14_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n40), 
	.D(FE_PHN2249_U_afifo_U_acore_U_sub_fifo_n258), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__13_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n8), 
	.D(FE_PHN2308_U_afifo_U_acore_U_sub_fifo_n259), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__12_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n41), 
	.D(FE_PHN1991_U_afifo_U_acore_U_sub_fifo_n260), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__11_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n42), 
	.D(FE_PHN2011_U_afifo_U_acore_U_sub_fifo_n261), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__9_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n43), 
	.D(FE_PHN2000_U_afifo_U_acore_U_sub_fifo_n263), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__8_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n44), 
	.D(FE_PHN1823_U_afifo_U_acore_U_sub_fifo_n264), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__7_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n45), 
	.D(FE_PHN2324_U_afifo_U_acore_U_sub_fifo_n265), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__49_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n2), 
	.D(FE_PHN1829_U_afifo_U_acore_U_sub_fifo_n273), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__48_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n102), 
	.D(FE_PHN5038_U_afifo_U_acore_U_sub_fifo_n274), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__47_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n103), 
	.D(FE_PHN2022_U_afifo_U_acore_U_sub_fifo_n275), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__46_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n104), 
	.D(FE_PHN2244_U_afifo_U_acore_U_sub_fifo_n276), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__45_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n105), 
	.D(FE_PHN1803_U_afifo_U_acore_U_sub_fifo_n277), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__44_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n106), 
	.D(FE_PHN3173_U_afifo_U_acore_U_sub_fifo_n278), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__43_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n107), 
	.D(FE_PHN2315_U_afifo_U_acore_U_sub_fifo_n279), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__42_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n108), 
	.D(FE_PHN3159_U_afifo_U_acore_U_sub_fifo_n280), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__41_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n109), 
	.D(FE_PHN1981_U_afifo_U_acore_U_sub_fifo_n281), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__40_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n110), 
	.D(FE_PHN1971_U_afifo_U_acore_U_sub_fifo_n282), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__39_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n111), 
	.D(FE_PHN2261_U_afifo_U_acore_U_sub_fifo_n283), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__38_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n112), 
	.D(FE_PHN2257_U_afifo_U_acore_U_sub_fifo_n284), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__37_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n113), 
	.D(FE_PHN1985_U_afifo_U_acore_U_sub_fifo_n285), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__36_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n114), 
	.D(FE_PHN2238_U_afifo_U_acore_U_sub_fifo_n286), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__35_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n115), 
	.D(FE_PHN3184_U_afifo_U_acore_U_sub_fifo_n287), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__34_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n116), 
	.D(FE_PHN2226_U_afifo_U_acore_U_sub_fifo_n288), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__33_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n117), 
	.D(FE_PHN2259_U_afifo_U_acore_U_sub_fifo_n289), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__32_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n118), 
	.D(FE_PHN2228_U_afifo_U_acore_U_sub_fifo_n290), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__31_ (.RN(FE_OFN29_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n119), 
	.D(FE_PHN1984_U_afifo_U_acore_U_sub_fifo_n291), 
	.CK(HCLK__L5_N39));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__30_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n120), 
	.D(FE_PHN3178_U_afifo_U_acore_U_sub_fifo_n292), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__29_ (.RN(FE_OFN32_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n121), 
	.D(FE_PHN2003_U_afifo_U_acore_U_sub_fifo_n293), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__28_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n122), 
	.D(FE_PHN5152_U_afifo_U_acore_U_sub_fifo_n294), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__27_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n123), 
	.D(FE_PHN3161_U_afifo_U_acore_U_sub_fifo_n295), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__26_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n124), 
	.D(FE_PHN4789_U_afifo_U_acore_U_sub_fifo_n296), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__25_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n125), 
	.D(FE_PHN4677_U_afifo_U_acore_U_sub_fifo_n297), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__24_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n126), 
	.D(FE_PHN2026_U_afifo_U_acore_U_sub_fifo_n298), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__23_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n127), 
	.D(FE_PHN1998_U_afifo_U_acore_U_sub_fifo_n299), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__22_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n128), 
	.D(FE_PHN2271_U_afifo_U_acore_U_sub_fifo_n300), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__21_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n129), 
	.D(FE_PHN2328_U_afifo_U_acore_U_sub_fifo_n301), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__20_ (.RN(FE_OFN149_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n130), 
	.D(FE_PHN2316_U_afifo_U_acore_U_sub_fifo_n302), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__19_ (.RN(FE_OFN58_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n131), 
	.D(FE_PHN1992_U_afifo_U_acore_U_sub_fifo_n303), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__18_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n132), 
	.D(FE_PHN1977_U_afifo_U_acore_U_sub_fifo_n304), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__17_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n133), 
	.D(FE_PHN3179_U_afifo_U_acore_U_sub_fifo_n305), 
	.CK(HCLK__L5_N37));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__16_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n134), 
	.D(FE_PHN2312_U_afifo_U_acore_U_sub_fifo_n306), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__15_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n135), 
	.D(FE_PHN5067_U_afifo_U_acore_U_sub_fifo_n307), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__14_ (.RN(FE_OFN47_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n136), 
	.D(FE_PHN5103_U_afifo_U_acore_U_sub_fifo_n308), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__13_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n137), 
	.D(FE_PHN2014_U_afifo_U_acore_U_sub_fifo_n309), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__12_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n138), 
	.D(FE_PHN3177_U_afifo_U_acore_U_sub_fifo_n310), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__11_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n139), 
	.D(FE_PHN2016_U_afifo_U_acore_U_sub_fifo_n311), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__9_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n140), 
	.D(FE_PHN2002_U_afifo_U_acore_U_sub_fifo_n313), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__8_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n141), 
	.D(FE_PHN1824_U_afifo_U_acore_U_sub_fifo_n314), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__7_ (.RN(FE_OFN168_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n142), 
	.D(FE_PHN1474_U_afifo_U_acore_U_sub_fifo_n315), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__6_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n143), 
	.D(FE_PHN5162_U_afifo_U_acore_U_sub_fifo_n316), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__5_ (.RN(FE_OFN170_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n144), 
	.D(FE_PHN1807_U_afifo_U_acore_U_sub_fifo_n317), 
	.CK(HCLK__L5_N38));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__4_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n145), 
	.D(FE_PHN3158_U_afifo_U_acore_U_sub_fifo_n318), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__3_ (.RN(FE_OFN34_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n146), 
	.D(FE_PHN2265_U_afifo_U_acore_U_sub_fifo_n319), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__2_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n147), 
	.D(FE_PHN1972_U_afifo_U_acore_U_sub_fifo_n320), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__0_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n148), 
	.D(FE_PHN3181_U_afifo_U_acore_U_sub_fifo_n322), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_in_ptr_reg_1_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n11), 
	.Q(U_afifo_U_acore_U_sub_fifo_in_ptr_1_), 
	.D(FE_PHN1471_U_afifo_U_acore_U_sub_fifo_n324), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_afifo_U_acore_U_sub_fifo_count_reg_0_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_afifo_U_acore_U_sub_fifo_n10), 
	.Q(U_afifo_U_acore_U_sub_fifo_count_0_), 
	.D(FE_PHN1100_U_afifo_U_acore_U_sub_fifo_n325), 
	.CK(HCLK__L5_N36));
   OAI21_X1 U_dfifo_U_dcore_U_sub_fifo_U435 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n448), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n57), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n603), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n12));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U434 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n310), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n117), 
	.A2(n60), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U433 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n309), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n116), 
	.A2(n59), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U432 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n308), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n115), 
	.A2(n52), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U431 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n307), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n114), 
	.A2(n58), 
	.A1(FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U430 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n306), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n113), 
	.A2(n57), 
	.A1(FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U429 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n305), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n112), 
	.A2(n56), 
	.A1(FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U428 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n304), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n111), 
	.A2(n55), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U427 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n303), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n110), 
	.A2(n54), 
	.A1(FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U426 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n302), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n109), 
	.A2(n53), 
	.A1(FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U425 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n301), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n108), 
	.A2(n67), 
	.A1(FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U424 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n300), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n107), 
	.A2(n66), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U423 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n299), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n106), 
	.A2(n65), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U422 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n298), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n105), 
	.A2(n64), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U421 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n297), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n104), 
	.A2(n63), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U420 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n296), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n103), 
	.A2(n62), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U419 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n295), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n102), 
	.A2(n61), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U418 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n294), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n101), 
	.A2(n83), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U417 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n293), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n100), 
	.A2(n82), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U416 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n292), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n99), 
	.A2(n81), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U415 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n291), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n98), 
	.A2(n80), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U414 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n290), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n97), 
	.A2(n79), 
	.A1(FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U413 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n289), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n96), 
	.A2(n78), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U412 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n288), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n95), 
	.A2(n77), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U411 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n287), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n94), 
	.A2(n76), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U410 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n286), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n93), 
	.A2(n75), 
	.A1(FE_OFN280_U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U409 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n285), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n92), 
	.A2(n74), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U408 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n284), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n91), 
	.A2(n85), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U407 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n283), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n90), 
	.A2(n84), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U406 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n282), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n89), 
	.A2(n73), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U405 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n281), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n88), 
	.A2(n72), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U404 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n280), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n87), 
	.A2(n71), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U403 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n279), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n86), 
	.A2(n70), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U402 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n276), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n52), 
	.A2(n60), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U401 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n275), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n51), 
	.A2(n59), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U400 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n274), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n50), 
	.A2(n52), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U399 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n273), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n49), 
	.A2(n58), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U398 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n272), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n48), 
	.A2(n57), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U397 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n271), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n47), 
	.A2(n56), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U396 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n270), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n46), 
	.A2(n55), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U395 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n269), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n45), 
	.A2(n54), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U394 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n268), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n44), 
	.A2(n53), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U393 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n267), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n43), 
	.A2(n67), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U392 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n266), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n42), 
	.A2(n66), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U391 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n265), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n41), 
	.A2(n65), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U390 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n264), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n40), 
	.A2(n64), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U389 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n263), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n39), 
	.A2(n63), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U388 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n262), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n38), 
	.A2(n62), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U387 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n261), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n37), 
	.A2(n61), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U386 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n260), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n36), 
	.A2(n83), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U385 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n259), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n35), 
	.A2(n82), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U384 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n258), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n34), 
	.A2(n81), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U383 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n257), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n33), 
	.A2(n80), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U382 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n256), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n32), 
	.A2(n79), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U381 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n255), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n31), 
	.A2(n78), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U380 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n254), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n30), 
	.A2(n77), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U379 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n253), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n29), 
	.A2(n76), 
	.A1(FE_OFN281_U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U378 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n252), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n28), 
	.A2(n75), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U377 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n251), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n27), 
	.A2(n74), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U376 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n250), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n26), 
	.A2(n85), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U375 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n249), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n25), 
	.A2(n84), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U374 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n248), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n24), 
	.A2(n73), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U373 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n247), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n23), 
	.A2(n72), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U372 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n246), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n22), 
	.A2(n71), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U371 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n245), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n21), 
	.A2(n70), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   OR2_X4 U_dfifo_U_dcore_U_sub_fifo_U370 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n567), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n602));
   OR2_X4 U_dfifo_U_dcore_U_sub_fifo_U369 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n567), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n604));
   OR3_X4 U_dfifo_U_dcore_U_sub_fifo_U368 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.A3(U_dfifo_U_dcore_U_sub_fifo_n602), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_in_ptr_2_));
   OR3_X4 U_dfifo_U_dcore_U_sub_fifo_U367 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.A3(U_dfifo_U_dcore_U_sub_fifo_n604), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_in_ptr_2_));
   AND2_X4 U_dfifo_U_dcore_U_sub_fifo_U366 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n18), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n460));
   AOI21_X1 U_dfifo_U_dcore_U_sub_fifo_U365 (.ZN(U_dfifo_U_dcore_m_sf_afull), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n54), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n13), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n17));
   INV_X1 U_dfifo_U_dcore_U_sub_fifo_U364 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n603), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n602));
   NOR3_X1 U_dfifo_U_dcore_U_sub_fifo_U363 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n456), 
	.A3(U_dfifo_U_dcore_U_sub_fifo_n13), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n609), 
	.A1(U_dfifo_U_dcore_n208));
   OAI21_X1 U_dfifo_U_dcore_U_sub_fifo_U362 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n449), 
	.B2(FE_PHN1791_U_dfifo_U_dcore_U_sub_fifo_n55), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n458), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n604));
   NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U359 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n460), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_out_ptr_1_));
   NOR2_X4 U_dfifo_U_dcore_U_sub_fifo_U358 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n56), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_));
   NOR2_X4 U_dfifo_U_dcore_U_sub_fifo_U357 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n56), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n18));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U356 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n514), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__25_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__25_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U355 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n512), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n92), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n27));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U354 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n513), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__25_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n512));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U353 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n490), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__18_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__18_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U352 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n488), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n99), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n34));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U351 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n489), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__18_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n488));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U350 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n466), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__10_), 
	.A2(FE_OFN271_U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__10_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U349 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n464), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n107), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n42));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U348 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n465), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__10_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n464));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U347 (.ZN(U_dfifo_U_dcore_m_sf_data_out[10]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1782_U_dfifo_U_dcore_U_sub_fifo_n73), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n465), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n466));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U346 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n487), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__17_), 
	.A2(FE_OFN271_U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__17_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U345 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n485), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n100), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n35));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U344 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n486), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__17_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n485));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U343 (.ZN(U_dfifo_U_dcore_m_sf_data_out[17]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1765_U_dfifo_U_dcore_U_sub_fifo_n66), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n486), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n487));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U342 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n564), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__9_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__9_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U341 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n561), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n108), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n43));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U340 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n563), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__9_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n561));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U339 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n529), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__2_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__2_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U338 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n527), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n115), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n50));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U337 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n528), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__2_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n527));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U336 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n511), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__24_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__24_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U335 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n509), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n93), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n28));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U334 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n510), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__24_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n509));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U333 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n478), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__14_), 
	.A2(FE_OFN271_U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__14_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U332 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n476), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n103), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n38));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U331 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n477), 
	.B2(FE_OFN267_U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__14_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n476));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U330 (.ZN(U_dfifo_U_dcore_m_sf_data_out[14]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1781_U_dfifo_U_dcore_U_sub_fifo_n69), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n477), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n478));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U329 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n469), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__11_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__11_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U328 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n467), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n106), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n41));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U327 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n468), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__11_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n467));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U326 (.ZN(U_dfifo_U_dcore_m_sf_data_out[11]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1772_U_dfifo_U_dcore_U_sub_fifo_n72), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n468), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n469));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U325 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n475), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__13_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__13_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U324 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n473), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n104), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n39));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U323 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n474), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__13_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n473));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U322 (.ZN(U_dfifo_U_dcore_m_sf_data_out[13]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1775_U_dfifo_U_dcore_U_sub_fifo_n70), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n474), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n475));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U321 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n472), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__12_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__12_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U320 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n470), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n105), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n40));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U319 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n471), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__12_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n470));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U318 (.ZN(U_dfifo_U_dcore_m_sf_data_out[12]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1776_U_dfifo_U_dcore_U_sub_fifo_n71), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n471), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n472));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U317 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n541), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__33_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__33_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U316 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n539), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n84), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n19));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U315 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n540), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__33_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n539));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U314 (.ZN(U_dfifo_U_dcore_m_sf_data_out[33]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1767_U_dfifo_U_dcore_U_sub_fifo_n58), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n540), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n541));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U313 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n517), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__26_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__26_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U312 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n515), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n91), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n26));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U311 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n516), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__26_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n515));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U310 (.ZN(U_dfifo_U_dcore_m_sf_data_out[26]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1778_U_dfifo_U_dcore_U_sub_fifo_n65), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n516), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n517));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U309 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n508), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__23_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__23_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U308 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n506), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n94), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n29));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U307 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n507), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__23_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n506));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U306 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n484), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__16_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__16_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U305 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n482), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n101), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n36));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U304 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n483), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__16_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n482));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U303 (.ZN(U_dfifo_U_dcore_m_sf_data_out[16]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1764_U_dfifo_U_dcore_U_sub_fifo_n67), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n483), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n484));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U302 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n481), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__15_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__15_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U301 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n479), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n102), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n37));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U300 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n480), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__15_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n479));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U299 (.ZN(U_dfifo_U_dcore_m_sf_data_out[15]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1766_U_dfifo_U_dcore_U_sub_fifo_n68), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n480), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n481));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U298 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n499), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__20_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__20_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U297 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n497), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n97), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n32));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U296 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n498), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__20_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n497));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U295 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n493), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__19_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__19_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U294 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n491), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n98), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n33));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U293 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n492), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__19_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n491));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U292 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n505), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__22_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__22_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U291 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n503), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n95), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n30));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U290 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n504), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__22_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n503));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U289 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n502), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__21_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__21_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U288 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n500), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n96), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n31));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U287 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n501), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__21_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n500));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U286 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n559), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__8_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__8_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U285 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n557), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n109), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n44));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U284 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n558), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__8_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n557));
   NAND2_X2 U_dfifo_U_dcore_U_sub_fifo_U282 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n604), 
	.A2(FE_PHN1791_U_dfifo_U_dcore_U_sub_fifo_n55), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n458));
   NAND2_X2 U_dfifo_U_dcore_U_sub_fifo_U249 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n602), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_in_ptr_0_), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n458));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U248 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n550), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__5_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__5_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U247 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n548), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n112), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n47));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U246 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n549), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__5_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n548));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U245 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n547), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__4_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__4_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U244 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n545), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n113), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n48));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U243 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n546), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__4_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n545));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U242 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n556), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__7_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__7_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U241 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n554), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n110), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n45));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U240 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n555), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__7_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n554));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U239 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n553), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__6_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__6_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U238 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n551), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n111), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n46));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U237 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n552), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__6_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n551));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U236 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n544), 
	.B2(FE_OFN265_U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__3_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__3_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U235 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n542), 
	.B2(FE_OFN282_U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n114), 
	.A2(FE_OFN289_U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n49));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U234 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n543), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__3_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n542));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U233 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n535), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__31_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__31_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U232 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n533), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n86), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n21));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U231 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n534), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__31_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n533));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U230 (.ZN(U_dfifo_U_dcore_m_sf_data_out[31]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1771_U_dfifo_U_dcore_U_sub_fifo_n60), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n534), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n535));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U229 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n538), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__32_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__32_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U228 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n536), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n85), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n20));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U227 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n537), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__32_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n536));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U226 (.ZN(U_dfifo_U_dcore_m_sf_data_out[32]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1774_U_dfifo_U_dcore_U_sub_fifo_n59), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n537), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n538));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U225 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n463), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__0_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__0_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U224 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n461), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n117), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n52));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U223 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n462), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__0_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n461));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U222 (.ZN(U_dfifo_U_dcore_m_sf_data_out[0]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1556_U_dfifo_U_dcore_U_sub_fifo_n83), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n462), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n463));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U221 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n364), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1781_U_dfifo_U_dcore_U_sub_fifo_n69), 
	.A2(n62), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U220 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n375), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1802_U_dfifo_U_dcore_U_sub_fifo_n80), 
	.A2(n58), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U219 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n361), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1765_U_dfifo_U_dcore_U_sub_fifo_n66), 
	.A2(n82), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U218 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n362), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1764_U_dfifo_U_dcore_U_sub_fifo_n67), 
	.A2(n83), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U217 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n347), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1771_U_dfifo_U_dcore_U_sub_fifo_n60), 
	.A2(n70), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U216 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n355), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1543_U_dfifo_U_dcore_U_sub_fifo_n120), 
	.A2(n76), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U215 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n373), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1779_U_dfifo_U_dcore_U_sub_fifo_n78), 
	.A2(n56), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U214 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n353), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1541_U_dfifo_U_dcore_U_sub_fifo_n118), 
	.A2(n74), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U213 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n359), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1540_U_dfifo_U_dcore_U_sub_fifo_n124), 
	.A2(n80), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U212 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n350), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1787_U_dfifo_U_dcore_U_sub_fifo_n63), 
	.A2(n73), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U211 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n349), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1785_U_dfifo_U_dcore_U_sub_fifo_n62), 
	.A2(n72), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U210 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n363), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1766_U_dfifo_U_dcore_U_sub_fifo_n68), 
	.A2(n61), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U209 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n345), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1767_U_dfifo_U_dcore_U_sub_fifo_n58), 
	.A2(n69), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U208 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n346), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1774_U_dfifo_U_dcore_U_sub_fifo_n59), 
	.A2(n68), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U207 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n368), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1782_U_dfifo_U_dcore_U_sub_fifo_n73), 
	.A2(n66), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U206 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n374), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1790_U_dfifo_U_dcore_U_sub_fifo_n79), 
	.A2(n57), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U205 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n371), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1760_U_dfifo_U_dcore_U_sub_fifo_n76), 
	.A2(n54), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U204 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n352), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1778_U_dfifo_U_dcore_U_sub_fifo_n65), 
	.A2(n85), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U203 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n376), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1788_U_dfifo_U_dcore_U_sub_fifo_n81), 
	.A2(n52), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U202 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n366), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1776_U_dfifo_U_dcore_U_sub_fifo_n71), 
	.A2(n64), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U201 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n351), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1773_U_dfifo_U_dcore_U_sub_fifo_n64), 
	.A2(n84), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U200 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n348), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1768_U_dfifo_U_dcore_U_sub_fifo_n61), 
	.A2(n71), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U199 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n365), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1775_U_dfifo_U_dcore_U_sub_fifo_n70), 
	.A2(n63), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U198 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n367), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1772_U_dfifo_U_dcore_U_sub_fifo_n72), 
	.A2(n65), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U197 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n356), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n121), 
	.A2(n77), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U196 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n372), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1753_U_dfifo_U_dcore_U_sub_fifo_n77), 
	.A2(n55), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U195 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n369), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1755_U_dfifo_U_dcore_U_sub_fifo_n74), 
	.A2(n67), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U194 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n377), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1795_U_dfifo_U_dcore_U_sub_fifo_n82), 
	.A2(n59), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U193 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n360), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1546_U_dfifo_U_dcore_U_sub_fifo_n125), 
	.A2(n81), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U192 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n354), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1539_U_dfifo_U_dcore_U_sub_fifo_n119), 
	.A2(n75), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U191 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n378), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1556_U_dfifo_U_dcore_U_sub_fifo_n83), 
	.A2(n60), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U190 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n357), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1542_U_dfifo_U_dcore_U_sub_fifo_n122), 
	.A2(n78), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U189 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n370), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1754_U_dfifo_U_dcore_U_sub_fifo_n75), 
	.A2(n53), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U188 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n358), 
	.B2(FE_OFN286_U_dfifo_U_dcore_U_sub_fifo_n10), 
	.B1(FE_PHN1545_U_dfifo_U_dcore_U_sub_fifo_n123), 
	.A2(n79), 
	.A1(FE_OFN275_U_dfifo_U_dcore_U_sub_fifo_n232));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U187 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n333), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n150), 
	.A2(n65), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U186 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n319), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n136), 
	.A2(n74), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U185 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n326), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n143), 
	.A2(n81), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U184 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n322), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n139), 
	.A2(n77), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U183 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n321), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n138), 
	.A2(n76), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U182 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n334), 
	.B2(FE_OFN288_U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n151), 
	.A2(n66), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U181 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n331), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n148), 
	.A2(n63), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U180 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n318), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n135), 
	.A2(n85), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U179 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n332), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n149), 
	.A2(FE_OFN296_n64), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U178 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n328), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n145), 
	.A2(n83), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U177 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n324), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n141), 
	.A2(n79), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U176 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n317), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n134), 
	.A2(n84), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U175 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n335), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n152), 
	.A2(n67), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U174 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n314), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n131), 
	.A2(n71), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U173 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n330), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n147), 
	.A2(n62), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U172 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n336), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n153), 
	.A2(FE_OFN290_n53), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U171 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n327), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n144), 
	.A2(n82), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U170 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n320), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n137), 
	.A2(n75), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U169 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n337), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n154), 
	.A2(n54), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U168 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n312), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n129), 
	.A2(n68), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U167 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n338), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n155), 
	.A2(FE_OFN291_n55), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U166 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n313), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n130), 
	.A2(n70), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U165 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n325), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n142), 
	.A2(n80), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U164 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n339), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n156), 
	.A2(FE_OFN292_n56), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U163 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n311), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n128), 
	.A2(n69), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U162 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n315), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n132), 
	.A2(n72), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U161 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n323), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n140), 
	.A2(n78), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U160 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n340), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n157), 
	.A2(n57), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U159 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n329), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n146), 
	.A2(FE_OFN295_n61), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U158 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n316), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n133), 
	.A2(n73), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U157 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n341), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n158), 
	.A2(n58), 
	.A1(FE_OFN278_U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U156 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n343), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n160), 
	.A2(n59), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U155 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n344), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n161), 
	.A2(FE_OFN294_n60), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U154 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n342), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n159), 
	.A2(n52), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n231));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U153 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n523), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__28_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__28_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U152 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n521), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n89), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n24));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U151 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n522), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__28_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n521));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U150 (.ZN(U_dfifo_U_dcore_m_sf_data_out[28]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1787_U_dfifo_U_dcore_U_sub_fifo_n63), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n522), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n523));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U149 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n520), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__27_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__27_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U148 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n518), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n90), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n25));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U147 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n519), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__27_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n518));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U146 (.ZN(U_dfifo_U_dcore_m_sf_data_out[27]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1773_U_dfifo_U_dcore_U_sub_fifo_n64), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n519), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n520));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U145 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n526), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__29_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__29_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U144 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n524), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n88), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n23));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U143 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n525), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__29_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n524));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U142 (.ZN(U_dfifo_U_dcore_m_sf_data_out[29]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1785_U_dfifo_U_dcore_U_sub_fifo_n62), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n525), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n526));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U141 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n532), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__30_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__30_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U140 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n530), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n87), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n22));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U139 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n531), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__30_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n530));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U138 (.ZN(U_dfifo_U_dcore_m_sf_data_out[30]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1768_U_dfifo_U_dcore_U_sub_fifo_n61), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n531), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n532));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U137 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n441), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n224), 
	.A2(n56), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U136 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n414), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n197), 
	.A2(n68), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U135 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n413), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n196), 
	.A2(n69), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U134 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n416), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n199), 
	.A2(n71), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U133 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n445), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n228), 
	.A2(n59), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U132 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n418), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n201), 
	.A2(n73), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U131 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n417), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n200), 
	.A2(n72), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U130 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n438), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n221), 
	.A2(n53), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U129 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n415), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n198), 
	.A2(n70), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U128 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n446), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n229), 
	.A2(n60), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U127 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n442), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n225), 
	.A2(n57), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U126 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n444), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n227), 
	.A2(n52), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U125 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n440), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n223), 
	.A2(n55), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U124 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n439), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n222), 
	.A2(n54), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U123 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n443), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n226), 
	.A2(n58), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U122 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n399), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n182), 
	.A2(n63), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U121 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n402), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n185), 
	.A2(n66), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U120 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n407), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n190), 
	.A2(n56), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U119 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n397), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n180), 
	.A2(n61), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U118 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n406), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n189), 
	.A2(n55), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U117 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n412), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n195), 
	.A2(n60), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U116 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n405), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n188), 
	.A2(n54), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U115 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n398), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n181), 
	.A2(n62), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U114 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n400), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n183), 
	.A2(n64), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U113 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n408), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n191), 
	.A2(n57), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U112 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n401), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n184), 
	.A2(n65), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U111 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n409), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n192), 
	.A2(n58), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U110 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n404), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n187), 
	.A2(n53), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U109 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n403), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n186), 
	.A2(n67), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U108 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n411), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n194), 
	.A2(n59), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U107 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n410), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n193), 
	.A2(n52), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U106 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n496), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_3__1_), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n560), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_mem_2__1_));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U105 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n494), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n116), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n51));
   AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U104 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n495), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n562), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_mem_0__1_), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n494));
   OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U103 (.ZN(U_dfifo_U_dcore_m_sf_data_out[1]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1795_U_dfifo_U_dcore_U_sub_fifo_n82), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n495), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n496));
   NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U102 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n607), 
	.A2(FE_PHN1584_U_dfifo_U_dcore_U_sub_fifo_n18), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n608));
   OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U101 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n451), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n608), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n56), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n607));
   OAI21_X2 U_dfifo_U_dcore_U_sub_fifo_U100 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n452), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n126), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n607), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n606));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U98 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n278), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n85), 
	.A2(n68), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U97 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n277), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n84), 
	.A2(n69), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n16));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U96 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n243), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n19), 
	.A2(n69), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U95 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n244), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n20), 
	.A2(n68), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n15));
   NAND2_X1 U_dfifo_U_dcore_U_sub_fifo_U94 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n567), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n57), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_));
   INV_X1 U_dfifo_U_dcore_U_sub_fifo_U93 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n608), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n609));
   NAND3_X1 U_dfifo_U_dcore_U_sub_fifo_U92 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n606), 
	.A3(U_dfifo_U_dcore_U_sub_fifo_n126), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n605), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n609));
   NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U88 (.ZN(U_dfifo_U_dcore_m_sf_full), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n17), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n241));
   NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U87 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n455), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n609), 
	.A1(U_dfifo_U_dcore_n24));
   NOR3_X4 U_dfifo_U_dcore_U_sub_fifo_U86 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n16), 
	.A3(U_dfifo_U_dcore_U_sub_fifo_n604), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n57), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_));
   NOR3_X4 U_dfifo_U_dcore_U_sub_fifo_U85 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n15), 
	.A3(U_dfifo_U_dcore_U_sub_fifo_n602), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n57), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_));
   INV_X4 U_dfifo_U_dcore_U_sub_fifo_U84 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n234), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n12));
   INV_X4 U_dfifo_U_dcore_U_sub_fifo_U83 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n233), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n11));
   NAND2_X2 U_dfifo_U_dcore_U_sub_fifo_U82 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n241), 
	.A2(FE_PHN1422_U_dfifo_U_dcore_U_sub_fifo_count_1_), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n13));
   NAND2_X4 U_dfifo_U_dcore_U_sub_fifo_U81 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n460), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_));
   NAND2_X4 U_dfifo_U_dcore_U_sub_fifo_U80 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n14), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n18), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_));
   NAND2_X4 U_dfifo_U_dcore_U_sub_fifo_U79 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n8), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U76 (.ZN(U_dfifo_U_dcore_m_sf_data_out[23]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1543_U_dfifo_U_dcore_U_sub_fifo_n120), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n507), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n508));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U75 (.ZN(U_dfifo_U_dcore_m_sf_data_out[22]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(U_dfifo_U_dcore_U_sub_fifo_n121), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n504), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n505));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U74 (.ZN(U_dfifo_U_dcore_m_sf_data_out[21]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1542_U_dfifo_U_dcore_U_sub_fifo_n122), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n501), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n502));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U73 (.ZN(U_dfifo_U_dcore_m_sf_data_out[20]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1545_U_dfifo_U_dcore_U_sub_fifo_n123), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n498), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n499));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U72 (.ZN(U_dfifo_U_dcore_m_sf_data_out[8]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1754_U_dfifo_U_dcore_U_sub_fifo_n75), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n558), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n559));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U71 (.ZN(U_dfifo_U_dcore_m_sf_data_out[5]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1779_U_dfifo_U_dcore_U_sub_fifo_n78), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n549), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n550));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U70 (.ZN(U_dfifo_U_dcore_m_sf_data_out[6]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1753_U_dfifo_U_dcore_U_sub_fifo_n77), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n552), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n553));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U69 (.ZN(U_dfifo_U_dcore_m_sf_data_out[4]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1790_U_dfifo_U_dcore_U_sub_fifo_n79), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n546), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n547));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U68 (.ZN(U_dfifo_U_dcore_m_sf_data_out[7]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1760_U_dfifo_U_dcore_U_sub_fifo_n76), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n555), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n556));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U67 (.ZN(U_dfifo_U_dcore_m_sf_data_out[3]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1802_U_dfifo_U_dcore_U_sub_fifo_n80), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n543), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n544));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U66 (.ZN(U_dfifo_U_dcore_m_sf_data_out[9]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1755_U_dfifo_U_dcore_U_sub_fifo_n74), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n563), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n564));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U65 (.ZN(U_dfifo_U_dcore_m_sf_data_out[24]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1539_U_dfifo_U_dcore_U_sub_fifo_n119), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n510), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n511));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U64 (.ZN(U_dfifo_U_dcore_m_sf_data_out[2]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1788_U_dfifo_U_dcore_U_sub_fifo_n81), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n528), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n529));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U63 (.ZN(U_dfifo_U_dcore_m_sf_data_out[25]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1541_U_dfifo_U_dcore_U_sub_fifo_n118), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n513), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n514));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U62 (.ZN(U_dfifo_U_dcore_m_sf_data_out[18]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1546_U_dfifo_U_dcore_U_sub_fifo_n125), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n489), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n490));
   OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U61 (.ZN(U_dfifo_U_dcore_m_sf_data_out[19]), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
	.C1(FE_PHN1540_U_dfifo_U_dcore_U_sub_fifo_n124), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n492), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n493));
   NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U60 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n609), 
	.A2(U_dfifo_U_dcore_m_sf_empty), 
	.A1(U_dfifo_U_dcore_n209));
   NOR2_X1 U_dfifo_U_dcore_U_sub_fifo_U59 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n565), 
	.A2(FE_PHN1595_U_dfifo_U_dcore_U_sub_fifo_count_0_), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n608));
   NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U58 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n458), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n455), 
	.A1(U_dfifo_U_dcore_n208));
   AOI21_X1 U_dfifo_U_dcore_U_sub_fifo_U57 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n453), 
	.B2(FE_PHN1584_U_dfifo_U_dcore_U_sub_fifo_n18), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n608), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n607));
   XOR2_X1 U_dfifo_U_dcore_U_sub_fifo_U56 (.Z(U_dfifo_U_dcore_U_sub_fifo_n454), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n458), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n459));
   XNOR2_X1 U_dfifo_U_dcore_U_sub_fifo_U55 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n242), 
	.B(U_dfifo_U_dcore_U_sub_fifo_n566), 
	.A(FE_PHN1422_U_dfifo_U_dcore_U_sub_fifo_count_1_));
   INV_X4 U_dfifo_U_dcore_U_sub_fifo_U54 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n231), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n9));
   INV_X4 U_dfifo_U_dcore_U_sub_fifo_U53 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n232), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n10));
   OAI21_X1 U_dfifo_U_dcore_U_sub_fifo_U52 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n447), 
	.B2(FE_PHN3715_U_dfifo_U_dcore_U_sub_fifo_n127), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_n603), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n10));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U51 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n419), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4892_U_dfifo_U_dcore_U_sub_fifo_n202), 
	.A2(n84), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U50 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n422), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4791_U_dfifo_U_dcore_U_sub_fifo_n205), 
	.A2(n75), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U49 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n421), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4741_U_dfifo_U_dcore_U_sub_fifo_n204), 
	.A2(n74), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U48 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n420), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN3761_U_dfifo_U_dcore_U_sub_fifo_n203), 
	.A2(n85), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U47 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n424), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4852_U_dfifo_U_dcore_U_sub_fifo_n207), 
	.A2(n77), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U46 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n425), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4764_U_dfifo_U_dcore_U_sub_fifo_n208), 
	.A2(n78), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U45 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n426), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4816_U_dfifo_U_dcore_U_sub_fifo_n209), 
	.A2(n79), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U44 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n427), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4929_U_dfifo_U_dcore_U_sub_fifo_n210), 
	.A2(n80), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U43 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n423), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4757_U_dfifo_U_dcore_U_sub_fifo_n206), 
	.A2(n76), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U42 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n428), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4786_U_dfifo_U_dcore_U_sub_fifo_n211), 
	.A2(n81), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U41 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n429), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4836_U_dfifo_U_dcore_U_sub_fifo_n212), 
	.A2(n82), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U40 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n430), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4975_U_dfifo_U_dcore_U_sub_fifo_n213), 
	.A2(n83), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U39 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n431), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4837_U_dfifo_U_dcore_U_sub_fifo_n214), 
	.A2(n61), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U38 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n432), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4773_U_dfifo_U_dcore_U_sub_fifo_n215), 
	.A2(n62), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U37 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n433), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4908_U_dfifo_U_dcore_U_sub_fifo_n216), 
	.A2(n63), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U36 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n434), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN3792_U_dfifo_U_dcore_U_sub_fifo_n217), 
	.A2(n64), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U35 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n435), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4817_U_dfifo_U_dcore_U_sub_fifo_n218), 
	.A2(n65), 
	.A1(FE_OFN273_U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U34 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n436), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4771_U_dfifo_U_dcore_U_sub_fifo_n219), 
	.A2(n66), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U33 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n437), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
	.B1(FE_PHN4762_U_dfifo_U_dcore_U_sub_fifo_n220), 
	.A2(n67), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n234));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U32 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n379), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN3827_U_dfifo_U_dcore_U_sub_fifo_n162), 
	.A2(n69), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U31 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n380), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4872_U_dfifo_U_dcore_U_sub_fifo_n163), 
	.A2(n68), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U30 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n381), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4903_U_dfifo_U_dcore_U_sub_fifo_n164), 
	.A2(n70), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U29 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n382), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4811_U_dfifo_U_dcore_U_sub_fifo_n165), 
	.A2(n71), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U28 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n383), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4846_U_dfifo_U_dcore_U_sub_fifo_n166), 
	.A2(n72), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U27 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n384), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4753_U_dfifo_U_dcore_U_sub_fifo_n167), 
	.A2(n73), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U26 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n385), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4825_U_dfifo_U_dcore_U_sub_fifo_n168), 
	.A2(n84), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U25 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n386), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4826_U_dfifo_U_dcore_U_sub_fifo_n169), 
	.A2(n85), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U24 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n387), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4803_U_dfifo_U_dcore_U_sub_fifo_n170), 
	.A2(n74), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U23 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n388), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN3944_U_dfifo_U_dcore_U_sub_fifo_n171), 
	.A2(n75), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U22 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n389), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4875_U_dfifo_U_dcore_U_sub_fifo_n172), 
	.A2(n76), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U21 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n390), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4800_U_dfifo_U_dcore_U_sub_fifo_n173), 
	.A2(n77), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U20 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n391), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4880_U_dfifo_U_dcore_U_sub_fifo_n174), 
	.A2(n78), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U19 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n392), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4799_U_dfifo_U_dcore_U_sub_fifo_n175), 
	.A2(n79), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U18 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n393), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4879_U_dfifo_U_dcore_U_sub_fifo_n176), 
	.A2(n80), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U17 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n394), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN3838_U_dfifo_U_dcore_U_sub_fifo_n177), 
	.A2(n81), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U16 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n395), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN5041_U_dfifo_U_dcore_U_sub_fifo_n178), 
	.A2(n82), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U15 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n396), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
	.B1(FE_PHN4848_U_dfifo_U_dcore_U_sub_fifo_n179), 
	.A2(n83), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_n233));
   NOR3_X2 U_dfifo_U_dcore_U_sub_fifo_U14 (.ZN(U_dfifo_U_dcore_m_sf_empty), 
	.A3(FE_PHN1422_U_dfifo_U_dcore_U_sub_fifo_count_1_), 
	.A2(FE_PHN1595_U_dfifo_U_dcore_U_sub_fifo_count_0_), 
	.A1(U_dfifo_U_dcore_U_sub_fifo_count_2_));
   MUX2_X1 U_dfifo_U_dcore_U_sub_fifo_U13 (.Z(U_dfifo_U_dcore_U_sub_fifo_n459), 
	.S(FE_PHN1595_U_dfifo_U_dcore_U_sub_fifo_count_0_), 
	.B(U_dfifo_U_dcore_n209), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n609));
   AOI21_X1 U_dfifo_U_dcore_U_sub_fifo_U12 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n566), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n565), 
	.B1(U_dfifo_U_dcore_n208), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n456));
   INV_X4 U_dfifo_U_dcore_U_sub_fifo_U11 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n7), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n15));
   INV_X4 U_dfifo_U_dcore_U_sub_fifo_U10 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n6), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n16));
   OAI221_X1 U_dfifo_U_dcore_U_sub_fifo_U8 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n450), 
	.C2(U_dfifo_U_dcore_U_sub_fifo_n5), 
	.C1(U_dfifo_U_dcore_U_sub_fifo_n17), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n1), 
	.B1(U_dfifo_U_dcore_U_sub_fifo_count_2_), 
	.A(U_dfifo_U_dcore_n24));
   AOI21_X1 U_dfifo_U_dcore_U_sub_fifo_U7 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n5), 
	.B2(FE_PHN1595_U_dfifo_U_dcore_U_sub_fifo_count_0_), 
	.B1(U_dfifo_U_dcore_n208), 
	.A(U_dfifo_U_dcore_U_sub_fifo_n4));
   OAI22_X1 U_dfifo_U_dcore_U_sub_fifo_U6 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n4), 
	.B2(U_dfifo_U_dcore_U_sub_fifo_n608), 
	.B1(U_dfifo_U_dcore_n208), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n3), 
	.A1(FE_PHN1422_U_dfifo_U_dcore_U_sub_fifo_count_1_));
   INV_X1 U_dfifo_U_dcore_U_sub_fifo_U5 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n3), 
	.A(U_dfifo_U_dcore_n209));
   NAND2_X1 U_dfifo_U_dcore_U_sub_fifo_U3 (.ZN(U_dfifo_U_dcore_U_sub_fifo_n1), 
	.A2(U_dfifo_U_dcore_U_sub_fifo_n456), 
	.A1(FE_PHN1422_U_dfifo_U_dcore_U_sub_fifo_count_1_));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_out_ptr_reg_0_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n18), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_), 
	.D(U_dfifo_U_dcore_U_sub_fifo_n453), 
	.CK(HCLK__L5_N4));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_out_ptr_reg_1_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n56), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_out_ptr_1_), 
	.D(FE_PHN1842_U_dfifo_U_dcore_U_sub_fifo_n451), 
	.CK(HCLK__L5_N4));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_out_ptr_reg_2_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n126), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_), 
	.D(FE_PHN1184_U_dfifo_U_dcore_U_sub_fifo_n452), 
	.CK(HCLK__L5_N4));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__5_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n78), 
	.D(FE_PHN2202_U_dfifo_U_dcore_U_sub_fifo_n373), 
	.CK(HCLK__L5_N15));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__6_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n77), 
	.D(FE_PHN2110_U_dfifo_U_dcore_U_sub_fifo_n372), 
	.CK(HCLK__L5_N18));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__7_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n76), 
	.D(FE_PHN1942_U_dfifo_U_dcore_U_sub_fifo_n371), 
	.CK(HCLK__L5_N15));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__8_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n75), 
	.D(FE_PHN1924_U_dfifo_U_dcore_U_sub_fifo_n370), 
	.CK(HCLK__L5_N15));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__9_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n74), 
	.D(FE_PHN2115_U_dfifo_U_dcore_U_sub_fifo_n369), 
	.CK(HCLK__L5_N15));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__10_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n73), 
	.D(FE_PHN2209_U_dfifo_U_dcore_U_sub_fifo_n368), 
	.CK(HCLK__L5_N16));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__11_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n72), 
	.D(FE_PHN1958_U_dfifo_U_dcore_U_sub_fifo_n367), 
	.CK(HCLK__L5_N18));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__12_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n71), 
	.D(FE_PHN2184_U_dfifo_U_dcore_U_sub_fifo_n366), 
	.CK(HCLK__L5_N18));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__13_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n70), 
	.D(FE_PHN2182_U_dfifo_U_dcore_U_sub_fifo_n365), 
	.CK(HCLK__L5_N18));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__14_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n69), 
	.D(FE_PHN1968_U_dfifo_U_dcore_U_sub_fifo_n364), 
	.CK(HCLK__L5_N16));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__15_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n68), 
	.D(FE_PHN2159_U_dfifo_U_dcore_U_sub_fifo_n363), 
	.CK(HCLK__L5_N18));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__16_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n67), 
	.D(FE_PHN1946_U_dfifo_U_dcore_U_sub_fifo_n362), 
	.CK(HCLK__L5_N18));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__17_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n66), 
	.D(FE_PHN2151_U_dfifo_U_dcore_U_sub_fifo_n361), 
	.CK(HCLK__L5_N16));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__18_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n125), 
	.D(FE_PHN1963_U_dfifo_U_dcore_U_sub_fifo_n360), 
	.CK(HCLK__L5_N16));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__19_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n124), 
	.D(FE_PHN1928_U_dfifo_U_dcore_U_sub_fifo_n359), 
	.CK(HCLK__L5_N15));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__20_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n123), 
	.D(FE_PHN1955_U_dfifo_U_dcore_U_sub_fifo_n358), 
	.CK(HCLK__L5_N15));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__21_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n122), 
	.D(FE_PHN1943_U_dfifo_U_dcore_U_sub_fifo_n357), 
	.CK(HCLK__L5_N6));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__22_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n121), 
	.D(FE_PHN1927_U_dfifo_U_dcore_U_sub_fifo_n356), 
	.CK(HCLK__L5_N14));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__23_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n120), 
	.D(FE_PHN1945_U_dfifo_U_dcore_U_sub_fifo_n355), 
	.CK(HCLK__L5_N16));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__24_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n119), 
	.D(FE_PHN1922_U_dfifo_U_dcore_U_sub_fifo_n354), 
	.CK(HCLK__L5_N16));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__25_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n118), 
	.D(FE_PHN1941_U_dfifo_U_dcore_U_sub_fifo_n353), 
	.CK(HCLK__L5_N14));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__26_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n65), 
	.D(FE_PHN1965_U_dfifo_U_dcore_U_sub_fifo_n352), 
	.CK(HCLK__L5_N14));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__27_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n64), 
	.D(FE_PHN1960_U_dfifo_U_dcore_U_sub_fifo_n351), 
	.CK(HCLK__L5_N18));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__28_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n63), 
	.D(FE_PHN2221_U_dfifo_U_dcore_U_sub_fifo_n350), 
	.CK(HCLK__L5_N14));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__29_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n62), 
	.D(FE_PHN1969_U_dfifo_U_dcore_U_sub_fifo_n349), 
	.CK(HCLK__L5_N14));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__30_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n61), 
	.D(FE_PHN1952_U_dfifo_U_dcore_U_sub_fifo_n348), 
	.CK(HCLK__L5_N14));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__31_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n60), 
	.D(FE_PHN1957_U_dfifo_U_dcore_U_sub_fifo_n347), 
	.CK(HCLK__L5_N14));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__32_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n59), 
	.D(FE_PHN1961_U_dfifo_U_dcore_U_sub_fifo_n346), 
	.CK(HCLK__L5_N14));
   DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__33_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n58), 
	.D(FE_PHN1949_U_dfifo_U_dcore_U_sub_fifo_n345), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_count_reg_1_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n54), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_count_1_), 
	.D(FE_PHN1591_U_dfifo_U_dcore_U_sub_fifo_n242), 
	.CK(HCLK__L5_N5));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__33_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n19), 
	.D(FE_PHN2320_U_dfifo_U_dcore_U_sub_fifo_n243), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__32_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n20), 
	.D(FE_PHN2305_U_dfifo_U_dcore_U_sub_fifo_n244), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__31_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n21), 
	.D(FE_PHN2309_U_dfifo_U_dcore_U_sub_fifo_n245), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__30_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n22), 
	.D(FE_PHN2334_U_dfifo_U_dcore_U_sub_fifo_n246), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__29_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n23), 
	.D(FE_PHN2296_U_dfifo_U_dcore_U_sub_fifo_n247), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__28_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n24), 
	.D(FE_PHN2331_U_dfifo_U_dcore_U_sub_fifo_n248), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__27_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n25), 
	.D(FE_PHN2332_U_dfifo_U_dcore_U_sub_fifo_n249), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__26_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n26), 
	.D(FE_PHN2323_U_dfifo_U_dcore_U_sub_fifo_n250), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__25_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n27), 
	.D(FE_PHN2288_U_dfifo_U_dcore_U_sub_fifo_n251), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__24_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n28), 
	.D(FE_PHN2293_U_dfifo_U_dcore_U_sub_fifo_n252), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__23_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n29), 
	.D(FE_PHN2352_U_dfifo_U_dcore_U_sub_fifo_n253), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__22_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n30), 
	.D(FE_PHN2341_U_dfifo_U_dcore_U_sub_fifo_n254), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__21_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n31), 
	.D(FE_PHN2342_U_dfifo_U_dcore_U_sub_fifo_n255), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__20_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n32), 
	.D(FE_PHN2326_U_dfifo_U_dcore_U_sub_fifo_n256), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__19_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n33), 
	.D(FE_PHN2353_U_dfifo_U_dcore_U_sub_fifo_n257), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__18_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n34), 
	.D(FE_PHN2344_U_dfifo_U_dcore_U_sub_fifo_n258), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__17_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n35), 
	.D(FE_PHN2318_U_dfifo_U_dcore_U_sub_fifo_n259), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__16_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n36), 
	.D(FE_PHN2369_U_dfifo_U_dcore_U_sub_fifo_n260), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__15_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n37), 
	.D(FE_PHN2319_U_dfifo_U_dcore_U_sub_fifo_n261), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__14_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n38), 
	.D(FE_PHN2335_U_dfifo_U_dcore_U_sub_fifo_n262), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__13_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n39), 
	.D(FE_PHN2325_U_dfifo_U_dcore_U_sub_fifo_n263), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__12_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n40), 
	.D(FE_PHN2023_U_dfifo_U_dcore_U_sub_fifo_n264), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__11_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n41), 
	.D(FE_PHN2349_U_dfifo_U_dcore_U_sub_fifo_n265), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__10_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n42), 
	.D(FE_PHN2310_U_dfifo_U_dcore_U_sub_fifo_n266), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__9_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n43), 
	.D(FE_PHN2339_U_dfifo_U_dcore_U_sub_fifo_n267), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__8_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n44), 
	.D(FE_PHN2357_U_dfifo_U_dcore_U_sub_fifo_n268), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__7_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n45), 
	.D(FE_PHN2361_U_dfifo_U_dcore_U_sub_fifo_n269), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__6_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n46), 
	.D(FE_PHN2360_U_dfifo_U_dcore_U_sub_fifo_n270), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__5_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n47), 
	.D(FE_PHN2374_U_dfifo_U_dcore_U_sub_fifo_n271), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__4_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n48), 
	.D(FE_PHN2375_U_dfifo_U_dcore_U_sub_fifo_n272), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__3_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n49), 
	.D(FE_PHN2304_U_dfifo_U_dcore_U_sub_fifo_n273), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__2_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n50), 
	.D(FE_PHN2340_U_dfifo_U_dcore_U_sub_fifo_n274), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__1_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n51), 
	.D(FE_PHN2363_U_dfifo_U_dcore_U_sub_fifo_n275), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__0_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n52), 
	.D(FE_PHN2336_U_dfifo_U_dcore_U_sub_fifo_n276), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__33_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n84), 
	.D(FE_PHN2338_U_dfifo_U_dcore_U_sub_fifo_n277), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__32_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n85), 
	.D(FE_PHN2366_U_dfifo_U_dcore_U_sub_fifo_n278), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__31_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n86), 
	.D(FE_PHN2350_U_dfifo_U_dcore_U_sub_fifo_n279), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__30_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n87), 
	.D(FE_PHN2291_U_dfifo_U_dcore_U_sub_fifo_n280), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__29_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n88), 
	.D(FE_PHN2285_U_dfifo_U_dcore_U_sub_fifo_n281), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__28_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n89), 
	.D(FE_PHN2329_U_dfifo_U_dcore_U_sub_fifo_n282), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__27_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n90), 
	.D(FE_PHN2358_U_dfifo_U_dcore_U_sub_fifo_n283), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__26_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n91), 
	.D(FE_PHN2317_U_dfifo_U_dcore_U_sub_fifo_n284), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__25_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n92), 
	.D(FE_PHN2280_U_dfifo_U_dcore_U_sub_fifo_n285), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__24_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n93), 
	.D(FE_PHN2337_U_dfifo_U_dcore_U_sub_fifo_n286), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__23_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n94), 
	.D(FE_PHN2313_U_dfifo_U_dcore_U_sub_fifo_n287), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__22_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n95), 
	.D(FE_PHN2289_U_dfifo_U_dcore_U_sub_fifo_n288), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__21_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n96), 
	.D(FE_PHN2314_U_dfifo_U_dcore_U_sub_fifo_n289), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__20_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n97), 
	.D(FE_PHN2345_U_dfifo_U_dcore_U_sub_fifo_n290), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__19_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n98), 
	.D(FE_PHN2284_U_dfifo_U_dcore_U_sub_fifo_n291), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__18_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n99), 
	.D(FE_PHN2354_U_dfifo_U_dcore_U_sub_fifo_n292), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__17_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n100), 
	.D(FE_PHN2298_U_dfifo_U_dcore_U_sub_fifo_n293), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__16_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n101), 
	.D(FE_PHN2370_U_dfifo_U_dcore_U_sub_fifo_n294), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__15_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n102), 
	.D(FE_PHN2368_U_dfifo_U_dcore_U_sub_fifo_n295), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__14_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n103), 
	.D(FE_PHN2301_U_dfifo_U_dcore_U_sub_fifo_n296), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__13_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n104), 
	.D(FE_PHN2283_U_dfifo_U_dcore_U_sub_fifo_n297), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__12_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n105), 
	.D(FE_PHN2311_U_dfifo_U_dcore_U_sub_fifo_n298), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__11_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n106), 
	.D(FE_PHN2327_U_dfifo_U_dcore_U_sub_fifo_n299), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__10_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n107), 
	.D(FE_PHN2306_U_dfifo_U_dcore_U_sub_fifo_n300), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__9_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n108), 
	.D(FE_PHN2303_U_dfifo_U_dcore_U_sub_fifo_n301), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__8_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n109), 
	.D(FE_PHN2322_U_dfifo_U_dcore_U_sub_fifo_n302), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__7_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n110), 
	.D(FE_PHN2372_U_dfifo_U_dcore_U_sub_fifo_n303), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__6_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n111), 
	.D(FE_PHN2299_U_dfifo_U_dcore_U_sub_fifo_n304), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__5_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n112), 
	.D(FE_PHN2365_U_dfifo_U_dcore_U_sub_fifo_n305), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__4_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n113), 
	.D(FE_PHN2371_U_dfifo_U_dcore_U_sub_fifo_n306), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__3_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n114), 
	.D(FE_PHN2356_U_dfifo_U_dcore_U_sub_fifo_n307), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__2_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n115), 
	.D(FE_PHN2297_U_dfifo_U_dcore_U_sub_fifo_n308), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__1_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n116), 
	.D(FE_PHN2367_U_dfifo_U_dcore_U_sub_fifo_n309), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__0_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n117), 
	.D(FE_PHN2307_U_dfifo_U_dcore_U_sub_fifo_n310), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__33_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n128), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__33_), 
	.D(FE_PHN2113_U_dfifo_U_dcore_U_sub_fifo_n311), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__32_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n129), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__32_), 
	.D(FE_PHN2124_U_dfifo_U_dcore_U_sub_fifo_n312), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__31_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n130), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__31_), 
	.D(FE_PHN2160_U_dfifo_U_dcore_U_sub_fifo_n313), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__30_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n131), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__30_), 
	.D(FE_PHN2205_U_dfifo_U_dcore_U_sub_fifo_n314), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__29_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n132), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__29_), 
	.D(FE_PHN2142_U_dfifo_U_dcore_U_sub_fifo_n315), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__28_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n133), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__28_), 
	.D(FE_PHN2108_U_dfifo_U_dcore_U_sub_fifo_n316), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__27_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n134), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__27_), 
	.D(FE_PHN2175_U_dfifo_U_dcore_U_sub_fifo_n317), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__26_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n135), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__26_), 
	.D(FE_PHN1951_U_dfifo_U_dcore_U_sub_fifo_n318), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__25_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n136), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__25_), 
	.D(FE_PHN2126_U_dfifo_U_dcore_U_sub_fifo_n319), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__24_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n137), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__24_), 
	.D(FE_PHN2128_U_dfifo_U_dcore_U_sub_fifo_n320), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__23_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n138), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__23_), 
	.D(FE_PHN2167_U_dfifo_U_dcore_U_sub_fifo_n321), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__22_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n139), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__22_), 
	.D(FE_PHN2137_U_dfifo_U_dcore_U_sub_fifo_n322), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__21_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n140), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__21_), 
	.D(FE_PHN2123_U_dfifo_U_dcore_U_sub_fifo_n323), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__20_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n141), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__20_), 
	.D(FE_PHN1936_U_dfifo_U_dcore_U_sub_fifo_n324), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__19_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n142), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__19_), 
	.D(FE_PHN2134_U_dfifo_U_dcore_U_sub_fifo_n325), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__18_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n143), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__18_), 
	.D(FE_PHN2144_U_dfifo_U_dcore_U_sub_fifo_n326), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__17_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n144), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__17_), 
	.D(FE_PHN1939_U_dfifo_U_dcore_U_sub_fifo_n327), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__16_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n145), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__16_), 
	.D(FE_PHN2131_U_dfifo_U_dcore_U_sub_fifo_n328), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__15_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n146), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__15_), 
	.D(FE_PHN1780_U_dfifo_U_dcore_U_sub_fifo_n329), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__14_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n147), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__14_), 
	.D(FE_PHN1964_U_dfifo_U_dcore_U_sub_fifo_n330), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__13_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n148), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__13_), 
	.D(FE_PHN1925_U_dfifo_U_dcore_U_sub_fifo_n331), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__12_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n149), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__12_), 
	.D(FE_PHN1758_U_dfifo_U_dcore_U_sub_fifo_n332), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__11_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n150), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__11_), 
	.D(FE_PHN2152_U_dfifo_U_dcore_U_sub_fifo_n333), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__10_ (.RN(FE_OFN176_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n151), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__10_), 
	.D(FE_PHN1932_U_dfifo_U_dcore_U_sub_fifo_n334), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__9_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n152), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__9_), 
	.D(FE_PHN1923_U_dfifo_U_dcore_U_sub_fifo_n335), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__8_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n153), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__8_), 
	.D(FE_PHN1752_U_dfifo_U_dcore_U_sub_fifo_n336), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__7_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n154), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__7_), 
	.D(FE_PHN2216_U_dfifo_U_dcore_U_sub_fifo_n337), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__6_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n155), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__6_), 
	.D(FE_PHN1770_U_dfifo_U_dcore_U_sub_fifo_n338), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__5_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n156), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__5_), 
	.D(FE_PHN1756_U_dfifo_U_dcore_U_sub_fifo_n339), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__4_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n157), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__4_), 
	.D(FE_PHN1937_U_dfifo_U_dcore_U_sub_fifo_n340), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__3_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n158), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__3_), 
	.D(FE_PHN1940_U_dfifo_U_dcore_U_sub_fifo_n341), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__2_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n159), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__2_), 
	.D(FE_PHN2129_U_dfifo_U_dcore_U_sub_fifo_n342), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__1_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n160), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__1_), 
	.D(FE_PHN1933_U_dfifo_U_dcore_U_sub_fifo_n343), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__0_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n161), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_0__0_), 
	.D(FE_PHN1761_U_dfifo_U_dcore_U_sub_fifo_n344), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__4_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n79), 
	.D(FE_PHN2229_U_dfifo_U_dcore_U_sub_fifo_n374), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__3_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n80), 
	.D(FE_PHN1997_U_dfifo_U_dcore_U_sub_fifo_n375), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__2_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n81), 
	.D(FE_PHN2222_U_dfifo_U_dcore_U_sub_fifo_n376), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__1_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n82), 
	.D(FE_PHN1990_U_dfifo_U_dcore_U_sub_fifo_n377), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__0_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n83), 
	.D(FE_PHN2004_U_dfifo_U_dcore_U_sub_fifo_n378), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__33_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n162), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__33_), 
	.D(FE_PHN2190_U_dfifo_U_dcore_U_sub_fifo_n379), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__32_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n163), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__32_), 
	.D(FE_PHN2185_U_dfifo_U_dcore_U_sub_fifo_n380), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__31_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n164), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__31_), 
	.D(FE_PHN2217_U_dfifo_U_dcore_U_sub_fifo_n381), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__30_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n165), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__30_), 
	.D(FE_PHN2178_U_dfifo_U_dcore_U_sub_fifo_n382), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__29_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n166), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__29_), 
	.D(FE_PHN2170_U_dfifo_U_dcore_U_sub_fifo_n383), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__28_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n167), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__28_), 
	.D(FE_PHN2192_U_dfifo_U_dcore_U_sub_fifo_n384), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__27_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n168), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__27_), 
	.D(FE_PHN2188_U_dfifo_U_dcore_U_sub_fifo_n385), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__26_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n169), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__26_), 
	.D(FE_PHN2211_U_dfifo_U_dcore_U_sub_fifo_n386), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__25_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n170), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__25_), 
	.D(FE_PHN2207_U_dfifo_U_dcore_U_sub_fifo_n387), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__24_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n171), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__24_), 
	.D(FE_PHN2214_U_dfifo_U_dcore_U_sub_fifo_n388), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__23_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n172), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__23_), 
	.D(FE_PHN2176_U_dfifo_U_dcore_U_sub_fifo_n389), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__22_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n173), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__22_), 
	.D(FE_PHN2174_U_dfifo_U_dcore_U_sub_fifo_n390), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__21_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n174), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__21_), 
	.D(FE_PHN2173_U_dfifo_U_dcore_U_sub_fifo_n391), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__20_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n175), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__20_), 
	.D(FE_PHN2169_U_dfifo_U_dcore_U_sub_fifo_n392), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__19_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n176), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__19_), 
	.D(FE_PHN2168_U_dfifo_U_dcore_U_sub_fifo_n393), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__18_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n177), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__18_), 
	.D(FE_PHN2204_U_dfifo_U_dcore_U_sub_fifo_n394), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__17_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n178), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__17_), 
	.D(FE_PHN2162_U_dfifo_U_dcore_U_sub_fifo_n395), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__16_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n179), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__16_), 
	.D(FE_PHN2235_U_dfifo_U_dcore_U_sub_fifo_n396), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__15_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n180), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__15_), 
	.D(FE_PHN1947_U_dfifo_U_dcore_U_sub_fifo_n397), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__14_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n181), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__14_), 
	.D(FE_PHN1954_U_dfifo_U_dcore_U_sub_fifo_n398), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__13_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n182), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__13_), 
	.D(FE_PHN1944_U_dfifo_U_dcore_U_sub_fifo_n399), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__12_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n183), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__12_), 
	.D(FE_PHN2132_U_dfifo_U_dcore_U_sub_fifo_n400), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__11_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n184), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__11_), 
	.D(FE_PHN2158_U_dfifo_U_dcore_U_sub_fifo_n401), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__10_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n185), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__10_), 
	.D(FE_PHN2135_U_dfifo_U_dcore_U_sub_fifo_n402), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__9_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n186), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__9_), 
	.D(FE_PHN2138_U_dfifo_U_dcore_U_sub_fifo_n403), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__8_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n187), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__8_), 
	.D(FE_PHN2112_U_dfifo_U_dcore_U_sub_fifo_n404), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__7_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n188), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__7_), 
	.D(FE_PHN2139_U_dfifo_U_dcore_U_sub_fifo_n405), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__6_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n189), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__6_), 
	.D(FE_PHN2122_U_dfifo_U_dcore_U_sub_fifo_n406), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__5_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n190), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__5_), 
	.D(FE_PHN1956_U_dfifo_U_dcore_U_sub_fifo_n407), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__4_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n191), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__4_), 
	.D(FE_PHN2116_U_dfifo_U_dcore_U_sub_fifo_n408), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__3_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n192), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__3_), 
	.D(FE_PHN2117_U_dfifo_U_dcore_U_sub_fifo_n409), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__2_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n193), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__2_), 
	.D(FE_PHN1926_U_dfifo_U_dcore_U_sub_fifo_n410), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__1_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n194), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__1_), 
	.D(FE_PHN2136_U_dfifo_U_dcore_U_sub_fifo_n411), 
	.CK(HCLK__L5_N5));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__0_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n195), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_2__0_), 
	.D(FE_PHN2121_U_dfifo_U_dcore_U_sub_fifo_n412), 
	.CK(HCLK__L5_N6));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__33_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n196), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__33_), 
	.D(FE_PHN2165_U_dfifo_U_dcore_U_sub_fifo_n413), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__32_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n197), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__32_), 
	.D(FE_PHN2127_U_dfifo_U_dcore_U_sub_fifo_n414), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__31_ (.RN(FE_OFN143_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n198), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__31_), 
	.D(FE_PHN1953_U_dfifo_U_dcore_U_sub_fifo_n415), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__30_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n199), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__30_), 
	.D(FE_PHN2153_U_dfifo_U_dcore_U_sub_fifo_n416), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__29_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n200), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__29_), 
	.D(FE_PHN1938_U_dfifo_U_dcore_U_sub_fifo_n417), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__28_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n201), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__28_), 
	.D(FE_PHN1930_U_dfifo_U_dcore_U_sub_fifo_n418), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__27_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n202), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__27_), 
	.D(FE_PHN2171_U_dfifo_U_dcore_U_sub_fifo_n419), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__26_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n203), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__26_), 
	.D(FE_PHN2155_U_dfifo_U_dcore_U_sub_fifo_n420), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__25_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n204), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__25_), 
	.D(FE_PHN2193_U_dfifo_U_dcore_U_sub_fifo_n421), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__24_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n205), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__24_), 
	.D(FE_PHN2218_U_dfifo_U_dcore_U_sub_fifo_n422), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__23_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n206), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__23_), 
	.D(FE_PHN2199_U_dfifo_U_dcore_U_sub_fifo_n423), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__22_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n207), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__22_), 
	.D(FE_PHN2177_U_dfifo_U_dcore_U_sub_fifo_n424), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__21_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n208), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__21_), 
	.D(FE_PHN2172_U_dfifo_U_dcore_U_sub_fifo_n425), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__20_ (.RN(FE_OFN136_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n209), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__20_), 
	.D(FE_PHN2197_U_dfifo_U_dcore_U_sub_fifo_n426), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__19_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n210), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__19_), 
	.D(FE_PHN2213_U_dfifo_U_dcore_U_sub_fifo_n427), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__18_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n211), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__18_), 
	.D(FE_PHN2195_U_dfifo_U_dcore_U_sub_fifo_n428), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__17_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n212), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__17_), 
	.D(FE_PHN2183_U_dfifo_U_dcore_U_sub_fifo_n429), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__16_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n213), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__16_), 
	.D(FE_PHN2220_U_dfifo_U_dcore_U_sub_fifo_n430), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__15_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n214), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__15_), 
	.D(FE_PHN2186_U_dfifo_U_dcore_U_sub_fifo_n431), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__14_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n215), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__14_), 
	.D(FE_PHN2206_U_dfifo_U_dcore_U_sub_fifo_n432), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__13_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n216), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__13_), 
	.D(FE_PHN2198_U_dfifo_U_dcore_U_sub_fifo_n433), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__12_ (.RN(FE_OFN69_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n217), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__12_), 
	.D(FE_PHN2201_U_dfifo_U_dcore_U_sub_fifo_n434), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__11_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n218), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__11_), 
	.D(FE_PHN2203_U_dfifo_U_dcore_U_sub_fifo_n435), 
	.CK(HCLK__L5_N18));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__10_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n219), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__10_), 
	.D(FE_PHN2191_U_dfifo_U_dcore_U_sub_fifo_n436), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__9_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n220), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__9_), 
	.D(FE_PHN2194_U_dfifo_U_dcore_U_sub_fifo_n437), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__8_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n221), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__8_), 
	.D(FE_PHN2130_U_dfifo_U_dcore_U_sub_fifo_n438), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__7_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n222), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__7_), 
	.D(FE_PHN2111_U_dfifo_U_dcore_U_sub_fifo_n439), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__6_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n223), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__6_), 
	.D(FE_PHN1935_U_dfifo_U_dcore_U_sub_fifo_n440), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__5_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n224), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__5_), 
	.D(FE_PHN2118_U_dfifo_U_dcore_U_sub_fifo_n441), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__4_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n225), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__4_), 
	.D(FE_PHN1931_U_dfifo_U_dcore_U_sub_fifo_n442), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__3_ (.RN(FE_OFN157_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n226), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__3_), 
	.D(FE_PHN2147_U_dfifo_U_dcore_U_sub_fifo_n443), 
	.CK(HCLK__L5_N15));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__2_ (.RN(FE_OFN67_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n227), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__2_), 
	.D(FE_PHN2119_U_dfifo_U_dcore_U_sub_fifo_n444), 
	.CK(HCLK__L5_N16));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__1_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n228), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__1_), 
	.D(FE_PHN2208_U_dfifo_U_dcore_U_sub_fifo_n445), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__0_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n229), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_mem_3__0_), 
	.D(FE_PHN1929_U_dfifo_U_dcore_U_sub_fifo_n446), 
	.CK(HCLK__L5_N14));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_in_ptr_reg_1_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n127), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_), 
	.D(FE_PHN1460_U_dfifo_U_dcore_U_sub_fifo_n447), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_in_ptr_reg_2_ (.RN(FE_OFN62_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n57), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_in_ptr_2_), 
	.D(FE_PHN4294_U_dfifo_U_dcore_U_sub_fifo_n448), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_in_ptr_reg_0_ (.RN(FE_OFN42_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n55), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_in_ptr_0_), 
	.D(U_dfifo_U_dcore_U_sub_fifo_n449), 
	.CK(HCLK__L5_N4));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_count_reg_2_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n17), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_count_2_), 
	.D(FE_PHN789_U_dfifo_U_dcore_U_sub_fifo_n450), 
	.CK(HCLK__L5_N5));
   DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_count_reg_0_ (.RN(FE_OFN43_HRESETn), 
	.QN(U_dfifo_U_dcore_U_sub_fifo_n13), 
	.Q(U_dfifo_U_dcore_U_sub_fifo_count_0_), 
	.D(U_dfifo_U_dcore_U_sub_fifo_n454), 
	.CK(HCLK__L5_N5));
   NOR2_X1 U3 (.ZN(n10), 
	.A2(U_ctl_n288), 
	.A1(FE_PHN1079_U_ctl_n400));
   AOI22_X1 U4 (.ZN(n11), 
	.B2(n10), 
	.B1(U_afifo_n140), 
	.A2(U_afifo_f_data2_12_), 
	.A1(U_afifo_n54));
   INV_X1 U5 (.ZN(U_afifo_m_data_in[12]), 
	.A(n11));
   AOI22_X1 U6 (.ZN(n12), 
	.B2(U_afifo_n54), 
	.B1(U_afifo_f_data2_16_), 
	.A2(U_afifo_n98), 
	.A1(haddr[6]));
   INV_X1 U7 (.ZN(U_afifo_m_data_in[16]), 
	.A(n12));
   AOI22_X1 U8 (.ZN(n13), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1817_U_afifo_f_data2_41_), 
	.A2(U_afifo_n99), 
	.A1(haddr[31]));
   INV_X1 U9 (.ZN(U_afifo_m_data_in[41]), 
	.A(FE_PHN1432_n13));
   AOI22_X1 U10 (.ZN(n14), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1859_U_afifo_f_data2_36_), 
	.A2(FE_OFN236_U_afifo_n93), 
	.A1(haddr[26]));
   INV_X1 U11 (.ZN(U_afifo_m_data_in[36]), 
	.A(n14));
   AOI22_X1 U12 (.ZN(n15), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1858_U_afifo_f_data2_28_), 
	.A2(U_afifo_n147), 
	.A1(haddr[18]));
   INV_X1 U13 (.ZN(U_afifo_m_data_in[28]), 
	.A(n15));
   AOI22_X1 U14 (.ZN(n16), 
	.B2(U_afifo_n54), 
	.B1(U_afifo_f_data2_17_), 
	.A2(U_afifo_n98), 
	.A1(haddr[7]));
   INV_X1 U15 (.ZN(U_afifo_m_data_in[17]), 
	.A(n16));
   AOI22_X1 U16 (.ZN(n17), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1869_U_afifo_f_data2_40_), 
	.A2(U_afifo_n140), 
	.A1(haddr[30]));
   INV_X1 U17 (.ZN(U_afifo_m_data_in[40]), 
	.A(FE_PHN1525_n17));
   AOI22_X1 U18 (.ZN(n18), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1870_U_afifo_f_data2_35_), 
	.A2(FE_OFN236_U_afifo_n93), 
	.A1(haddr[25]));
   INV_X1 U19 (.ZN(U_afifo_m_data_in[35]), 
	.A(n18));
   AOI22_X1 U20 (.ZN(n19), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1883_U_afifo_f_data2_31_), 
	.A2(U_afifo_n99), 
	.A1(haddr[21]));
   INV_X1 U21 (.ZN(U_afifo_m_data_in[31]), 
	.A(n19));
   AOI22_X1 U22 (.ZN(n20), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1867_U_afifo_f_data2_27_), 
	.A2(U_afifo_n147), 
	.A1(haddr[17]));
   INV_X1 U23 (.ZN(U_afifo_m_data_in[27]), 
	.A(n20));
   INV_X1 U24 (.ZN(n21), 
	.A(U_ctl_n308));
   NOR3_X1 U25 (.ZN(n22), 
	.A3(n21), 
	.A2(U_ctl_n97), 
	.A1(U_ctl_fr_prv_1wrap));
   NOR4_X1 U26 (.ZN(n23), 
	.A4(m_df_push_n), 
	.A3(n22), 
	.A2(hiu_rw), 
	.A1(miu_pop_n));
   OAI221_X1 U27 (.ZN(U_ctl_n304), 
	.C2(U_dfifo_m_aempty), 
	.C1(U_dfifo_m_empty), 
	.B2(U_dfifo_n5), 
	.B1(U_dfifo_m_empty), 
	.A(n23));
   AOI22_X1 U28 (.ZN(n24), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1871_U_afifo_f_data2_39_), 
	.A2(U_afifo_n98), 
	.A1(haddr[29]));
   INV_X1 U29 (.ZN(U_afifo_m_data_in[39]), 
	.A(n24));
   AOI22_X1 U30 (.ZN(n25), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1857_U_afifo_f_data2_34_), 
	.A2(FE_OFN236_U_afifo_n93), 
	.A1(haddr[24]));
   INV_X1 U31 (.ZN(U_afifo_m_data_in[34]), 
	.A(FE_PHN1777_n25));
   AOI22_X1 U32 (.ZN(n26), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1856_U_afifo_f_data2_33_), 
	.A2(U_afifo_n140), 
	.A1(haddr[23]));
   INV_X1 U33 (.ZN(U_afifo_m_data_in[33]), 
	.A(n26));
   AOI22_X1 U34 (.ZN(n27), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1873_U_afifo_f_data2_26_), 
	.A2(U_afifo_n147), 
	.A1(haddr[16]));
   INV_X1 U35 (.ZN(U_afifo_m_data_in[26]), 
	.A(FE_PHN1798_n27));
   AOI22_X1 U36 (.ZN(n28), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1876_U_afifo_f_data2_24_), 
	.A2(U_afifo_n99), 
	.A1(haddr[14]));
   INV_X1 U37 (.ZN(U_afifo_m_data_in[24]), 
	.A(n28));
   OAI22_X2 U38 (.ZN(hiu_burst_size[5]), 
	.B2(U_afifo_U_acore_n32), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n8), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   AOI22_X1 U39 (.ZN(n29), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1878_U_afifo_f_data2_37_), 
	.A2(U_afifo_n98), 
	.A1(haddr[27]));
   INV_X1 U40 (.ZN(U_afifo_m_data_in[37]), 
	.A(FE_PHN1689_n29));
   AOI22_X1 U41 (.ZN(n30), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1861_U_afifo_f_data2_30_), 
	.A2(U_afifo_n140), 
	.A1(haddr[20]));
   INV_X1 U42 (.ZN(U_afifo_m_data_in[30]), 
	.A(n30));
   AOI22_X1 U43 (.ZN(n31), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1866_U_afifo_f_data2_29_), 
	.A2(FE_OFN236_U_afifo_n93), 
	.A1(haddr[19]));
   INV_X1 U44 (.ZN(U_afifo_m_data_in[29]), 
	.A(n31));
   AOI22_X1 U45 (.ZN(n32), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1880_U_afifo_f_data2_20_), 
	.A2(U_afifo_n147), 
	.A1(haddr[10]));
   INV_X1 U46 (.ZN(U_afifo_m_data_in[20]), 
	.A(n32));
   AOI22_X1 U47 (.ZN(n33), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1862_U_afifo_f_data2_2_), 
	.A2(U_afifo_n99), 
	.A1(m_af_data1_in_2_));
   INV_X1 U48 (.ZN(U_afifo_m_data_in[2]), 
	.A(n33));
   INV_X1 U49 (.ZN(n34), 
	.A(U_rbuf_n123));
   AOI21_X1 U50 (.ZN(U_rbuf_n161), 
	.B2(n34), 
	.B1(U_rbuf_n34), 
	.A(miu_push_n));
   OAI22_X2 U51 (.ZN(hiu_burst_size[0]), 
	.B2(FE_PHN1847_U_afifo_U_acore_n181), 
	.B1(FE_OFN26_U_afifo_U_acore_n38), 
	.A2(U_afifo_U_acore_n4), 
	.A1(FE_OFN250_U_afifo_U_acore_n1));
   AOI22_X1 U55 (.ZN(n37), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1865_U_afifo_f_data2_25_), 
	.A2(U_afifo_n98), 
	.A1(haddr[15]));
   INV_X1 U56 (.ZN(U_afifo_m_data_in[25]), 
	.A(FE_PHN1838_n37));
   AOI22_X1 U57 (.ZN(n38), 
	.B2(U_afifo_n54), 
	.B1(FE_PHN1874_U_afifo_f_data2_23_), 
	.A2(U_afifo_n99), 
	.A1(haddr[13]));
   INV_X1 U58 (.ZN(U_afifo_m_data_in[23]), 
	.A(n38));
   AOI22_X1 U59 (.ZN(n39), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1864_U_afifo_f_data2_22_), 
	.A2(FE_OFN236_U_afifo_n93), 
	.A1(haddr[12]));
   INV_X1 U60 (.ZN(U_afifo_m_data_in[22]), 
	.A(FE_PHN1762_n39));
   AOI22_X1 U61 (.ZN(n40), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1853_U_afifo_f_data2_21_), 
	.A2(U_afifo_n140), 
	.A1(haddr[11]));
   INV_X1 U62 (.ZN(U_afifo_m_data_in[21]), 
	.A(n40));
   AOI22_X1 U63 (.ZN(n41), 
	.B2(FE_OFN237_U_afifo_n54), 
	.B1(FE_PHN1860_U_afifo_f_data2_19_), 
	.A2(U_afifo_n147), 
	.A1(haddr[9]));
   INV_X1 U64 (.ZN(U_afifo_m_data_in[19]), 
	.A(n41));
   AOI211_X1 U67 (.ZN(U_ctl_n118), 
	.C2(U_ctl_n145), 
	.C1(U_ctl_n395), 
	.B(U_ctl_n323), 
	.A(1'b0));
   OAI22_X1 U70 (.ZN(U_afifo_n21), 
	.B2(1'b0), 
	.B1(FE_PHN2433_U_afifo_n164), 
	.A2(1'b1), 
	.A1(1'b0));
   OAI21_X1 U72 (.ZN(U_afifo_n12), 
	.B2(1'b0), 
	.B1(FE_PHN2434_U_afifo_n158), 
	.A(1'b1));
   INV_X2 U73 (.ZN(U_afifo_m_data_in[48]), 
	.A(U_afifo_n15));
   INV_X2 U76 (.ZN(U_rbuf_n181), 
	.A(miu_data[0]));
   INV_X2 U77 (.ZN(U_rbuf_n182), 
	.A(miu_data[1]));
   INV_X2 U78 (.ZN(U_rbuf_n184), 
	.A(miu_data[3]));
   INV_X2 U79 (.ZN(U_rbuf_n186), 
	.A(miu_data[5]));
   INV_X2 U80 (.ZN(U_rbuf_n187), 
	.A(miu_data[6]));
   INV_X2 U81 (.ZN(U_rbuf_n188), 
	.A(miu_data[7]));
   INV_X2 U82 (.ZN(U_rbuf_n190), 
	.A(miu_data[9]));
   INV_X2 U83 (.ZN(U_rbuf_n191), 
	.A(miu_data[10]));
   INV_X2 U84 (.ZN(U_rbuf_n193), 
	.A(miu_data[12]));
   AND2_X2 U89 (.ZN(n50), 
	.A2(U_rbuf_f_top_data_13_), 
	.A1(U_rbuf_n145));
endmodule

module DW_memctl_miu (
	hclk, 
	hclk_2x, 
	hresetn, 
	scan_mode, 
	hiu_mem_req, 
	hiu_reg_req, 
	hiu_rw, 
	hiu_burst_size, 
	hiu_wrapped_burst, 
	hiu_terminate, 
	hiu_addr, 
	hiu_haddr, 
	hiu_hsize, 
	hiu_wr_data, 
	s_rd_data, 
	miu_burst_done, 
	miu_pop_n, 
	miu_push_n, 
	miu_col_addr_width, 
	miu_data_width, 
	m_addr, 
	s_addr, 
	s_bank_addr, 
	s_ras_n, 
	s_cas_n, 
	s_sel_n, 
	s_cke, 
	sf_cke, 
	s_we_n, 
	s_wr_data, 
	s_dqm, 
	s_dout_valid, 
	s_rd_ready, 
	s_rd_start, 
	s_rd_pop, 
	s_rd_end, 
	s_rd_dqs_mask, 
	s_cas_latency, 
	s_read_pipe, 
	sf_cas_latency, 
	s_sa, 
	s_scl, 
	s_dqs, 
	s_rp_n, 
	s_sda_out, 
	s_sda_in, 
	s_sda_oe_n, 
	sm_addr, 
	sm_oe_n, 
	sm_we_n, 
	sm_bs_n, 
	sm_dout_valid, 
	sm_rp_n, 
	sm_wp_n, 
	sm_adv_n, 
	sm_rd_data, 
	sm_wr_data, 
	remap, 
	sm_clken, 
	sm_ready, 
	sm_data_width_set0, 
	sm_access, 
	m_wr_data, 
	m_dout_valid, 
	m_precharge_bit, 
	s_ebi_req, 
	s_ebi_gnt, 
	sm_ebi_req, 
	sm_ebi_gnt, 
	power_down, 
	sf_power_down, 
	sm_power_down, 
	clear_sr_dp, 
	sf_clear_dp, 
	big_endian, 
	miu_rd_data_out, 
	gpi, 
	gpo, 
	debug_ad_bank_addr, 
	debug_ad_row_addr, 
	debug_ad_sf_bank_addr, 
	debug_ad_sf_row_addr, 
	debug_ad_sf_col_addr, 
	debug_sm_burst_done, 
	debug_sm_pop_n, 
	debug_sm_push_n, 
	debug_smc_cs, 
	debug_ref_req, 
	debug_ad_col_addr_15_, 
	debug_ad_col_addr_14_, 
	debug_ad_col_addr_11_, 
	debug_ad_col_addr_10_, 
	debug_ad_col_addr_9_, 
	debug_ad_col_addr_8_, 
	debug_ad_col_addr_7_, 
	debug_ad_col_addr_6_, 
	debug_ad_col_addr_5_, 
	debug_ad_col_addr_4_, 
	debug_ad_col_addr_3_, 
	debug_ad_col_addr_2_, 
	debug_ad_col_addr_1_, 
	debug_ad_col_addr_0_, 
	debug_ad_col_addr_13__BAR_BAR, 
	debug_ad_col_addr_12__BAR_BAR, 
	FE_OFN28_HRESETn, 
	FE_OFN31_HRESETn, 
	FE_OFN35_HRESETn, 
	FE_OFN46_HRESETn, 
	FE_OFN51_HRESETn, 
	FE_OFN53_HRESETn, 
	FE_OFN57_HRESETn, 
	HCLK__L5_N11, 
	HCLK__L5_N12, 
	HCLK__L5_N17, 
	HCLK__L5_N28, 
	HCLK__L5_N29, 
	HCLK__L5_N30, 
	HCLK__L5_N31, 
	HCLK__L5_N32, 
	HCLK__L5_N33, 
	HCLK__L5_N34, 
	HCLK__L5_N35, 
	HCLK__L5_N36, 
	HCLK__L5_N6, 
	FE_OFN151_HRESETn, 
	FE_OFN160_HRESETn, 
	FE_OFN191_HRESETn, 
	FE_OFN214_hiu_burst_size_4_, 
	FE_OFN217_hiu_burst_size_2_, 
	FE_OFN220_hiu_burst_size_0_);
   input hclk;
   input hclk_2x;
   input hresetn;
   input scan_mode;
   input hiu_mem_req;
   input hiu_reg_req;
   input hiu_rw;
   input [5:0] hiu_burst_size;
   input hiu_wrapped_burst;
   input hiu_terminate;
   input [31:0] hiu_addr;
   input [3:0] hiu_haddr;
   input [2:0] hiu_hsize;
   input [31:0] hiu_wr_data;
   input [31:0] s_rd_data;
   output miu_burst_done;
   output miu_pop_n;
   output miu_push_n;
   output [3:0] miu_col_addr_width;
   output [1:0] miu_data_width;
   output [15:0] m_addr;
   output [15:0] s_addr;
   output [1:0] s_bank_addr;
   output s_ras_n;
   output s_cas_n;
   output [0:0] s_sel_n;
   output s_cke;
   output sf_cke;
   output s_we_n;
   output [15:0] s_wr_data;
   output [1:0] s_dqm;
   output [1:0] s_dout_valid;
   input s_rd_ready;
   output s_rd_start;
   output s_rd_pop;
   output s_rd_end;
   output s_rd_dqs_mask;
   output [2:0] s_cas_latency;
   output [2:0] s_read_pipe;
   output [2:0] sf_cas_latency;
   output [2:0] s_sa;
   output s_scl;
   output [1:0] s_dqs;
   output s_rp_n;
   output s_sda_out;
   input s_sda_in;
   output s_sda_oe_n;
   output [22:0] sm_addr;
   output sm_oe_n;
   output sm_we_n;
   output [3:0] sm_bs_n;
   output [3:0] sm_dout_valid;
   output sm_rp_n;
   output [2:0] sm_wp_n;
   output sm_adv_n;
   input [31:0] sm_rd_data;
   output [31:0] sm_wr_data;
   input remap;
   input sm_clken;
   input sm_ready;
   input [2:0] sm_data_width_set0;
   output sm_access;
   output [15:0] m_wr_data;
   output [1:0] m_dout_valid;
   output m_precharge_bit;
   output s_ebi_req;
   input s_ebi_gnt;
   output sm_ebi_req;
   input sm_ebi_gnt;
   input power_down;
   input sf_power_down;
   input sm_power_down;
   input clear_sr_dp;
   input sf_clear_dp;
   input big_endian;
   output [31:0] miu_rd_data_out;
   input [7:0] gpi;
   output [7:0] gpo;
   output [1:0] debug_ad_bank_addr;
   output [15:0] debug_ad_row_addr;
   output [1:0] debug_ad_sf_bank_addr;
   output [15:0] debug_ad_sf_row_addr;
   output [15:0] debug_ad_sf_col_addr;
   output debug_sm_burst_done;
   output debug_sm_pop_n;
   output debug_sm_push_n;
   output [3:0] debug_smc_cs;
   output debug_ref_req;
   output debug_ad_col_addr_15_;
   output debug_ad_col_addr_14_;
   output debug_ad_col_addr_11_;
   output debug_ad_col_addr_10_;
   output debug_ad_col_addr_9_;
   output debug_ad_col_addr_8_;
   output debug_ad_col_addr_7_;
   output debug_ad_col_addr_6_;
   output debug_ad_col_addr_5_;
   output debug_ad_col_addr_4_;
   output debug_ad_col_addr_3_;
   output debug_ad_col_addr_2_;
   output debug_ad_col_addr_1_;
   output debug_ad_col_addr_0_;
   output debug_ad_col_addr_13__BAR_BAR;
   output debug_ad_col_addr_12__BAR_BAR;
   input FE_OFN28_HRESETn;
   input FE_OFN31_HRESETn;
   input FE_OFN35_HRESETn;
   input FE_OFN46_HRESETn;
   input FE_OFN51_HRESETn;
   input FE_OFN53_HRESETn;
   input FE_OFN57_HRESETn;
   input HCLK__L5_N11;
   input HCLK__L5_N12;
   input HCLK__L5_N17;
   input HCLK__L5_N28;
   input HCLK__L5_N29;
   input HCLK__L5_N30;
   input HCLK__L5_N31;
   input HCLK__L5_N32;
   input HCLK__L5_N33;
   input HCLK__L5_N34;
   input HCLK__L5_N35;
   input HCLK__L5_N36;
   input HCLK__L5_N6;
   input FE_OFN151_HRESETn;
   input FE_OFN160_HRESETn;
   input FE_OFN191_HRESETn;
   input FE_OFN214_hiu_burst_size_4_;
   input FE_OFN217_hiu_burst_size_2_;
   input FE_OFN220_hiu_burst_size_0_;

   // Internal wires
   wire FE_PHN5253_U_cr_N551;
   wire FE_PHN5237_U_cr_n455;
   wire FE_PHN5234_U_cr_N551;
   wire FE_PHN5176_U_dsdc_n1637;
   wire FE_PHN5174_U_dsdc_n1436;
   wire FE_PHN5171_n27;
   wire FE_PHN5144_U_dsdc_n226;
   wire FE_PHN5142_U_dsdc_n378;
   wire FE_PHN5112_U_cr_N556;
   wire FE_PHN5110_U_cr_N398;
   wire FE_PHN5102_U_addrdec_N133;
   wire FE_PHN5064_s_read_pipe_0_;
   wire FE_PHN5056_U_dsdc_n376;
   wire FE_PHN5047_U_dsdc_n228;
   wire FE_PHN5042_U_dsdc_N4228;
   wire FE_PHN5012_U_dsdc_n371;
   wire FE_PHN5011_U_cr_N559;
   wire FE_PHN4966_U_cr_n65;
   wire FE_PHN4962_U_dsdc_n230;
   wire FE_PHN4952_U_cr_n108;
   wire FE_PHN4938_U_dmc_n12;
   wire FE_PHN4934_U_refctl_count_next_1_;
   wire FE_PHN4922_U_cr_N564;
   wire FE_PHN4915_U_cr_n51;
   wire FE_PHN4914_U_cr_n59;
   wire FE_PHN4913_U_cr_N404;
   wire FE_PHN4894_U_cr_n48;
   wire FE_PHN4893_U_cr_N473;
   wire FE_PHN4878_U_dsdc_n366;
   wire FE_PHN4871_U_cr_n46;
   wire FE_PHN4855_U_cr_n49;
   wire FE_PHN4851_U_cr_N691;
   wire FE_PHN4849_U_cr_N395;
   wire FE_PHN4845_U_cr_n47;
   wire FE_PHN4842_U_cr_N636;
   wire FE_PHN4841_U_cr_N313;
   wire FE_PHN4818_U_cr_N469;
   wire FE_PHN4805_U_cr_N468;
   wire FE_PHN4798_U_cr_n50;
   wire FE_PHN4792_U_cr_N635;
   wire FE_PHN4787_U_cr_N736;
   wire FE_PHN4785_U_dsdc_N4229;
   wire FE_PHN4777_U_dsdc_n214;
   wire FE_PHN4776_U_cr_N558;
   wire FE_PHN4775_U_cr_N476;
   wire FE_PHN4763_U_cr_N479;
   wire FE_PHN4760_U_cr_N397;
   wire FE_PHN4759_U_cr_N745;
   wire FE_PHN4736_U_cr_N403;
   wire FE_PHN4728_U_cr_N551;
   wire FE_PHN4727_U_refctl_ref_req_next;
   wire FE_PHN4718_U_dsdc_n389;
   wire FE_PHN4717_U_dsdc_n268;
   wire FE_PHN4716_U_dsdc_n261;
   wire FE_PHN4715_U_dsdc_n276;
   wire FE_PHN4714_cr_t_xsr_1_;
   wire FE_PHN4713_U_dmc_data_cnt_nxt_5_;
   wire FE_PHN4678_U_dsdc_N4428;
   wire FE_PHN4676_U_dsdc_N4381;
   wire FE_PHN4645_U_cr_N302;
   wire FE_PHN4627_U_cr_N405;
   wire FE_PHN4625_U_dsdc_n1637;
   wire FE_PHN4623_U_dsdc_n1436;
   wire FE_PHN4620_U_cr_s_sda_d;
   wire FE_PHN4618_U_cr_n20;
   wire FE_PHN4617_U_cr_n18;
   wire FE_PHN4616_n27;
   wire FE_PHN4614_U_dsdc_n409;
   wire FE_PHN4613_U_dsdc_n386;
   wire FE_PHN4612_U_cr_n285;
   wire FE_PHN4610_U_dsdc_rcar_cnt1_nxt_0_;
   wire FE_PHN4609_U_cr_N301;
   wire FE_PHN4606_U_dsdc_N4347;
   wire FE_PHN4605_U_dsdc_N4339;
   wire FE_PHN4604_U_dsdc_N4341;
   wire FE_PHN4603_U_dsdc_n295;
   wire FE_PHN4600_U_dsdc_n393;
   wire FE_PHN4599_U_dsdc_n221;
   wire FE_PHN4598_U_dsdc_N4345;
   wire FE_PHN4594_U_cr_N409;
   wire FE_PHN4593_U_dsdc_N4337;
   wire FE_PHN4592_U_dsdc_n390;
   wire FE_PHN4591_U_dsdc_N4349;
   wire FE_PHN4589_U_cr_n286;
   wire FE_PHN4587_U_dsdc_N4140;
   wire FE_PHN4582_U_dsdc_n294;
   wire FE_PHN4581_U_dsdc_N4492;
   wire FE_PHN4578_U_dsdc_N4343;
   wire FE_PHN4574_U_cr_N563;
   wire FE_PHN4568_U_cr_N553;
   wire FE_PHN4558_U_dsdc_N4384;
   wire FE_PHN4551_U_dsdc_N4389;
   wire FE_PHN4547_U_dsdc_N4440;
   wire FE_PHN4546_U_dsdc_N4434;
   wire FE_PHN4543_U_refctl_count_next_0_;
   wire FE_PHN4542_U_dsdc_N4351;
   wire FE_PHN4537_U_dsdc_N4340;
   wire FE_PHN4530_U_dsdc_N4397;
   wire FE_PHN4528_U_dsdc_N4477;
   wire FE_PHN4527_U_dsdc_N4388;
   wire FE_PHN4522_U_dsdc_n300;
   wire FE_PHN4521_U_dsdc_N4436;
   wire FE_PHN4520_U_dsdc_N4433;
   wire FE_PHN4519_U_dsdc_N4336;
   wire FE_PHN4513_U_dsdc_N4383;
   wire FE_PHN4507_U_dsdc_N4444;
   wire FE_PHN4503_U_dsdc_N4473;
   wire FE_PHN4502_U_dsdc_N4442;
   wire FE_PHN4501_U_dsdc_N4431;
   wire FE_PHN4498_U_dsdc_N4481;
   wire FE_PHN4497_U_dsdc_wrapped_pop_flag_nxt;
   wire FE_PHN4491_U_dsdc_N4491;
   wire FE_PHN4489_U_dsdc_N4430;
   wire FE_PHN4483_U_cr_N638;
   wire FE_PHN4480_U_dsdc_N4441;
   wire FE_PHN4473_U_dsdc_N4482;
   wire FE_PHN4470_U_cr_N646;
   wire FE_PHN4469_U_dsdc_N4439;
   wire FE_PHN4465_U_dsdc_N4488;
   wire FE_PHN4464_U_cr_n19;
   wire FE_PHN4461_U_dsdc_N4350;
   wire FE_PHN4455_U_dsdc_N4395;
   wire FE_PHN4445_U_dsdc_N4479;
   wire FE_PHN4443_U_dsdc_N4435;
   wire FE_PHN4442_U_dsdc_N4438;
   wire FE_PHN4435_U_dsdc_N4478;
   wire FE_PHN4434_U_dsdc_N4398;
   wire FE_PHN4429_U_cr_N644;
   wire FE_PHN4428_U_cr_N692;
   wire FE_PHN4424_U_dsdc_N4342;
   wire FE_PHN4423_U_dsdc_N4487;
   wire FE_PHN4415_U_dsdc_N4391;
   wire FE_PHN4414_U_dsdc_N4386;
   wire FE_PHN4410_U_refctl_count_next_4_;
   wire FE_PHN4409_U_cr_N305;
   wire FE_PHN4408_U_dsdc_N4390;
   wire FE_PHN4398_U_cr_N303;
   wire FE_PHN4397_U_dsdc_n279;
   wire FE_PHN4395_U_dsdc_wtr_cnt_nxt_0_;
   wire FE_PHN4391_U_dsdc_n209;
   wire FE_PHN4390_U_dsdc_N4483;
   wire FE_PHN4389_U_dsdc_N4392;
   wire FE_PHN4388_U_dsdc_N4394;
   wire FE_PHN4381_U_dsdc_N4489;
   wire FE_PHN4365_U_dsdc_N4485;
   wire FE_PHN4360_U_cr_N640;
   wire FE_PHN4359_U_dsdc_N4445;
   wire FE_PHN4354_U_dsdc_N4385;
   wire FE_PHN4353_U_dsdc_N4338;
   wire FE_PHN4349_U_dsdc_N4480;
   wire FE_PHN4345_U_dsdc_N4486;
   wire FE_PHN4344_U_dsdc_N4344;
   wire FE_PHN4342_U_dsdc_N4393;
   wire FE_PHN4339_U_dsdc_N4437;
   wire FE_PHN4328_U_dsdc_N4443;
   wire FE_PHN4323_U_dsdc_N4346;
   wire FE_PHN4315_U_dsdc_N4348;
   wire FE_PHN4308_U_dsdc_n213;
   wire FE_PHN4307_U_dsdc_N4396;
   wire FE_PHN4306_U_dsdc_N4490;
   wire FE_PHN4304_U_dsdc_N4484;
   wire FE_PHN4293_U_dsdc_n293;
   wire FE_PHN4286_U_dsdc_N4432;
   wire FE_PHN4277_U_dsdc_N4387;
   wire FE_PHN4265_U_cr_n29;
   wire FE_PHN4246_U_dsdc_n356;
   wire FE_PHN4204_U_cr_N556;
   wire FE_PHN4152_s_read_pipe_0_;
   wire FE_PHN4110_U_cr_n53;
   wire FE_PHN4075_U_dsdc_n185;
   wire FE_PHN4045_U_cr_n46;
   wire FE_PHN4029_U_cr_N306;
   wire FE_PHN4013_U_cr_n108;
   wire FE_PHN4006_U_cr_n49;
   wire FE_PHN3988_U_cr_n60;
   wire FE_PHN3968_U_cr_n51;
   wire FE_PHN3951_U_dsdc_N4139;
   wire FE_PHN3938_U_cr_n48;
   wire FE_PHN3889_U_cr_n47;
   wire FE_PHN3876_U_cr_n50;
   wire FE_PHN3870_U_dmc_n12;
   wire FE_PHN3867_U_cr_N559;
   wire FE_PHN3844_U_cr_N472;
   wire FE_PHN3833_U_cr_N642;
   wire FE_PHN3831_U_cr_N696;
   wire FE_PHN3830_U_cr_N691;
   wire FE_PHN3826_U_cr_n83;
   wire FE_PHN3816_U_cr_N473;
   wire FE_PHN3810_U_cr_N636;
   wire FE_PHN3800_U_cr_N397;
   wire FE_PHN3786_U_cr_N469;
   wire FE_PHN3781_U_cr_N468;
   wire FE_PHN3777_U_cr_N697;
   wire FE_PHN3776_U_cr_N736;
   wire FE_PHN3771_U_cr_N635;
   wire FE_PHN3768_U_cr_N637;
   wire FE_PHN3766_U_cr_N402;
   wire FE_PHN3760_U_cr_N471;
   wire FE_PHN3759_U_cr_N394;
   wire FE_PHN3758_U_cr_N560;
   wire FE_PHN3757_U_cr_n82;
   wire FE_PHN3751_U_cr_N478;
   wire FE_PHN3745_U_cr_N558;
   wire FE_PHN3739_U_cr_N476;
   wire FE_PHN3738_U_cr_N474;
   wire FE_PHN3737_U_cr_N737;
   wire FE_PHN3736_U_cr_N645;
   wire FE_PHN3724_U_cr_N396;
   wire FE_PHN3722_U_cr_N699;
   wire FE_PHN3714_U_cr_N694;
   wire FE_PHN3713_U_cr_N299;
   wire FE_PHN3712_U_cr_N555;
   wire FE_PHN3707_U_cr_N479;
   wire FE_PHN3704_U_cr_n90;
   wire FE_PHN3702_U_cr_N695;
   wire FE_PHN3698_U_cr_N740;
   wire FE_PHN3697_U_cr_n89;
   wire FE_PHN3692_U_cr_N298;
   wire FE_PHN3687_U_cr_n91;
   wire FE_PHN3686_U_cr_N745;
   wire FE_PHN3684_U_cr_N643;
   wire FE_PHN3683_U_cr_N310;
   wire FE_PHN3680_U_cr_N693;
   wire FE_PHN3672_U_cr_n88;
   wire FE_PHN3669_U_cr_N477;
   wire FE_PHN3666_U_cr_N700;
   wire FE_PHN3665_U_cr_N470;
   wire FE_PHN3660_U_cr_N647;
   wire FE_PHN3659_U_cr_N639;
   wire FE_PHN3657_U_cr_N698;
   wire FE_PHN3651_U_cr_N554;
   wire FE_PHN3645_U_cr_N738;
   wire FE_PHN3643_U_cr_N641;
   wire FE_PHN3640_U_cr_N475;
   wire FE_PHN3638_U_cr_N739;
   wire FE_PHN3628_U_cr_n92;
   wire FE_PHN3619_U_cr_n94;
   wire FE_PHN3614_U_cr_N550;
   wire FE_PHN3613_U_dsdc_n405;
   wire FE_PHN3607_U_refctl_count_next_2_;
   wire FE_PHN3600_U_cr_n59;
   wire FE_PHN3588_U_cr_n149;
   wire FE_PHN3579_U_cr_N467;
   wire FE_PHN3575_U_cr_N401;
   wire FE_PHN3549_U_cr_n165;
   wire FE_PHN3515_U_cr_N551;
   wire FE_PHN3514_U_cr_n148;
   wire FE_PHN3513_U_dsdc_bm_ras_cnt_3__0_;
   wire FE_PHN3511_U_dsdc_bm_ras_cnt_0__0_;
   wire FE_PHN3510_U_dsdc_bm_ras_cnt_2__0_;
   wire FE_PHN3509_U_dsdc_bm_rc_cnt_2__0_;
   wire FE_PHN3508_U_dsdc_bm_rc_cnt_1__0_;
   wire FE_PHN3507_U_dsdc_bm_ras_cnt_1__0_;
   wire FE_PHN3505_U_cr_n45;
   wire FE_PHN3503_U_dsdc_rp_cnt1_nxt_0_;
   wire FE_PHN3485_U_cr_n77;
   wire FE_PHN3480_U_cr_n80;
   wire FE_PHN3479_U_cr_N404;
   wire FE_PHN3476_U_cr_n75;
   wire FE_PHN3475_U_cr_n74;
   wire FE_PHN3473_U_dsdc_n2095;
   wire FE_PHN3467_U_dsdc_n1924;
   wire FE_PHN3464_U_dsdc_n319;
   wire FE_PHN3463_U_dsdc_n1594;
   wire FE_PHN3461_U_dsdc_n394;
   wire FE_PHN3456_U_cr_N690;
   wire FE_PHN3454_U_dmc_n40;
   wire FE_PHN3452_U_dsdc_n410;
   wire FE_PHN3450_U_dsdc_wtr_cnt_nxt_1_;
   wire FE_PHN3449_U_refctl_next_state_0_;
   wire FE_PHN3446_U_dsdc_n269;
   wire FE_PHN3445_U_dsdc_n391;
   wire FE_PHN3443_U_dsdc_n282;
   wire FE_PHN3442_U_dsdc_n240;
   wire FE_PHN3440_U_dsdc_n265;
   wire FE_PHN3432_U_dsdc_n296;
   wire FE_PHN3431_U_dsdc_n256;
   wire FE_PHN3427_U_dsdc_rp_cnt2_nxt_2_;
   wire FE_PHN3415_U_dsdc_n266;
   wire FE_PHN3407_U_dsdc_n267;
   wire FE_PHN3399_U_dsdc_n412;
   wire FE_PHN3389_U_cr_N734;
   wire FE_PHN3379_U_cr_N733;
   wire FE_PHN3378_U_cr_N735;
   wire FE_PHN3373_U_addrdec_n347;
   wire FE_PHN3371_U_dsdc_n1231;
   wire FE_PHN3370_U_dsdc_n271;
   wire FE_PHN3355_U_dsdc_n406;
   wire FE_PHN3352_U_cr_n87;
   wire FE_PHN3349_U_cr_n86;
   wire FE_PHN3346_U_dsdc_n277;
   wire FE_PHN3345_U_dmc_n13;
   wire FE_PHN3343_U_refctl_count_next_3_;
   wire FE_PHN3337_U_dsdc_N4429;
   wire FE_PHN3328_U_dsdc_N4476;
   wire FE_PHN3327_U_dsdc_wr_cnt_nxt_0_;
   wire FE_PHN3326_U_refctl_count_next_15_;
   wire FE_PHN3325_U_dsdc_n262;
   wire FE_PHN3324_U_dsdc_num_init_ref_cnt_nxt_1_;
   wire FE_PHN3322_U_dsdc_n270;
   wire FE_PHN3321_U_dsdc_n263;
   wire FE_PHN3320_U_dsdc_n222;
   wire FE_PHN3319_U_dsdc_n255;
   wire FE_PHN3318_U_dsdc_n264;
   wire FE_PHN3317_U_dsdc_n259;
   wire FE_PHN3316_U_dsdc_n260;
   wire FE_PHN3315_U_dsdc_n211;
   wire FE_PHN3314_U_dsdc_n261;
   wire FE_PHN3313_U_dsdc_rp_cnt1_0_;
   wire FE_PHN3312_U_dsdc_n257;
   wire FE_PHN3311_U_dsdc_n268;
   wire FE_PHN3309_U_dsdc_cas_latency_cnt_2_;
   wire FE_PHN3305_U_refctl_count_next_1_;
   wire FE_PHN3299_U_dsdc_n274;
   wire FE_PHN3298_U_dsdc_n389;
   wire FE_PHN3297_U_dsdc_n283;
   wire FE_PHN3293_U_dsdc_n276;
   wire FE_PHN3292_cr_t_xsr_1_;
   wire FE_PHN3291_U_dmc_data_cnt_nxt_5_;
   wire FE_PHN3289_U_dsdc_n275;
   wire FE_PHN3288_U_dsdc_N4229;
   wire FE_PHN3287_U_cr_N576;
   wire FE_PHN3286_U_cr_n85;
   wire FE_PHN3283_cr_reg_data_out_24_;
   wire FE_PHN3268_U_dsdc_init_cnt_10_;
   wire FE_PHN3260_U_dsdc_n1212;
   wire FE_PHN3259_U_dsdc_n1205;
   wire FE_PHN3258_U_dsdc_n1184;
   wire FE_PHN3256_U_dsdc_n1198;
   wire FE_PHN3255_U_dsdc_n1241;
   wire FE_PHN3252_U_dsdc_n1191;
   wire FE_PHN3250_U_cr_N311;
   wire FE_PHN3249_U_cr_N312;
   wire FE_PHN3247_U_dsdc_n1177;
   wire FE_PHN3245_U_dsdc_N4462;
   wire FE_PHN3244_U_dsdc_n227;
   wire FE_PHN3242_U_dsdc_N4332;
   wire FE_PHN3241_U_dsdc_n212;
   wire FE_PHN3240_cr_t_rcar_2_;
   wire FE_PHN3239_U_dsdc_n230;
   wire FE_PHN3238_U_dsdc_rp_cnt1_nxt_1_;
   wire FE_PHN3237_U_cr_N562;
   wire FE_PHN3235_U_dsdc_n201;
   wire FE_PHN3234_U_dsdc_n228;
   wire FE_PHN3233_U_dsdc_n377;
   wire FE_PHN3232_U_dsdc_n370;
   wire FE_PHN3231_U_dsdc_n379;
   wire FE_PHN3230_U_cr_n81;
   wire FE_PHN3229_U_cr_n65;
   wire FE_PHN3228_U_dsdc_n368;
   wire FE_PHN3227_U_dsdc_n372;
   wire FE_PHN3224_U_cr_N410;
   wire FE_PHN3223_U_cr_N313;
   wire FE_PHN3222_U_dsdc_n375;
   wire FE_PHN3221_U_dsdc_n381;
   wire FE_PHN3220_U_cr_N408;
   wire FE_PHN3216_U_dsdc_n373;
   wire FE_PHN3215_U_cr_n76;
   wire FE_PHN3212_U_cr_n93;
   wire FE_PHN3208_U_dsdc_n2096;
   wire FE_PHN3197_U_dmc_n59;
   wire FE_PHN3196_U_cr_n99;
   wire FE_PHN3195_U_dsdc_n417;
   wire FE_PHN3194_U_dsdc_cas_cnt_nxt_3_;
   wire FE_PHN3193_U_dmc_n1;
   wire FE_PHN3192_U_cr_n128;
   wire FE_PHN3191_U_dsdc_n388;
   wire FE_PHN3189_U_dsdc_N4334;
   wire FE_PHN3188_U_addrdec_N119;
   wire FE_PHN3187_U_dsdc_rcar_cnt1_nxt_3_;
   wire FE_PHN3186_U_dsdc_num_init_ref_cnt_nxt_0_;
   wire FE_PHN3185_U_cr_n73;
   wire FE_PHN3183_U_dsdc_N4228;
   wire FE_PHN3182_U_dsdc_N4368;
   wire FE_PHN3170_U_dsdc_n371;
   wire FE_PHN3169_U_dsdc_n367;
   wire FE_PHN3168_U_dsdc_n380;
   wire FE_PHN3167_U_dsdc_n366;
   wire FE_PHN3166_U_dsdc_n374;
   wire FE_PHN3165_U_dsdc_n378;
   wire FE_PHN3164_U_addrdec_N130;
   wire FE_PHN3162_U_dsdc_n369;
   wire FE_PHN3160_U_dsdc_n423;
   wire FE_PHN3156_U_dsdc_n281;
   wire FE_PHN3127_U_dsdc_n414;
   wire FE_PHN3126_cr_block_size1_6_;
   wire FE_PHN3123_U_dsdc_n407;
   wire FE_PHN3119_U_dsdc_n411;
   wire FE_PHN3115_U_dsdc_n297;
   wire FE_PHN3113_U_cr_n63;
   wire FE_PHN3112_U_dsdc_n415;
   wire FE_PHN3111_cr_s_data_width_early_0_;
   wire FE_PHN3110_U_dsdc_num_init_ref_cnt_nxt_2_;
   wire FE_PHN3109_U_dsdc_N4415;
   wire FE_PHN3108_U_dsdc_N4321;
   wire FE_PHN3107_U_cr_n44;
   wire FE_PHN3106_U_cr_n43;
   wire FE_PHN3105_U_dsdc_n_2090_;
   wire FE_PHN3104_U_dsdc_N4174;
   wire FE_PHN3087_U_dsdc_cas_cnt_nxt_2_;
   wire FE_PHN3086_U_dsdc_n1275;
   wire FE_PHN3085_U_dsdc_rp_cnt2_nxt_0_;
   wire FE_PHN3083_U_dsdc_n280;
   wire FE_PHN3082_U_dsdc_n418;
   wire FE_PHN3081_U_dsdc_n416;
   wire FE_PHN3080_U_dsdc_n431;
   wire FE_PHN3079_U_dsdc_rcar_cnt2_nxt_3_;
   wire FE_PHN3077_U_dsdc_n460;
   wire FE_PHN3075_cr_push_n;
   wire FE_PHN3054_cr_row_addr_width_2_;
   wire FE_PHN3053_U_dsdc_n231;
   wire FE_PHN3052_U_cr_N302;
   wire FE_PHN3051_U_cr_N403;
   wire FE_PHN3049_U_refctl_ref_req_next;
   wire FE_PHN3047_U_dsdc_wr_cnt_nxt_2_;
   wire FE_PHN3046_ctl_sd_in_sf_mode;
   wire FE_PHN3045_U_dsdc_rp_cnt1_nxt_2_;
   wire FE_PHN3044_U_dsdc_n376;
   wire FE_PHN3043_U_cr_N413;
   wire FE_PHN3041_cr_t_init_0_;
   wire FE_PHN3034_U_dsdc_N4381;
   wire FE_PHN3033_U_dsdc_N4428;
   wire FE_PHN3031_n4;
   wire FE_PHN3030_n6;
   wire FE_PHN3029_n5;
   wire FE_PHN3028_U_dsdc_term_cnt_nxt_4_;
   wire FE_PHN3013_U_dsdc_N4475;
   wire FE_PHN3012_U_cr_n147;
   wire FE_PHN3011_U_dsdc_term_cnt_nxt_2_;
   wire FE_PHN2978_U_dsdc_N4141;
   wire FE_PHN2977_U_cr_N315;
   wire FE_PHN2975_U_dsdc_n216;
   wire FE_PHN2971_U_dsdc_n214;
   wire FE_PHN2964_U_cr_N405;
   wire FE_PHN2941_U_dsdc_term_cnt_nxt_0_;
   wire FE_PHN2929_cr_reg_data_out_15_;
   wire FE_PHN2915_U_cr_N566;
   wire FE_PHN2910_U_dsdc_n1637;
   wire FE_PHN2909_U_dsdc_n1436;
   wire FE_PHN2905_U_cr_s_sda_d;
   wire FE_PHN2455_U_cr_n20;
   wire FE_PHN2432_n27;
   wire FE_PHN2431_U_addrdec_N129;
   wire FE_PHN2427_U_addrdec_n347;
   wire FE_PHN2425_U_dsdc_N4341;
   wire FE_PHN2424_U_dsdc_N4347;
   wire FE_PHN2423_U_dsdc_N4345;
   wire FE_PHN2422_U_addrdec_n348;
   wire FE_PHN2419_U_dsdc_N4343;
   wire FE_PHN2418_U_dsdc_N4440;
   wire FE_PHN2417_U_dsdc_N4477;
   wire FE_PHN2416_U_dsdc_N4492;
   wire FE_PHN2414_U_dsdc_N4389;
   wire FE_PHN2413_U_dsdc_N4397;
   wire FE_PHN2411_U_dsdc_N4430;
   wire FE_PHN2410_U_dsdc_N4336;
   wire FE_PHN2409_U_dsdc_N4491;
   wire FE_PHN2408_U_dsdc_N4351;
   wire FE_PHN2407_U_dsdc_N4433;
   wire FE_PHN2406_U_dsdc_N4444;
   wire FE_PHN2405_U_dsdc_N4438;
   wire FE_PHN2404_U_dsdc_N4388;
   wire FE_PHN2402_U_dsdc_N4483;
   wire FE_PHN2401_U_dsdc_N4342;
   wire FE_PHN2400_U_dsdc_N4488;
   wire FE_PHN2399_U_dsdc_N4384;
   wire FE_PHN2398_U_dsdc_N4391;
   wire FE_PHN2397_U_dsdc_N4480;
   wire FE_PHN2396_U_dsdc_N4386;
   wire FE_PHN2395_U_dsdc_N4395;
   wire FE_PHN2394_U_dsdc_N4390;
   wire FE_PHN2393_U_dsdc_N4478;
   wire FE_PHN2392_U_dsdc_N4392;
   wire FE_PHN2391_U_dsdc_N4385;
   wire FE_PHN2390_U_dsdc_N4437;
   wire FE_PHN2389_U_dsdc_N4432;
   wire FE_PHN2388_U_dsdc_N4338;
   wire FE_PHN2387_U_dsdc_N4486;
   wire FE_PHN2386_U_dsdc_N4396;
   wire FE_PHN2384_U_dsdc_N4393;
   wire FE_PHN2383_U_dsdc_N4443;
   wire FE_PHN2382_U_dsdc_N4344;
   wire FE_PHN2381_U_dsdc_N4348;
   wire FE_PHN2380_U_dsdc_N4490;
   wire FE_PHN2377_U_dsdc_N4366;
   wire FE_PHN2373_U_dsdc_N4387;
   wire FE_PHN2146_U_addrdec_N131;
   wire FE_PHN2051_U_cr_n18;
   wire FE_PHN2044_U_dsdc_n273;
   wire FE_PHN2040_U_dsdc_n271;
   wire FE_PHN2038_U_dsdc_n277;
   wire FE_PHN2037_U_dsdc_rcar_cnt1_nxt_0_;
   wire FE_PHN2036_U_dsdc_cas_latency_cnt_0_;
   wire FE_PHN2034_U_dsdc_bm_ras_cnt_max_0_;
   wire FE_PHN2033_U_dsdc_n262;
   wire FE_PHN2032_U_dsdc_n270;
   wire FE_PHN2031_U_dsdc_n264;
   wire FE_PHN2030_U_dsdc_n255;
   wire FE_PHN2029_U_dsdc_n263;
   wire FE_PHN2027_U_dsdc_n268;
   wire FE_PHN2025_U_addrdec_N107;
   wire FE_PHN1921_U_dsdc_n1084;
   wire FE_PHN1918_U_cr_n285;
   wire FE_PHN1917_U_cr_N304;
   wire FE_PHN1916_U_cr_N556;
   wire FE_PHN1913_U_cr_N389;
   wire FE_PHN1911_U_cr_N399;
   wire FE_PHN1897_U_dsdc_n1002;
   wire FE_PHN1896_U_dsdc_r_burst_size_1_;
   wire FE_PHN1895_U_dsdc_n996;
   wire FE_PHN1893_U_dsdc_n1392;
   wire FE_PHN1892_U_dsdc_r_burst_size_3_;
   wire FE_PHN1891_U_dsdc_bm_ras_cnt_3__2_;
   wire FE_PHN1890_U_dsdc_r_burst_size_5_;
   wire FE_PHN1889_U_dsdc_bm_ras_cnt_1__2_;
   wire FE_PHN1888_U_dsdc_r_burst_size_4_;
   wire FE_PHN1887_U_dsdc_n166;
   wire FE_PHN1868_U_addrdec_n309;
   wire FE_PHN1855_cr_block_size1_7_;
   wire FE_PHN1854_U_addrdec_n346;
   wire FE_PHN1848_U_cr_N464;
   wire FE_PHN1845_U_cr_N465;
   wire FE_PHN1747_U_cr_N555;
   wire FE_PHN1746_U_cr_N554;
   wire FE_PHN1745_U_cr_N557;
   wire FE_PHN1740_U_cr_N564;
   wire FE_PHN1739_U_cr_N392;
   wire FE_PHN1738_U_cr_N402;
   wire FE_PHN1737_U_cr_N390;
   wire FE_PHN1736_U_cr_N394;
   wire FE_PHN1735_U_cr_N395;
   wire FE_PHN1734_U_cr_N396;
   wire FE_PHN1733_U_cr_N563;
   wire FE_PHN1732_U_cr_N479;
   wire FE_PHN1731_U_cr_N560;
   wire FE_PHN1730_U_cr_N472;
   wire FE_PHN1729_U_cr_N397;
   wire FE_PHN1728_U_cr_N475;
   wire FE_PHN1727_U_cr_N473;
   wire FE_PHN1726_U_cr_N558;
   wire FE_PHN1725_U_cr_N400;
   wire FE_PHN1724_U_cr_N398;
   wire FE_PHN1723_U_cr_N644;
   wire FE_PHN1722_U_cr_N647;
   wire FE_PHN1721_U_cr_N641;
   wire FE_PHN1720_U_cr_N643;
   wire FE_PHN1719_U_cr_N476;
   wire FE_PHN1718_U_cr_N640;
   wire FE_PHN1716_U_cr_n82;
   wire FE_PHN1715_U_cr_N642;
   wire FE_PHN1714_U_cr_N635;
   wire FE_PHN1713_U_cr_N636;
   wire FE_PHN1712_U_cr_N738;
   wire FE_PHN1711_U_cr_N471;
   wire FE_PHN1710_U_cr_n83;
   wire FE_PHN1709_U_cr_N739;
   wire FE_PHN1708_U_cr_N468;
   wire FE_PHN1707_U_cr_N740;
   wire FE_PHN1706_U_cr_N301;
   wire FE_PHN1705_U_cr_N470;
   wire FE_PHN1704_U_cr_N469;
   wire FE_PHN1703_U_cr_N691;
   wire FE_PHN1702_U_cr_N693;
   wire FE_PHN1701_U_cr_N737;
   wire FE_PHN1700_U_cr_N300;
   wire FE_PHN1699_U_cr_N299;
   wire FE_PHN1698_U_cr_N696;
   wire FE_PHN1697_U_cr_N697;
   wire FE_PHN1696_U_cr_N698;
   wire FE_PHN1695_U_cr_N700;
   wire FE_PHN1694_U_cr_n89;
   wire FE_PHN1693_U_cr_n91;
   wire FE_PHN1692_U_cr_N745;
   wire FE_PHN1690_U_cr_n92;
   wire FE_PHN1683_U_dsdc_N4229;
   wire FE_PHN1663_U_refctl_count_0_;
   wire FE_PHN1662_U_addrdec_n58;
   wire FE_PHN1661_U_cr_N574;
   wire FE_PHN1659_U_dsdc_n386;
   wire FE_PHN1658_U_dsdc_n403;
   wire FE_PHN1656_U_cr_N577;
   wire FE_PHN1647_U_cr_n86;
   wire FE_PHN1645_U_cr_n65;
   wire FE_PHN1643_U_cr_N688;
   wire FE_PHN1642_U_cr_n119;
   wire FE_PHN1641_U_addrdec_n345;
   wire FE_PHN1640_U_cr_N576;
   wire FE_PHN1639_U_cr_N733;
   wire FE_PHN1638_U_cr_N689;
   wire FE_PHN1637_U_cr_N734;
   wire FE_PHN1634_U_cr_n167;
   wire FE_PHN1628_U_cr_n286;
   wire FE_PHN1623_U_dsdc_n366;
   wire FE_PHN1617_U_cr_N406;
   wire FE_PHN1608_cr_reg_data_out_18_;
   wire FE_PHN1597_U_dmc_n1;
   wire FE_PHN1596_U_dsdc_n1091;
   wire FE_PHN1594_U_addrdec_N133;
   wire FE_PHN1593_U_dsdc_bm_bank_status_1_;
   wire FE_PHN1590_U_dsdc_N4322;
   wire FE_PHN1589_U_cr_N552;
   wire FE_PHN1587_U_cr_N391;
   wire FE_PHN1585_U_dsdc_n1094;
   wire FE_PHN1583_U_refctl_n80;
   wire FE_PHN1582_U_dsdc_N4340;
   wire FE_PHN1581_U_dsdc_N4482;
   wire FE_PHN1580_U_dsdc_N4436;
   wire FE_PHN1578_U_dsdc_N4434;
   wire FE_PHN1576_U_dsdc_N4481;
   wire FE_PHN1575_U_dsdc_N4435;
   wire FE_PHN1574_U_refctl_n78;
   wire FE_PHN1573_U_dsdc_N4487;
   wire FE_PHN1572_U_dsdc_N4485;
   wire FE_PHN1570_U_dsdc_N4346;
   wire FE_PHN1569_U_cr_N735;
   wire FE_PHN1568_U_cr_N466;
   wire FE_PHN1567_U_cr_N690;
   wire FE_PHN1557_U_refctl_count_next_1_;
   wire FE_PHN1555_U_cr_N571;
   wire FE_PHN1549_U_refctl_n89;
   wire FE_PHN1548_U_refctl_n85;
   wire FE_PHN1537_U_cr_N553;
   wire FE_PHN1536_U_cr_N478;
   wire FE_PHN1535_U_cr_N477;
   wire FE_PHN1534_U_cr_N637;
   wire FE_PHN1533_U_cr_N639;
   wire FE_PHN1532_U_cr_N638;
   wire FE_PHN1531_U_cr_N694;
   wire FE_PHN1530_U_cr_N695;
   wire FE_PHN1529_U_dsdc_n215;
   wire FE_PHN1528_U_cr_n88;
   wire FE_PHN1526_U_cr_N407;
   wire FE_PHN1524_U_cr_N408;
   wire FE_PHN1523_U_cr_N409;
   wire FE_PHN1522_U_cr_n94;
   wire FE_PHN1521_U_dsdc_n423;
   wire FE_PHN1520_U_cr_n75;
   wire FE_PHN1519_U_cr_n74;
   wire FE_PHN1518_U_cr_n76;
   wire FE_PHN1517_U_cr_n78;
   wire FE_PHN1516_U_cr_n79;
   wire FE_PHN1514_U_cr_N311;
   wire FE_PHN1504_U_cr_N551;
   wire FE_PHN1497_U_dsdc_n1238;
   wire FE_PHN1496_U_dsdc_N4369;
   wire FE_PHN1495_U_dsdc_N4416;
   wire FE_PHN1494_U_refctl_next_state_0_;
   wire FE_PHN1493_U_dsdc_n282;
   wire FE_PHN1492_U_dsdc_n1180;
   wire FE_PHN1491_U_dsdc_N4140;
   wire FE_PHN1489_U_dsdc_N4429;
   wire FE_PHN1487_U_dsdc_n1194;
   wire FE_PHN1486_U_dsdc_N4476;
   wire FE_PHN1485_U_dsdc_N4442;
   wire FE_PHN1484_U_dsdc_n319;
   wire FE_PHN1483_U_dsdc_n280;
   wire FE_PHN1482_U_cr_n151;
   wire FE_PHN1481_U_dsdc_N4489;
   wire FE_PHN1480_U_dsdc_n259;
   wire FE_PHN1479_U_dsdc_n260;
   wire FE_PHN1478_U_dsdc_n261;
   wire FE_PHN1477_U_cr_stmg0r_0_;
   wire FE_PHN1476_U_refctl_count_next_15_;
   wire FE_PHN1475_cr_s_data_width_early_0_;
   wire FE_PHN1473_U_cr_n27;
   wire FE_PHN1470_U_dsdc_write_start_nxt;
   wire FE_PHN1456_U_cr_N310;
   wire FE_PHN1455_U_cr_N303;
   wire FE_PHN1449_U_cr_N561;
   wire FE_PHN1447_U_dsdc_N429;
   wire FE_PHN1445_U_dsdc_n157;
   wire FE_PHN1444_U_cr_N646;
   wire FE_PHN1430_U_dsdc_N4228;
   wire FE_PHN1427_cr_reg_data_out_17_;
   wire FE_PHN1424_U_refctl_count_12_;
   wire FE_PHN1421_U_refctl_count_10_;
   wire FE_PHN1420_U_refctl_count_8_;
   wire FE_PHN1419_U_refctl_count_6_;
   wire FE_PHN1418_U_dmc_data_cnt_2_;
   wire FE_PHN1416_U_dsdc_r_col_addr_1_;
   wire FE_PHN1415_U_refctl_n86;
   wire FE_PHN1414_U_refctl_count_next_14_;
   wire FE_PHN1413_U_dsdc_N4281;
   wire FE_PHN1412_U_cr_N634;
   wire FE_PHN1411_U_refctl_n91;
   wire FE_PHN1410_U_dsdc_N4413;
   wire FE_PHN1409_U_cr_n85;
   wire FE_PHN1407_U_cr_n104;
   wire FE_PHN1403_U_refctl_count_next_5_;
   wire FE_PHN1402_U_dsdc_n1462;
   wire FE_PHN1401_U_cr_cr_cs_1_;
   wire FE_PHN1400_U_cr_n197;
   wire FE_PHN1388_U_cr_N393;
   wire FE_PHN1387_U_cr_N401;
   wire FE_PHN1386_U_cr_N474;
   wire FE_PHN1384_U_cr_N467;
   wire FE_PHN1383_U_cr_N736;
   wire FE_PHN1382_U_cr_N692;
   wire FE_PHN1381_U_dsdc_wr_cnt_nxt_1_;
   wire FE_PHN1380_U_cr_N699;
   wire FE_PHN1378_U_cr_n90;
   wire FE_PHN1376_U_cr_N648;
   wire FE_PHN1375_U_cr_N649;
   wire FE_PHN1372_cr_reg_data_out_26_;
   wire FE_PHN1371_cr_reg_data_out_19_;
   wire FE_PHN1369_cr_reg_data_out_23_;
   wire FE_PHN1343_U_dsdc_n1276;
   wire FE_PHN1340_U_dmc_data_cnt_nxt_1_;
   wire FE_PHN1338_U_dsdc_cas_cnt_nxt_5_;
   wire FE_PHN1337_U_dsdc_n363;
   wire FE_PHN1336_U_dsdc_n364;
   wire FE_PHN1335_U_dsdc_n1281;
   wire FE_PHN1334_U_dsdc_n365;
   wire FE_PHN1333_U_dsdc_n382;
   wire FE_PHN1329_U_dsdc_N4339;
   wire FE_PHN1328_U_dsdc_n417;
   wire FE_PHN1326_U_dsdc_n258;
   wire FE_PHN1323_U_dsdc_n393;
   wire FE_PHN1322_U_dsdc_N4337;
   wire FE_PHN1321_U_dsdc_n390;
   wire FE_PHN1315_U_dsdc_N4414;
   wire FE_PHN1311_U_dsdc_N4427;
   wire FE_PHN1310_U_dsdc_N4474;
   wire FE_PHN1306_U_dsdc_N4380;
   wire FE_PHN1303_U_dsdc_N4383;
   wire FE_PHN1300_U_dsdc_N4439;
   wire FE_PHN1299_U_dsdc_N4350;
   wire FE_PHN1295_U_dsdc_n418;
   wire FE_PHN1294_U_dsdc_N4333;
   wire FE_PHN1292_U_dsdc_N4479;
   wire FE_PHN1291_U_dsdc_N4431;
   wire FE_PHN1288_U_dsdc_N4319;
   wire FE_PHN1287_U_dsdc_N4473;
   wire FE_PHN1279_U_dsdc_N4484;
   wire FE_PHN1275_U_dsdc_N4426;
   wire FE_PHN1271_U_dsdc_N4379;
   wire FE_PHN1269_U_dsdc_n257;
   wire FE_PHN1268_U_dsdc_N4332;
   wire FE_PHN1262_U_dsdc_N4139;
   wire FE_PHN1256_U_cr_N573;
   wire FE_PHN1254_U_cr_n55;
   wire FE_PHN1253_U_cr_N306;
   wire FE_PHN1252_U_cr_N307;
   wire FE_PHN1251_U_refctl_ref_req_next;
   wire FE_PHN1249_U_dsdc_add_x_2600_1_n8;
   wire FE_PHN1247_U_dsdc_n373;
   wire FE_PHN1243_U_cr_N655;
   wire FE_PHN1242_U_dsdc_wtr_cnt_nxt_1_;
   wire FE_PHN1240_U_cr_N312;
   wire FE_PHN1236_cr_reg_data_out_25_;
   wire FE_PHN1235_cr_reg_data_out_5_;
   wire FE_PHN1234_cr_reg_data_out_4_;
   wire FE_PHN1230_cr_reg_data_out_11_;
   wire FE_PHN1228_U_dmc_data_cnt_3_;
   wire FE_PHN1227_U_dsdc_cas_cnt_2_;
   wire FE_PHN1224_ctl_sd_in_sf_mode;
   wire FE_PHN1222_U_dsdc_bm_rc_cnt_2__2_;
   wire FE_PHN1221_U_dsdc_bm_rc_cnt_1__2_;
   wire FE_PHN1220_U_dsdc_n407;
   wire FE_PHN1219_U_dsdc_bm_rc_cnt_3__2_;
   wire FE_PHN1218_U_dsdc_cas_cnt_nxt_1_;
   wire FE_PHN1217_U_dmc_data_cnt_nxt_2_;
   wire FE_PHN1216_U_dsdc_n413;
   wire FE_PHN1215_U_dsdc_n409;
   wire FE_PHN1214_U_dsdc_n411;
   wire FE_PHN1213_U_dsdc_rcar_cnt2_nxt_0_;
   wire FE_PHN1212_U_dsdc_cas_latency_cnt_1_;
   wire FE_PHN1211_U_dmc_data_cnt_nxt_5_;
   wire FE_PHN1210_U_dsdc_n388;
   wire FE_PHN1209_U_dsdc_N4349;
   wire FE_PHN1208_U_dsdc_rcar_cnt1_nxt_1_;
   wire FE_PHN1207_U_refctl_count_next_11_;
   wire FE_PHN1206_U_dsdc_N4398;
   wire FE_PHN1205_U_dsdc_N4441;
   wire FE_PHN1204_U_dsdc_N4445;
   wire FE_PHN1203_U_refctl_count_next_9_;
   wire FE_PHN1202_U_dsdc_N4394;
   wire FE_PHN1201_U_refctl_count_next_13_;
   wire FE_PHN1200_U_dsdc_n1161;
   wire FE_PHN1199_U_dsdc_rp_cnt1_nxt_2_;
   wire FE_PHN1198_U_dsdc_rp_cnt1_nxt_0_;
   wire FE_PHN1185_U_refctl_count_next_7_;
   wire FE_PHN1176_U_cr_n84;
   wire FE_PHN1173_U_dsdc_wr_cnt_nxt_0_;
   wire FE_PHN1171_U_cr_n297;
   wire FE_PHN1170_U_cr_N313;
   wire FE_PHN1169_cr_reg_data_out_24_;
   wire FE_PHN1168_U_cr_N413;
   wire FE_PHN1167_cr_reg_data_out_1_;
   wire FE_PHN1166_cr_reg_data_out_29_;
   wire FE_PHN1165_cr_reg_data_out_14_;
   wire FE_PHN1163_U_cr_n482;
   wire FE_PHN1161_U_dsdc_n1339;
   wire FE_PHN1160_U_dmc_n48;
   wire FE_PHN1158_U_dsdc_bm_ras_cnt_max_1_;
   wire FE_PHN1156_U_dsdc_n1182;
   wire FE_PHN1155_U_dsdc_n1210;
   wire FE_PHN1154_U_dsdc_n1196;
   wire FE_PHN1153_U_dsdc_cas_latency_cnt_3_;
   wire FE_PHN1152_U_dsdc_r_row_addr_5_;
   wire FE_PHN1151_U_dsdc_r_row_addr_8_;
   wire FE_PHN1150_U_cr_sctlr_14_;
   wire FE_PHN1149_U_dsdc_r_row_addr_12_;
   wire FE_PHN1148_U_dsdc_r_row_addr_10_;
   wire FE_PHN1147_U_dsdc_r_row_addr_4_;
   wire FE_PHN1146_U_dsdc_r_row_addr_6_;
   wire FE_PHN1144_U_dsdc_wrapped_pop_flag_nxt;
   wire FE_PHN1143_U_dsdc_num_init_ref_cnt_nxt_2_;
   wire FE_PHN1140_U_refctl_count_next_2_;
   wire FE_PHN1127_U_cr_N305;
   wire FE_PHN1124_U_cr_N645;
   wire FE_PHN1123_U_dsdc_n372;
   wire FE_PHN1122_U_dsdc_n371;
   wire FE_PHN1121_U_dsdc_n367;
   wire FE_PHN1120_U_dsdc_n369;
   wire FE_PHN1119_U_cr_N653;
   wire FE_PHN1118_U_cr_N654;
   wire FE_PHN1117_cr_reg_data_out_20_;
   wire FE_PHN1116_U_cr_N415;
   wire FE_PHN1103_U_cr_n455;
   wire FE_PHN1101_U_dsdc_n1275;
   wire FE_PHN1099_U_dsdc_n404;
   wire FE_PHN1098_U_dsdc_N4334;
   wire FE_PHN1097_U_dsdc_N4428;
   wire FE_PHN1096_U_dsdc_N4381;
   wire FE_PHN1095_U_dsdc_n392;
   wire FE_PHN1094_U_dsdc_n394;
   wire FE_PHN1093_U_dsdc_n340;
   wire FE_PHN1092_U_dsdc_N4128;
   wire FE_PHN1091_U_refctl_count_next_3_;
   wire FE_PHN1090_U_dsdc_N4460;
   wire FE_PHN1089_U_refctl_count_next_4_;
   wire FE_PHN1088_U_cr_n558;
   wire FE_PHN1087_U_dsdc_rp_cnt1_nxt_1_;
   wire FE_PHN1083_U_cr_N650;
   wire FE_PHN1082_U_cr_n77;
   wire FE_PHN1081_U_dsdc_n1671;
   wire FE_PHN1080_cr_reg_data_out_0_;
   wire FE_PHN1077_cr_reg_data_out_22_;
   wire FE_PHN1076_U_cr_N418;
   wire FE_PHN1064_cr_row_addr_width_3_;
   wire FE_PHN1062_U_dsdc_init_cnt_3_;
   wire FE_PHN1061_U_dsdc_N4475;
   wire FE_PHN1060_U_dsdc_N4321;
   wire FE_PHN1059_U_dsdc_N4462;
   wire FE_PHN1058_U_dsdc_N4141;
   wire FE_PHN1057_U_dsdc_N4415;
   wire FE_PHN1056_U_dmc_terminate;
   wire FE_PHN1055_U_dsdc_N4368;
   wire FE_PHN1054_U_dsdc_rp_cnt2_nxt_0_;
   wire FE_PHN1053_U_dsdc_rcar_cnt1_nxt_3_;
   wire FE_PHN1052_U_cr_n127;
   wire FE_PHN1051_U_dsdc_rcar_cnt1_nxt_2_;
   wire FE_PHN1050_U_dsdc_n218;
   wire FE_PHN1048_U_cr_N550;
   wire FE_PHN1047_U_dsdc_n405;
   wire FE_PHN1046_U_dsdc_n380;
   wire FE_PHN1045_U_dsdc_n376;
   wire FE_PHN1044_U_cr_N652;
   wire FE_PHN1043_U_cr_N412;
   wire FE_PHN1042_cr_reg_data_out_28_;
   wire FE_PHN1041_cr_reg_data_out_2_;
   wire FE_PHN1040_U_cr_N419;
   wire FE_PHN1035_U_dsdc_n327;
   wire FE_PHN1034_cr_bank_addr_width_1_;
   wire FE_PHN1033_U_dsdc_xsr_cnt_1_;
   wire FE_PHN1032_U_dsdc_init_cnt_9_;
   wire FE_PHN1031_U_dsdc_init_cnt_7_;
   wire FE_PHN1030_U_dsdc_xsr_cnt_3_;
   wire FE_PHN1029_U_dsdc_n414;
   wire FE_PHN1028_U_dsdc_N4127;
   wire FE_PHN1026_U_dsdc_N4367;
   wire FE_PHN1023_U_dsdc_n387;
   wire FE_PHN1020_U_dsdc_n1085;
   wire FE_PHN1017_U_cr_N651;
   wire FE_PHN1016_U_dsdc_n281;
   wire FE_PHN1015_U_cr_n295;
   wire FE_PHN1014_U_cr_N567;
   wire FE_PHN1013_U_cr_n73;
   wire FE_PHN1012_U_dsdc_n_2088_;
   wire FE_PHN1001_U_dsdc_n391;
   wire FE_PHN1000_U_dmc_n14;
   wire FE_PHN998_U_dsdc_n221;
   wire FE_PHN997_U_dsdc_N4320;
   wire FE_PHN996_U_dsdc_num_init_ref_cnt_nxt_0_;
   wire FE_PHN995_U_dsdc_N4283;
   wire FE_PHN994_U_dsdc_n212;
   wire FE_PHN992_U_dsdc_n209;
   wire FE_PHN990_U_dsdc_n_2089_;
   wire FE_PHN989_U_dsdc_n214;
   wire FE_PHN988_U_cr_N298;
   wire FE_PHN987_U_dsdc_n370;
   wire FE_PHN986_U_dsdc_n368;
   wire FE_PHN985_U_dsdc_n377;
   wire FE_PHN984_U_dsdc_n381;
   wire FE_PHN983_U_dsdc_n378;
   wire FE_PHN982_U_cr_n93;
   wire FE_PHN981_U_dsdc_n329;
   wire FE_PHN980_cr_reg_data_out_16_;
   wire FE_PHN979_cr_reg_data_out_30_;
   wire FE_PHN978_U_cr_N416;
   wire FE_PHN977_U_cr_N417;
   wire FE_PHN971_U_dsdc_init_cnt_5_;
   wire FE_PHN970_U_dsdc_init_cnt_11_;
   wire FE_PHN969_U_dsdc_n1727;
   wire FE_PHN968_U_dsdc_n415;
   wire FE_PHN967_U_dmc_n4;
   wire FE_PHN966_U_dsdc_n416;
   wire FE_PHN964_U_dsdc_n431;
   wire FE_PHN961_U_dsdc_n231;
   wire FE_PHN960_U_dsdc_rcar_cnt2_nxt_3_;
   wire FE_PHN959_U_dsdc_n226;
   wire FE_PHN958_U_dsdc_n353;
   wire FE_PHN957_U_cr_N559;
   wire FE_PHN955_s_read_pipe_1_;
   wire FE_PHN953_U_dsdc_n375;
   wire FE_PHN952_U_cr_N410;
   wire FE_PHN951_U_dsdc_n216;
   wire FE_PHN949_cr_reg_data_out_21_;
   wire FE_PHN948_U_cr_n442;
   wire FE_PHN945_U_dsdc_n1175;
   wire FE_PHN944_U_dmc_n54;
   wire FE_PHN943_U_dmc_n7;
   wire FE_PHN942_U_dsdc_n408;
   wire FE_PHN940_U_dsdc_n294;
   wire FE_PHN938_U_dsdc_n406;
   wire FE_PHN937_U_dsdc_n297;
   wire FE_PHN934_U_dsdc_n_2090_;
   wire FE_PHN933_U_dsdc_wtr_cnt_nxt_0_;
   wire FE_PHN932_U_cr_N315;
   wire FE_PHN931_U_dsdc_n2094;
   wire FE_PHN927_U_addrdec_N108;
   wire FE_PHN926_U_cr_n98;
   wire FE_PHN925_U_dsdc_n410;
   wire FE_PHN924_U_dsdc_rp_cnt2_nxt_2_;
   wire FE_PHN922_U_dsdc_n412;
   wire FE_PHN921_U_dsdc_N4461;
   wire FE_PHN918_cr_bank_addr_width_0_;
   wire FE_PHN917_U_dsdc_n223;
   wire FE_PHN916_U_cr_cr_cs_2_;
   wire FE_PHN907_U_dsdc_cas_latency_1_;
   wire FE_PHN906_U_dsdc_n379;
   wire FE_PHN905_U_dsdc_n374;
   wire FE_PHN902_U_dmc_data_cnt_4_;
   wire FE_PHN901_U_dsdc_n295;
   wire FE_PHN900_U_dsdc_rcar_cnt2_nxt_1_;
   wire FE_PHN899_U_dsdc_n227;
   wire FE_PHN898_U_dsdc_n213;
   wire FE_PHN897_U_dsdc_n352;
   wire FE_PHN896_U_dsdc_n389;
   wire FE_PHN895_U_dsdc_n283;
   wire FE_PHN894_U_dsdc_n1464;
   wire FE_PHN893_U_dsdc_n1092;
   wire FE_PHN891_U_dsdc_wr_cnt_nxt_2_;
   wire FE_PHN889_U_cr_N411;
   wire FE_PHN887_n4;
   wire FE_PHN886_n6;
   wire FE_PHN884_n1;
   wire FE_PHN883_n2;
   wire FE_PHN882_U_dsdc_n2097;
   wire FE_PHN881_n3;
   wire FE_PHN880_cr_reg_data_out_12_;
   wire FE_PHN866_U_dmc_n13;
   wire FE_PHN865_U_dsdc_n296;
   wire FE_PHN864_U_dsdc_n222;
   wire FE_PHN863_U_dsdc_n211;
   wire FE_PHN862_U_dsdc_n230;
   wire FE_PHN855_cr_reg_data_out_8_;
   wire FE_PHN854_U_dsdc_n2093;
   wire FE_PHN853_cr_reg_data_out_13_;
   wire FE_PHN850_cr_reg_data_out_7_;
   wire FE_PHN843_U_dsdc_num_init_ref_cnt_1_;
   wire FE_PHN842_U_dsdc_n220;
   wire FE_PHN841_U_dsdc_bm_ras_cnt_max_3_;
   wire FE_PHN840_U_cr_n99;
   wire FE_PHN838_U_dsdc_rp_cnt2_nxt_1_;
   wire FE_PHN837_U_cr_cr_cs_0_;
   wire FE_PHN836_U_dsdc_n287;
   wire FE_PHN835_U_dsdc_term_cnt_nxt_4_;
   wire FE_PHN834_U_dsdc_term_cnt_nxt_3_;
   wire FE_PHN833_U_dsdc_term_cnt_nxt_2_;
   wire FE_PHN832_cr_reg_data_out_9_;
   wire FE_PHN831_cr_reg_data_out_6_;
   wire FE_PHN816_U_dsdc_n359;
   wire FE_PHN814_U_dsdc_n228;
   wire FE_PHN807_U_cr_N420;
   wire FE_PHN800_U_cr_n96;
   wire FE_PHN799_U_dsdc_n225;
   wire FE_PHN797_U_dsdc_num_init_ref_cnt_nxt_1_;
   wire FE_PHN796_U_dsdc_N4174;
   wire FE_PHN792_U_dsdc_n219;
   wire FE_PHN791_U_dsdc_n1491;
   wire FE_PHN790_U_dsdc_n289;
   wire FE_PHN788_U_dsdc_n554;
   wire FE_PHN787_n90;
   wire FE_PHN786_U_dsdc_n291;
   wire FE_PHN781_U_dsdc_n224;
   wire FE_PHN777_U_dmc_N23;
   wire FE_PHN773_U_dsdc_n1823;
   wire FE_PHN772_U_dsdc_n2095;
   wire FE_PHN771_U_dsdc_n1540;
   wire FE_PHN767_U_dsdc_term_cnt_nxt_1_;
   wire FE_PHN764_U_dsdc_n210;
   wire FE_PHN759_U_cr_N565;
   wire FE_PHN758_U_dsdc_n2096;
   wire FE_PHN757_U_dsdc_auto_ref_en_nxt;
   wire FE_PHN751_U_dsdc_rcar_cnt2_nxt_2_;
   wire FE_PHN745_U_dsdc_n229;
   wire FE_PHN742_U_dsdc_wtr_cnt_nxt_2_;
   wire FE_PHN740_U_dsdc_term_cnt_nxt_0_;
   wire FE_PHN726_n7;
   wire FE_PHN725_cr_reg_data_out_10_;
   wire FE_PHN713_U_dmc_N24;
   wire FE_PHN710_cr_reg_data_out_3_;
   wire FE_PHN706_U_dsdc_n290;
   wire FE_PHN698_U_cr_N414;
   wire FE_PHN697_U_dsdc_n288;
   wire FE_PHN696_U_dsdc_n286;
   wire FE_PHN694_cr_reg_data_out_15_;
   wire FE_PHN691_n5;
   wire FE_PHN683_U_dsdc_n1394;
   wire FE_PHN678_U_dsdc_n896;
   wire FE_PHN672_U_dsdc_n1436;
   wire FE_PHN671_U_dsdc_n1637;
   wire FE_OFN371_cr_t_ras_min_3_;
   wire FE_OFN365_n95;
   wire FE_OFN360_U_addrdec_n26;
   wire FE_OFN357_U_addrdec_n40;
   wire FE_OFN353_U_addrdec_n272;
   wire FE_OFN348_U_cr_n169;
   wire FE_OFN347_U_cr_n290;
   wire FE_OFN345_U_cr_n291;
   wire FE_OFN336_U_cr_n527;
   wire FE_OFN333_U_cr_n528;
   wire FE_OFN332_U_cr_n529;
   wire FE_OFN326_U_cr_n531;
   wire FE_OFN319_U_cr_n548;
   wire FE_OFN316_U_dsdc_n310;
   wire FE_OFN314_U_dsdc_n313;
   wire FE_OFN311_U_dsdc_n620;
   wire FE_OFN304_U_dsdc_n2014;
   wire FE_OFN303_U_dsdc_n2038;
   wire FE_OFN227_hiu_data_25_;
   wire FE_OFN226_hiu_data_26_;
   wire FE_OFN224_hiu_data_29_;
   wire FE_OFN223_hiu_data_30_;
   wire FE_OFN221_hiu_burst_size_0_;
   wire FE_OFN218_hiu_burst_size_2_;
   wire FE_OFN215_hiu_burst_size_4_;
   wire FE_OFN211_debug_ad_col_addr_13_;
   wire FE_OFN189_HRESETn;
   wire FE_OFN188_HRESETn;
   wire FE_OFN187_HRESETn;
   wire FE_OFN186_HRESETn;
   wire FE_OFN183_HRESETn;
   wire FE_OFN173_HRESETn;
   wire FE_OFN172_HRESETn;
   wire FE_OFN148_HRESETn;
   wire FE_OFN142_HRESETn;
   wire FE_OFN141_HRESETn;
   wire FE_OFN64_HRESETn;
   wire FE_OFN63_HRESETn;
   wire FE_OFN59_HRESETn;
   wire FE_OFN50_HRESETn;
   wire FE_OFN45_HRESETn;
   wire FE_OFN44_HRESETn;
   wire FE_OFN39_HRESETn;
   wire FE_OFN36_HRESETn;
   wire FE_OFN25_ctl_push_n;
   wire FE_OFN23_U_cr_n64;
   wire FE_OFN1_U_cr_n541;
   wire FE_OFN0_U_cr_n314;
   wire n27;
   wire n44;
   wire debug_ad_col_addr_13_;
   wire debug_ad_col_addr_12_;
   wire ad_static_mem_req;
   wire cr_do_self_ref_rp;
   wire ctl_burst_done;
   wire ctl_pop_n;
   wire cr_pop_n;
   wire dmc_pop_n;
   wire ctl_push_n;
   wire cr_push_reg_n;
   wire dmc_push_n;
   wire sdram_req_i;
   wire ctl_auto_ref_en;
   wire ctl_ext_mode_reg_done;
   wire ctl_ref_ack;
   wire cr_push_n;
   wire ad_sdram_type_0_;
   wire ad_sdram_chip_select_0_;
   wire cr_s_ready_valid;
   wire cr_do_initialize;
   wire cr_do_power_down;
   wire cr_mode_reg_update;
   wire cr_exn_mode_reg_update;
   wire cr_delayed_precharge;
   wire cr_ref_all_before_sr;
   wire cr_ref_all_after_sr;
   wire ctl_init_done;
   wire ctl_mode_reg_done;
   wire ctl_sd_in_sf_mode;
   wire cr_s_data_width_early_0_;
   wire N28;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n14;
   wire n19;
   wire n21;
   wire U_dsdc_n2085;
   wire U_dsdc_n2084;
   wire U_dsdc_n2083;
   wire U_dsdc_n2082;
   wire U_dsdc_n2081;
   wire U_dsdc_n2080;
   wire U_dsdc_n2079;
   wire U_dsdc_n2078;
   wire U_dsdc_n2077;
   wire U_dsdc_n2076;
   wire U_dsdc_n2075;
   wire U_dsdc_n2074;
   wire U_dsdc_n2073;
   wire U_dsdc_n2072;
   wire U_dsdc_n2071;
   wire U_dsdc_n2070;
   wire U_dsdc_n2069;
   wire U_dsdc_n2068;
   wire U_dsdc_n2067;
   wire U_dsdc_n2066;
   wire U_dsdc_n2065;
   wire U_dsdc_n2064;
   wire U_dsdc_n2063;
   wire U_dsdc_n2062;
   wire U_dsdc_n2061;
   wire U_dsdc_n2060;
   wire U_dsdc_n2059;
   wire U_dsdc_n2058;
   wire U_dsdc_n2057;
   wire U_dsdc_n2056;
   wire U_dsdc_n2055;
   wire U_dsdc_n2052;
   wire U_dsdc_n2051;
   wire U_dsdc_n2050;
   wire U_dsdc_n2049;
   wire U_dsdc_n2048;
   wire U_dsdc_n2047;
   wire U_dsdc_n2046;
   wire U_dsdc_n2045;
   wire U_dsdc_n2044;
   wire U_dsdc_n2043;
   wire U_dsdc_n2042;
   wire U_dsdc_n2041;
   wire U_dsdc_n2040;
   wire U_dsdc_n2039;
   wire U_dsdc_n2038;
   wire U_dsdc_n2037;
   wire U_dsdc_n2036;
   wire U_dsdc_n2035;
   wire U_dsdc_n2034;
   wire U_dsdc_n2033;
   wire U_dsdc_n2032;
   wire U_dsdc_n2031;
   wire U_dsdc_n2030;
   wire U_dsdc_n2029;
   wire U_dsdc_n2028;
   wire U_dsdc_n2027;
   wire U_dsdc_n2026;
   wire U_dsdc_n2025;
   wire U_dsdc_n2024;
   wire U_dsdc_n2023;
   wire U_dsdc_n2014;
   wire U_dsdc_n2013;
   wire U_dsdc_n2012;
   wire U_dsdc_n2007;
   wire U_dsdc_n1991;
   wire U_dsdc_n1980;
   wire U_dsdc_n1979;
   wire U_dsdc_n1978;
   wire U_dsdc_n1977;
   wire U_dsdc_n1976;
   wire U_dsdc_n1975;
   wire U_dsdc_n1974;
   wire U_dsdc_n1973;
   wire U_dsdc_n1972;
   wire U_dsdc_n1971;
   wire U_dsdc_n1970;
   wire U_dsdc_n1969;
   wire U_dsdc_n1968;
   wire U_dsdc_n1967;
   wire U_dsdc_n1966;
   wire U_dsdc_n1965;
   wire U_dsdc_n1964;
   wire U_dsdc_n1963;
   wire U_dsdc_n1962;
   wire U_dsdc_n1961;
   wire U_dsdc_n1960;
   wire U_dsdc_n1959;
   wire U_dsdc_n1958;
   wire U_dsdc_n1957;
   wire U_dsdc_n1956;
   wire U_dsdc_n1954;
   wire U_dsdc_n1953;
   wire U_dsdc_n1951;
   wire U_dsdc_n1948;
   wire U_dsdc_n1947;
   wire U_dsdc_n1946;
   wire U_dsdc_n1945;
   wire U_dsdc_n1944;
   wire U_dsdc_n1943;
   wire U_dsdc_n1942;
   wire U_dsdc_n1941;
   wire U_dsdc_n1940;
   wire U_dsdc_n1939;
   wire U_dsdc_n1938;
   wire U_dsdc_n1937;
   wire U_dsdc_n1936;
   wire U_dsdc_n1935;
   wire U_dsdc_n1934;
   wire U_dsdc_n1933;
   wire U_dsdc_n1932;
   wire U_dsdc_n1931;
   wire U_dsdc_n1930;
   wire U_dsdc_n1929;
   wire U_dsdc_n1928;
   wire U_dsdc_n1927;
   wire U_dsdc_n1926;
   wire U_dsdc_n1925;
   wire U_dsdc_n1924;
   wire U_dsdc_n1923;
   wire U_dsdc_n1922;
   wire U_dsdc_n1921;
   wire U_dsdc_n1920;
   wire U_dsdc_n1919;
   wire U_dsdc_n1918;
   wire U_dsdc_n1917;
   wire U_dsdc_n1916;
   wire U_dsdc_n1915;
   wire U_dsdc_n1914;
   wire U_dsdc_n1913;
   wire U_dsdc_n1912;
   wire U_dsdc_n1911;
   wire U_dsdc_n1910;
   wire U_dsdc_n1909;
   wire U_dsdc_n1908;
   wire U_dsdc_n1907;
   wire U_dsdc_n1906;
   wire U_dsdc_n1905;
   wire U_dsdc_n1904;
   wire U_dsdc_n1903;
   wire U_dsdc_n1902;
   wire U_dsdc_n1901;
   wire U_dsdc_n1900;
   wire U_dsdc_n1899;
   wire U_dsdc_n1898;
   wire U_dsdc_n1897;
   wire U_dsdc_n1896;
   wire U_dsdc_n1895;
   wire U_dsdc_n1894;
   wire U_dsdc_n1893;
   wire U_dsdc_n1892;
   wire U_dsdc_n1891;
   wire U_dsdc_n1890;
   wire U_dsdc_n1889;
   wire U_dsdc_n1888;
   wire U_dsdc_n1887;
   wire U_dsdc_n1886;
   wire U_dsdc_n1885;
   wire U_dsdc_n1884;
   wire U_dsdc_n1883;
   wire U_dsdc_n1882;
   wire U_dsdc_n1881;
   wire U_dsdc_n1880;
   wire U_dsdc_n1879;
   wire U_dsdc_n1878;
   wire U_dsdc_n1877;
   wire U_dsdc_n1876;
   wire U_dsdc_n1875;
   wire U_dsdc_n1874;
   wire U_dsdc_n1872;
   wire U_dsdc_n1871;
   wire U_dsdc_n1870;
   wire U_dsdc_n1869;
   wire U_dsdc_n1868;
   wire U_dsdc_n1867;
   wire U_dsdc_n1866;
   wire U_dsdc_n1865;
   wire U_dsdc_n1864;
   wire U_dsdc_n1863;
   wire U_dsdc_n1862;
   wire U_dsdc_n1861;
   wire U_dsdc_n1860;
   wire U_dsdc_n1859;
   wire U_dsdc_n1858;
   wire U_dsdc_n1857;
   wire U_dsdc_n1856;
   wire U_dsdc_n1855;
   wire U_dsdc_n1854;
   wire U_dsdc_n1853;
   wire U_dsdc_n1852;
   wire U_dsdc_n1851;
   wire U_dsdc_n1850;
   wire U_dsdc_n1849;
   wire U_dsdc_n1848;
   wire U_dsdc_n1847;
   wire U_dsdc_n1846;
   wire U_dsdc_n1844;
   wire U_dsdc_n1843;
   wire U_dsdc_n1842;
   wire U_dsdc_n1841;
   wire U_dsdc_n1840;
   wire U_dsdc_n1839;
   wire U_dsdc_n1837;
   wire U_dsdc_n1836;
   wire U_dsdc_n1834;
   wire U_dsdc_n1833;
   wire U_dsdc_n1832;
   wire U_dsdc_n1831;
   wire U_dsdc_n1830;
   wire U_dsdc_n1829;
   wire U_dsdc_n1828;
   wire U_dsdc_n1827;
   wire U_dsdc_n1826;
   wire U_dsdc_n1825;
   wire U_dsdc_n1824;
   wire U_dsdc_n1823;
   wire U_dsdc_n1822;
   wire U_dsdc_n1821;
   wire U_dsdc_n1820;
   wire U_dsdc_n1817;
   wire U_dsdc_n1815;
   wire U_dsdc_n1813;
   wire U_dsdc_n1812;
   wire U_dsdc_n1805;
   wire U_dsdc_n1804;
   wire U_dsdc_n1803;
   wire U_dsdc_n1802;
   wire U_dsdc_n1801;
   wire U_dsdc_n1800;
   wire U_dsdc_n1799;
   wire U_dsdc_n1798;
   wire U_dsdc_n1797;
   wire U_dsdc_n1796;
   wire U_dsdc_n1795;
   wire U_dsdc_n1794;
   wire U_dsdc_n1793;
   wire U_dsdc_n1792;
   wire U_dsdc_n1791;
   wire U_dsdc_n1790;
   wire U_dsdc_n1789;
   wire U_dsdc_n1788;
   wire U_dsdc_n1787;
   wire U_dsdc_n1786;
   wire U_dsdc_n1785;
   wire U_dsdc_n1784;
   wire U_dsdc_n1783;
   wire U_dsdc_n1782;
   wire U_dsdc_n1781;
   wire U_dsdc_n1780;
   wire U_dsdc_n1779;
   wire U_dsdc_n1778;
   wire U_dsdc_n1777;
   wire U_dsdc_n1776;
   wire U_dsdc_n1775;
   wire U_dsdc_n1774;
   wire U_dsdc_n1773;
   wire U_dsdc_n1772;
   wire U_dsdc_n1771;
   wire U_dsdc_n1770;
   wire U_dsdc_n1769;
   wire U_dsdc_n1768;
   wire U_dsdc_n1767;
   wire U_dsdc_n1766;
   wire U_dsdc_n1765;
   wire U_dsdc_n1764;
   wire U_dsdc_n1763;
   wire U_dsdc_n1762;
   wire U_dsdc_n1761;
   wire U_dsdc_n1760;
   wire U_dsdc_n1759;
   wire U_dsdc_n1758;
   wire U_dsdc_n1757;
   wire U_dsdc_n1756;
   wire U_dsdc_n1755;
   wire U_dsdc_n1754;
   wire U_dsdc_n1753;
   wire U_dsdc_n1752;
   wire U_dsdc_n1751;
   wire U_dsdc_n1750;
   wire U_dsdc_n1749;
   wire U_dsdc_n1748;
   wire U_dsdc_n1747;
   wire U_dsdc_n1746;
   wire U_dsdc_n1745;
   wire U_dsdc_n1744;
   wire U_dsdc_n1743;
   wire U_dsdc_n1742;
   wire U_dsdc_n1741;
   wire U_dsdc_n1740;
   wire U_dsdc_n1739;
   wire U_dsdc_n1738;
   wire U_dsdc_n1737;
   wire U_dsdc_n1736;
   wire U_dsdc_n1735;
   wire U_dsdc_n1734;
   wire U_dsdc_n1733;
   wire U_dsdc_n1732;
   wire U_dsdc_n1731;
   wire U_dsdc_n1730;
   wire U_dsdc_n1729;
   wire U_dsdc_n1728;
   wire U_dsdc_n1727;
   wire U_dsdc_n1726;
   wire U_dsdc_n1725;
   wire U_dsdc_n1724;
   wire U_dsdc_n1723;
   wire U_dsdc_n1722;
   wire U_dsdc_n1721;
   wire U_dsdc_n1720;
   wire U_dsdc_n1719;
   wire U_dsdc_n1718;
   wire U_dsdc_n1717;
   wire U_dsdc_n1716;
   wire U_dsdc_n1715;
   wire U_dsdc_n1714;
   wire U_dsdc_n1713;
   wire U_dsdc_n1712;
   wire U_dsdc_n1711;
   wire U_dsdc_n1710;
   wire U_dsdc_n1709;
   wire U_dsdc_n1708;
   wire U_dsdc_n1707;
   wire U_dsdc_n1706;
   wire U_dsdc_n1705;
   wire U_dsdc_n1704;
   wire U_dsdc_n1703;
   wire U_dsdc_n1702;
   wire U_dsdc_n1701;
   wire U_dsdc_n1700;
   wire U_dsdc_n1699;
   wire U_dsdc_n1698;
   wire U_dsdc_n1697;
   wire U_dsdc_n1696;
   wire U_dsdc_n1695;
   wire U_dsdc_n1694;
   wire U_dsdc_n1693;
   wire U_dsdc_n1692;
   wire U_dsdc_n1691;
   wire U_dsdc_n1690;
   wire U_dsdc_n1689;
   wire U_dsdc_n1688;
   wire U_dsdc_n1687;
   wire U_dsdc_n1686;
   wire U_dsdc_n1685;
   wire U_dsdc_n1684;
   wire U_dsdc_n1683;
   wire U_dsdc_n1682;
   wire U_dsdc_n1681;
   wire U_dsdc_n1680;
   wire U_dsdc_n1679;
   wire U_dsdc_n1678;
   wire U_dsdc_n1677;
   wire U_dsdc_n1676;
   wire U_dsdc_n1675;
   wire U_dsdc_n1674;
   wire U_dsdc_n1673;
   wire U_dsdc_n1672;
   wire U_dsdc_n1671;
   wire U_dsdc_n1670;
   wire U_dsdc_n1669;
   wire U_dsdc_n1668;
   wire U_dsdc_n1667;
   wire U_dsdc_n1666;
   wire U_dsdc_n1662;
   wire U_dsdc_n1661;
   wire U_dsdc_n1660;
   wire U_dsdc_n1659;
   wire U_dsdc_n1658;
   wire U_dsdc_n1657;
   wire U_dsdc_n1656;
   wire U_dsdc_n1655;
   wire U_dsdc_n1654;
   wire U_dsdc_n1653;
   wire U_dsdc_n1652;
   wire U_dsdc_n1651;
   wire U_dsdc_n1650;
   wire U_dsdc_n1649;
   wire U_dsdc_n1648;
   wire U_dsdc_n1647;
   wire U_dsdc_n1646;
   wire U_dsdc_n1645;
   wire U_dsdc_n1644;
   wire U_dsdc_n1643;
   wire U_dsdc_n1642;
   wire U_dsdc_n1641;
   wire U_dsdc_n1640;
   wire U_dsdc_n1639;
   wire U_dsdc_n1638;
   wire U_dsdc_n1637;
   wire U_dsdc_n1636;
   wire U_dsdc_n1635;
   wire U_dsdc_n1634;
   wire U_dsdc_n1633;
   wire U_dsdc_n1632;
   wire U_dsdc_n1631;
   wire U_dsdc_n1630;
   wire U_dsdc_n1629;
   wire U_dsdc_n1628;
   wire U_dsdc_n1627;
   wire U_dsdc_n1625;
   wire U_dsdc_n1624;
   wire U_dsdc_n1623;
   wire U_dsdc_n1622;
   wire U_dsdc_n1621;
   wire U_dsdc_n1620;
   wire U_dsdc_n1619;
   wire U_dsdc_n1618;
   wire U_dsdc_n1617;
   wire U_dsdc_n1616;
   wire U_dsdc_n1615;
   wire U_dsdc_n1614;
   wire U_dsdc_n1612;
   wire U_dsdc_n1611;
   wire U_dsdc_n1610;
   wire U_dsdc_n1609;
   wire U_dsdc_n1608;
   wire U_dsdc_n1606;
   wire U_dsdc_n1605;
   wire U_dsdc_n1604;
   wire U_dsdc_n1603;
   wire U_dsdc_n1602;
   wire U_dsdc_n1601;
   wire U_dsdc_n1600;
   wire U_dsdc_n1598;
   wire U_dsdc_n1597;
   wire U_dsdc_n1596;
   wire U_dsdc_n1594;
   wire U_dsdc_n1593;
   wire U_dsdc_n1592;
   wire U_dsdc_n1591;
   wire U_dsdc_n1590;
   wire U_dsdc_n1589;
   wire U_dsdc_n1588;
   wire U_dsdc_n1587;
   wire U_dsdc_n1586;
   wire U_dsdc_n1585;
   wire U_dsdc_n1584;
   wire U_dsdc_n1583;
   wire U_dsdc_n1582;
   wire U_dsdc_n1581;
   wire U_dsdc_n1580;
   wire U_dsdc_n1579;
   wire U_dsdc_n1578;
   wire U_dsdc_n1577;
   wire U_dsdc_n1576;
   wire U_dsdc_n1575;
   wire U_dsdc_n1574;
   wire U_dsdc_n1573;
   wire U_dsdc_n1572;
   wire U_dsdc_n1571;
   wire U_dsdc_n1570;
   wire U_dsdc_n1569;
   wire U_dsdc_n1568;
   wire U_dsdc_n1567;
   wire U_dsdc_n1566;
   wire U_dsdc_n1565;
   wire U_dsdc_n1564;
   wire U_dsdc_n1563;
   wire U_dsdc_n1562;
   wire U_dsdc_n1561;
   wire U_dsdc_n1560;
   wire U_dsdc_n1559;
   wire U_dsdc_n1558;
   wire U_dsdc_n1557;
   wire U_dsdc_n1556;
   wire U_dsdc_n1546;
   wire U_dsdc_n1545;
   wire U_dsdc_n1544;
   wire U_dsdc_n1543;
   wire U_dsdc_n1542;
   wire U_dsdc_n1541;
   wire U_dsdc_n1540;
   wire U_dsdc_n1539;
   wire U_dsdc_n1538;
   wire U_dsdc_n1537;
   wire U_dsdc_n1536;
   wire U_dsdc_n1535;
   wire U_dsdc_n1534;
   wire U_dsdc_n1533;
   wire U_dsdc_n1532;
   wire U_dsdc_n1531;
   wire U_dsdc_n1530;
   wire U_dsdc_n1529;
   wire U_dsdc_n1528;
   wire U_dsdc_n1527;
   wire U_dsdc_n1526;
   wire U_dsdc_n1525;
   wire U_dsdc_n1524;
   wire U_dsdc_n1523;
   wire U_dsdc_n1522;
   wire U_dsdc_n1521;
   wire U_dsdc_n1520;
   wire U_dsdc_n1519;
   wire U_dsdc_n1518;
   wire U_dsdc_n1517;
   wire U_dsdc_n1516;
   wire U_dsdc_n1515;
   wire U_dsdc_n1514;
   wire U_dsdc_n1513;
   wire U_dsdc_n1512;
   wire U_dsdc_n1511;
   wire U_dsdc_n1510;
   wire U_dsdc_n1509;
   wire U_dsdc_n1508;
   wire U_dsdc_n1507;
   wire U_dsdc_n1506;
   wire U_dsdc_n1505;
   wire U_dsdc_n1504;
   wire U_dsdc_n1503;
   wire U_dsdc_n1502;
   wire U_dsdc_n1501;
   wire U_dsdc_n1500;
   wire U_dsdc_n1499;
   wire U_dsdc_n1498;
   wire U_dsdc_n1497;
   wire U_dsdc_n1496;
   wire U_dsdc_n1495;
   wire U_dsdc_n1493;
   wire U_dsdc_n1492;
   wire U_dsdc_n1491;
   wire U_dsdc_n1490;
   wire U_dsdc_n1489;
   wire U_dsdc_n1488;
   wire U_dsdc_n1487;
   wire U_dsdc_n1486;
   wire U_dsdc_n1485;
   wire U_dsdc_n1484;
   wire U_dsdc_n1483;
   wire U_dsdc_n1482;
   wire U_dsdc_n1481;
   wire U_dsdc_n1480;
   wire U_dsdc_n1479;
   wire U_dsdc_n1478;
   wire U_dsdc_n1477;
   wire U_dsdc_n1476;
   wire U_dsdc_n1475;
   wire U_dsdc_n1474;
   wire U_dsdc_n1473;
   wire U_dsdc_n1472;
   wire U_dsdc_n1471;
   wire U_dsdc_n1470;
   wire U_dsdc_n1469;
   wire U_dsdc_n1468;
   wire U_dsdc_n1467;
   wire U_dsdc_n1466;
   wire U_dsdc_n1465;
   wire U_dsdc_n1464;
   wire U_dsdc_n1462;
   wire U_dsdc_n1461;
   wire U_dsdc_n1460;
   wire U_dsdc_n1458;
   wire U_dsdc_n1455;
   wire U_dsdc_n1454;
   wire U_dsdc_n1452;
   wire U_dsdc_n1451;
   wire U_dsdc_n1450;
   wire U_dsdc_n1449;
   wire U_dsdc_n1448;
   wire U_dsdc_n1447;
   wire U_dsdc_n1446;
   wire U_dsdc_n1445;
   wire U_dsdc_n1444;
   wire U_dsdc_n1438;
   wire U_dsdc_n1437;
   wire U_dsdc_n1436;
   wire U_dsdc_n1435;
   wire U_dsdc_n1434;
   wire U_dsdc_n1433;
   wire U_dsdc_n1432;
   wire U_dsdc_n1431;
   wire U_dsdc_n1430;
   wire U_dsdc_n1429;
   wire U_dsdc_n1428;
   wire U_dsdc_n1427;
   wire U_dsdc_n1426;
   wire U_dsdc_n1425;
   wire U_dsdc_n1424;
   wire U_dsdc_n1423;
   wire U_dsdc_n1422;
   wire U_dsdc_n1421;
   wire U_dsdc_n1420;
   wire U_dsdc_n1419;
   wire U_dsdc_n1418;
   wire U_dsdc_n1417;
   wire U_dsdc_n1416;
   wire U_dsdc_n1415;
   wire U_dsdc_n1414;
   wire U_dsdc_n1413;
   wire U_dsdc_n1412;
   wire U_dsdc_n1411;
   wire U_dsdc_n1410;
   wire U_dsdc_n1409;
   wire U_dsdc_n1403;
   wire U_dsdc_n1398;
   wire U_dsdc_n1397;
   wire U_dsdc_n1396;
   wire U_dsdc_n1395;
   wire U_dsdc_n1394;
   wire U_dsdc_n1393;
   wire U_dsdc_n1392;
   wire U_dsdc_n1391;
   wire U_dsdc_n1390;
   wire U_dsdc_n1389;
   wire U_dsdc_n1388;
   wire U_dsdc_n1387;
   wire U_dsdc_n1386;
   wire U_dsdc_n1385;
   wire U_dsdc_n1384;
   wire U_dsdc_n1383;
   wire U_dsdc_n1382;
   wire U_dsdc_n1381;
   wire U_dsdc_n1380;
   wire U_dsdc_n1379;
   wire U_dsdc_n1377;
   wire U_dsdc_n1376;
   wire U_dsdc_n1375;
   wire U_dsdc_n1374;
   wire U_dsdc_n1373;
   wire U_dsdc_n1372;
   wire U_dsdc_n1371;
   wire U_dsdc_n1370;
   wire U_dsdc_n1369;
   wire U_dsdc_n1368;
   wire U_dsdc_n1367;
   wire U_dsdc_n1366;
   wire U_dsdc_n1365;
   wire U_dsdc_n1364;
   wire U_dsdc_n1363;
   wire U_dsdc_n1362;
   wire U_dsdc_n1361;
   wire U_dsdc_n1360;
   wire U_dsdc_n1359;
   wire U_dsdc_n1358;
   wire U_dsdc_n1357;
   wire U_dsdc_n1356;
   wire U_dsdc_n1355;
   wire U_dsdc_n1354;
   wire U_dsdc_n1353;
   wire U_dsdc_n1352;
   wire U_dsdc_n1351;
   wire U_dsdc_n1350;
   wire U_dsdc_n1349;
   wire U_dsdc_n1348;
   wire U_dsdc_n1347;
   wire U_dsdc_n1346;
   wire U_dsdc_n1345;
   wire U_dsdc_n1344;
   wire U_dsdc_n1343;
   wire U_dsdc_n1342;
   wire U_dsdc_n1341;
   wire U_dsdc_n1340;
   wire U_dsdc_n1339;
   wire U_dsdc_n1338;
   wire U_dsdc_n1337;
   wire U_dsdc_n1336;
   wire U_dsdc_n1335;
   wire U_dsdc_n1334;
   wire U_dsdc_n1333;
   wire U_dsdc_n1332;
   wire U_dsdc_n1331;
   wire U_dsdc_n1330;
   wire U_dsdc_n1329;
   wire U_dsdc_n1328;
   wire U_dsdc_n1327;
   wire U_dsdc_n1326;
   wire U_dsdc_n1325;
   wire U_dsdc_n1324;
   wire U_dsdc_n1323;
   wire U_dsdc_n1322;
   wire U_dsdc_n1321;
   wire U_dsdc_n1320;
   wire U_dsdc_n1319;
   wire U_dsdc_n1318;
   wire U_dsdc_n1317;
   wire U_dsdc_n1316;
   wire U_dsdc_n1315;
   wire U_dsdc_n1314;
   wire U_dsdc_n1313;
   wire U_dsdc_n1312;
   wire U_dsdc_n1311;
   wire U_dsdc_n1310;
   wire U_dsdc_n1309;
   wire U_dsdc_n1308;
   wire U_dsdc_n1307;
   wire U_dsdc_n1306;
   wire U_dsdc_n1305;
   wire U_dsdc_n1304;
   wire U_dsdc_n1303;
   wire U_dsdc_n1302;
   wire U_dsdc_n1301;
   wire U_dsdc_n1300;
   wire U_dsdc_n1299;
   wire U_dsdc_n1298;
   wire U_dsdc_n1297;
   wire U_dsdc_n1296;
   wire U_dsdc_n1295;
   wire U_dsdc_n1294;
   wire U_dsdc_n1293;
   wire U_dsdc_n1292;
   wire U_dsdc_n1291;
   wire U_dsdc_n1290;
   wire U_dsdc_n1289;
   wire U_dsdc_n1288;
   wire U_dsdc_n1287;
   wire U_dsdc_n1286;
   wire U_dsdc_n1285;
   wire U_dsdc_n1284;
   wire U_dsdc_n1283;
   wire U_dsdc_n1282;
   wire U_dsdc_n1281;
   wire U_dsdc_n1280;
   wire U_dsdc_n1279;
   wire U_dsdc_n1278;
   wire U_dsdc_n1277;
   wire U_dsdc_n1276;
   wire U_dsdc_n1275;
   wire U_dsdc_n1274;
   wire U_dsdc_n1273;
   wire U_dsdc_n1272;
   wire U_dsdc_n1271;
   wire U_dsdc_n1270;
   wire U_dsdc_n1269;
   wire U_dsdc_n1268;
   wire U_dsdc_n1267;
   wire U_dsdc_n1266;
   wire U_dsdc_n1264;
   wire U_dsdc_n1263;
   wire U_dsdc_n1262;
   wire U_dsdc_n1261;
   wire U_dsdc_n1260;
   wire U_dsdc_n1259;
   wire U_dsdc_n1258;
   wire U_dsdc_n1254;
   wire U_dsdc_n1253;
   wire U_dsdc_n1252;
   wire U_dsdc_n1251;
   wire U_dsdc_n1250;
   wire U_dsdc_n1249;
   wire U_dsdc_n1248;
   wire U_dsdc_n1247;
   wire U_dsdc_n1246;
   wire U_dsdc_n1245;
   wire U_dsdc_n1244;
   wire U_dsdc_n1243;
   wire U_dsdc_n1241;
   wire U_dsdc_n1239;
   wire U_dsdc_n1238;
   wire U_dsdc_n1237;
   wire U_dsdc_n1235;
   wire U_dsdc_n1234;
   wire U_dsdc_n1233;
   wire U_dsdc_n1231;
   wire U_dsdc_n1229;
   wire U_dsdc_n1228;
   wire U_dsdc_n1227;
   wire U_dsdc_n1225;
   wire U_dsdc_n1224;
   wire U_dsdc_n1223;
   wire U_dsdc_n1222;
   wire U_dsdc_n1221;
   wire U_dsdc_n1220;
   wire U_dsdc_n1219;
   wire U_dsdc_n1218;
   wire U_dsdc_n1217;
   wire U_dsdc_n1216;
   wire U_dsdc_n1215;
   wire U_dsdc_n1214;
   wire U_dsdc_n1213;
   wire U_dsdc_n1212;
   wire U_dsdc_n1211;
   wire U_dsdc_n1210;
   wire U_dsdc_n1209;
   wire U_dsdc_n1208;
   wire U_dsdc_n1207;
   wire U_dsdc_n1206;
   wire U_dsdc_n1205;
   wire U_dsdc_n1204;
   wire U_dsdc_n1203;
   wire U_dsdc_n1202;
   wire U_dsdc_n1201;
   wire U_dsdc_n1200;
   wire U_dsdc_n1199;
   wire U_dsdc_n1198;
   wire U_dsdc_n1197;
   wire U_dsdc_n1196;
   wire U_dsdc_n1195;
   wire U_dsdc_n1194;
   wire U_dsdc_n1193;
   wire U_dsdc_n1192;
   wire U_dsdc_n1191;
   wire U_dsdc_n1190;
   wire U_dsdc_n1189;
   wire U_dsdc_n1188;
   wire U_dsdc_n1187;
   wire U_dsdc_n1186;
   wire U_dsdc_n1185;
   wire U_dsdc_n1184;
   wire U_dsdc_n1183;
   wire U_dsdc_n1182;
   wire U_dsdc_n1181;
   wire U_dsdc_n1180;
   wire U_dsdc_n1179;
   wire U_dsdc_n1178;
   wire U_dsdc_n1177;
   wire U_dsdc_n1176;
   wire U_dsdc_n1175;
   wire U_dsdc_n1174;
   wire U_dsdc_n1173;
   wire U_dsdc_n1172;
   wire U_dsdc_n1171;
   wire U_dsdc_n1170;
   wire U_dsdc_n1169;
   wire U_dsdc_n1168;
   wire U_dsdc_n1167;
   wire U_dsdc_n1166;
   wire U_dsdc_n1165;
   wire U_dsdc_n1164;
   wire U_dsdc_n1163;
   wire U_dsdc_n1162;
   wire U_dsdc_n1161;
   wire U_dsdc_n1160;
   wire U_dsdc_n1159;
   wire U_dsdc_n1158;
   wire U_dsdc_n1157;
   wire U_dsdc_n1156;
   wire U_dsdc_n1155;
   wire U_dsdc_n1154;
   wire U_dsdc_n1153;
   wire U_dsdc_n1152;
   wire U_dsdc_n1151;
   wire U_dsdc_n1150;
   wire U_dsdc_n1149;
   wire U_dsdc_n1148;
   wire U_dsdc_n1147;
   wire U_dsdc_n1146;
   wire U_dsdc_n1145;
   wire U_dsdc_n1144;
   wire U_dsdc_n1143;
   wire U_dsdc_n1137;
   wire U_dsdc_n1136;
   wire U_dsdc_n1134;
   wire U_dsdc_n1132;
   wire U_dsdc_n1130;
   wire U_dsdc_n1127;
   wire U_dsdc_n1124;
   wire U_dsdc_n1123;
   wire U_dsdc_n1122;
   wire U_dsdc_n1117;
   wire U_dsdc_n1116;
   wire U_dsdc_n1115;
   wire U_dsdc_n1112;
   wire U_dsdc_n1111;
   wire U_dsdc_n1110;
   wire U_dsdc_n1109;
   wire U_dsdc_n1104;
   wire U_dsdc_n1103;
   wire U_dsdc_n1098;
   wire U_dsdc_n1097;
   wire U_dsdc_n1095;
   wire U_dsdc_n1094;
   wire U_dsdc_n1093;
   wire U_dsdc_n1092;
   wire U_dsdc_n1091;
   wire U_dsdc_n1090;
   wire U_dsdc_n1089;
   wire U_dsdc_n1088;
   wire U_dsdc_n1087;
   wire U_dsdc_n1085;
   wire U_dsdc_n1084;
   wire U_dsdc_n1082;
   wire U_dsdc_n1081;
   wire U_dsdc_n1079;
   wire U_dsdc_n1076;
   wire U_dsdc_n1075;
   wire U_dsdc_n1073;
   wire U_dsdc_n1069;
   wire U_dsdc_n1064;
   wire U_dsdc_n1063;
   wire U_dsdc_n1062;
   wire U_dsdc_n1061;
   wire U_dsdc_n1060;
   wire U_dsdc_n1059;
   wire U_dsdc_n1058;
   wire U_dsdc_n1053;
   wire U_dsdc_n1052;
   wire U_dsdc_n1051;
   wire U_dsdc_n1044;
   wire U_dsdc_n1043;
   wire U_dsdc_n1042;
   wire U_dsdc_n1041;
   wire U_dsdc_n1040;
   wire U_dsdc_n1038;
   wire U_dsdc_n1037;
   wire U_dsdc_n1033;
   wire U_dsdc_n1032;
   wire U_dsdc_n1031;
   wire U_dsdc_n1028;
   wire U_dsdc_n1027;
   wire U_dsdc_n1026;
   wire U_dsdc_n1025;
   wire U_dsdc_n1024;
   wire U_dsdc_n1023;
   wire U_dsdc_n1022;
   wire U_dsdc_n1021;
   wire U_dsdc_n1020;
   wire U_dsdc_n1019;
   wire U_dsdc_n1018;
   wire U_dsdc_n1017;
   wire U_dsdc_n1016;
   wire U_dsdc_n1015;
   wire U_dsdc_n1014;
   wire U_dsdc_n1013;
   wire U_dsdc_n1012;
   wire U_dsdc_n1011;
   wire U_dsdc_n1010;
   wire U_dsdc_n1009;
   wire U_dsdc_n1008;
   wire U_dsdc_n1007;
   wire U_dsdc_n1006;
   wire U_dsdc_n1005;
   wire U_dsdc_n1004;
   wire U_dsdc_n1003;
   wire U_dsdc_n1002;
   wire U_dsdc_n1001;
   wire U_dsdc_n1000;
   wire U_dsdc_n999;
   wire U_dsdc_n998;
   wire U_dsdc_n997;
   wire U_dsdc_n996;
   wire U_dsdc_n995;
   wire U_dsdc_n994;
   wire U_dsdc_n993;
   wire U_dsdc_n992;
   wire U_dsdc_n991;
   wire U_dsdc_n990;
   wire U_dsdc_n989;
   wire U_dsdc_n988;
   wire U_dsdc_n987;
   wire U_dsdc_n986;
   wire U_dsdc_n985;
   wire U_dsdc_n984;
   wire U_dsdc_n983;
   wire U_dsdc_n982;
   wire U_dsdc_n981;
   wire U_dsdc_n980;
   wire U_dsdc_n979;
   wire U_dsdc_n978;
   wire U_dsdc_n977;
   wire U_dsdc_n976;
   wire U_dsdc_n975;
   wire U_dsdc_n974;
   wire U_dsdc_n972;
   wire U_dsdc_n967;
   wire U_dsdc_n966;
   wire U_dsdc_n964;
   wire U_dsdc_n963;
   wire U_dsdc_n960;
   wire U_dsdc_n959;
   wire U_dsdc_n958;
   wire U_dsdc_n957;
   wire U_dsdc_n956;
   wire U_dsdc_n945;
   wire U_dsdc_n940;
   wire U_dsdc_n939;
   wire U_dsdc_n937;
   wire U_dsdc_n936;
   wire U_dsdc_n935;
   wire U_dsdc_n934;
   wire U_dsdc_n933;
   wire U_dsdc_n921;
   wire U_dsdc_n915;
   wire U_dsdc_n914;
   wire U_dsdc_n913;
   wire U_dsdc_n910;
   wire U_dsdc_n904;
   wire U_dsdc_n903;
   wire U_dsdc_n901;
   wire U_dsdc_n900;
   wire U_dsdc_n899;
   wire U_dsdc_n896;
   wire U_dsdc_n894;
   wire U_dsdc_n893;
   wire U_dsdc_n892;
   wire U_dsdc_n891;
   wire U_dsdc_n890;
   wire U_dsdc_n889;
   wire U_dsdc_n887;
   wire U_dsdc_n886;
   wire U_dsdc_n885;
   wire U_dsdc_n884;
   wire U_dsdc_n883;
   wire U_dsdc_n881;
   wire U_dsdc_n880;
   wire U_dsdc_n879;
   wire U_dsdc_n871;
   wire U_dsdc_n869;
   wire U_dsdc_n868;
   wire U_dsdc_n867;
   wire U_dsdc_n866;
   wire U_dsdc_n865;
   wire U_dsdc_n864;
   wire U_dsdc_n856;
   wire U_dsdc_n852;
   wire U_dsdc_n848;
   wire U_dsdc_n847;
   wire U_dsdc_n846;
   wire U_dsdc_n845;
   wire U_dsdc_n844;
   wire U_dsdc_n843;
   wire U_dsdc_n842;
   wire U_dsdc_n841;
   wire U_dsdc_n840;
   wire U_dsdc_n839;
   wire U_dsdc_n838;
   wire U_dsdc_n837;
   wire U_dsdc_n836;
   wire U_dsdc_n835;
   wire U_dsdc_n834;
   wire U_dsdc_n833;
   wire U_dsdc_n832;
   wire U_dsdc_n831;
   wire U_dsdc_n830;
   wire U_dsdc_n829;
   wire U_dsdc_n828;
   wire U_dsdc_n827;
   wire U_dsdc_n826;
   wire U_dsdc_n825;
   wire U_dsdc_n821;
   wire U_dsdc_n819;
   wire U_dsdc_n818;
   wire U_dsdc_n817;
   wire U_dsdc_n816;
   wire U_dsdc_n815;
   wire U_dsdc_n814;
   wire U_dsdc_n813;
   wire U_dsdc_n812;
   wire U_dsdc_n810;
   wire U_dsdc_n809;
   wire U_dsdc_n808;
   wire U_dsdc_n807;
   wire U_dsdc_n806;
   wire U_dsdc_n805;
   wire U_dsdc_n804;
   wire U_dsdc_n803;
   wire U_dsdc_n802;
   wire U_dsdc_n801;
   wire U_dsdc_n800;
   wire U_dsdc_n799;
   wire U_dsdc_n798;
   wire U_dsdc_n797;
   wire U_dsdc_n796;
   wire U_dsdc_n795;
   wire U_dsdc_n794;
   wire U_dsdc_n793;
   wire U_dsdc_n792;
   wire U_dsdc_n791;
   wire U_dsdc_n790;
   wire U_dsdc_n789;
   wire U_dsdc_n788;
   wire U_dsdc_n787;
   wire U_dsdc_n786;
   wire U_dsdc_n785;
   wire U_dsdc_n784;
   wire U_dsdc_n783;
   wire U_dsdc_n782;
   wire U_dsdc_n778;
   wire U_dsdc_n777;
   wire U_dsdc_n776;
   wire U_dsdc_n775;
   wire U_dsdc_n774;
   wire U_dsdc_n773;
   wire U_dsdc_n772;
   wire U_dsdc_n770;
   wire U_dsdc_n767;
   wire U_dsdc_n766;
   wire U_dsdc_n765;
   wire U_dsdc_n764;
   wire U_dsdc_n763;
   wire U_dsdc_n762;
   wire U_dsdc_n761;
   wire U_dsdc_n760;
   wire U_dsdc_n759;
   wire U_dsdc_n758;
   wire U_dsdc_n757;
   wire U_dsdc_n756;
   wire U_dsdc_n755;
   wire U_dsdc_n754;
   wire U_dsdc_n753;
   wire U_dsdc_n752;
   wire U_dsdc_n751;
   wire U_dsdc_n750;
   wire U_dsdc_n749;
   wire U_dsdc_n748;
   wire U_dsdc_n747;
   wire U_dsdc_n746;
   wire U_dsdc_n745;
   wire U_dsdc_n744;
   wire U_dsdc_n741;
   wire U_dsdc_n740;
   wire U_dsdc_n739;
   wire U_dsdc_n738;
   wire U_dsdc_n737;
   wire U_dsdc_n736;
   wire U_dsdc_n735;
   wire U_dsdc_n734;
   wire U_dsdc_n733;
   wire U_dsdc_n732;
   wire U_dsdc_n731;
   wire U_dsdc_n730;
   wire U_dsdc_n729;
   wire U_dsdc_n728;
   wire U_dsdc_n727;
   wire U_dsdc_n726;
   wire U_dsdc_n725;
   wire U_dsdc_n724;
   wire U_dsdc_n723;
   wire U_dsdc_n722;
   wire U_dsdc_n721;
   wire U_dsdc_n720;
   wire U_dsdc_n718;
   wire U_dsdc_n717;
   wire U_dsdc_n716;
   wire U_dsdc_n715;
   wire U_dsdc_n714;
   wire U_dsdc_n713;
   wire U_dsdc_n712;
   wire U_dsdc_n711;
   wire U_dsdc_n710;
   wire U_dsdc_n708;
   wire U_dsdc_n705;
   wire U_dsdc_n704;
   wire U_dsdc_n703;
   wire U_dsdc_n693;
   wire U_dsdc_n692;
   wire U_dsdc_n691;
   wire U_dsdc_n690;
   wire U_dsdc_n689;
   wire U_dsdc_n688;
   wire U_dsdc_n687;
   wire U_dsdc_n686;
   wire U_dsdc_n685;
   wire U_dsdc_n684;
   wire U_dsdc_n683;
   wire U_dsdc_n682;
   wire U_dsdc_n676;
   wire U_dsdc_n675;
   wire U_dsdc_n674;
   wire U_dsdc_n673;
   wire U_dsdc_n672;
   wire U_dsdc_n670;
   wire U_dsdc_n669;
   wire U_dsdc_n668;
   wire U_dsdc_n667;
   wire U_dsdc_n666;
   wire U_dsdc_n663;
   wire U_dsdc_n662;
   wire U_dsdc_n661;
   wire U_dsdc_n660;
   wire U_dsdc_n659;
   wire U_dsdc_n658;
   wire U_dsdc_n657;
   wire U_dsdc_n654;
   wire U_dsdc_n653;
   wire U_dsdc_n652;
   wire U_dsdc_n651;
   wire U_dsdc_n650;
   wire U_dsdc_n649;
   wire U_dsdc_n648;
   wire U_dsdc_n646;
   wire U_dsdc_n645;
   wire U_dsdc_n644;
   wire U_dsdc_n643;
   wire U_dsdc_n642;
   wire U_dsdc_n641;
   wire U_dsdc_n621;
   wire U_dsdc_n620;
   wire U_dsdc_n619;
   wire U_dsdc_n618;
   wire U_dsdc_n617;
   wire U_dsdc_n616;
   wire U_dsdc_n615;
   wire U_dsdc_n614;
   wire U_dsdc_n613;
   wire U_dsdc_n612;
   wire U_dsdc_n611;
   wire U_dsdc_n610;
   wire U_dsdc_n609;
   wire U_dsdc_n608;
   wire U_dsdc_n607;
   wire U_dsdc_n606;
   wire U_dsdc_n604;
   wire U_dsdc_n603;
   wire U_dsdc_n602;
   wire U_dsdc_n601;
   wire U_dsdc_n600;
   wire U_dsdc_n599;
   wire U_dsdc_n598;
   wire U_dsdc_n597;
   wire U_dsdc_n596;
   wire U_dsdc_n595;
   wire U_dsdc_n594;
   wire U_dsdc_n593;
   wire U_dsdc_n592;
   wire U_dsdc_n591;
   wire U_dsdc_n590;
   wire U_dsdc_n589;
   wire U_dsdc_n588;
   wire U_dsdc_n587;
   wire U_dsdc_n586;
   wire U_dsdc_n585;
   wire U_dsdc_n584;
   wire U_dsdc_n583;
   wire U_dsdc_n582;
   wire U_dsdc_n581;
   wire U_dsdc_n580;
   wire U_dsdc_n579;
   wire U_dsdc_n578;
   wire U_dsdc_n577;
   wire U_dsdc_n576;
   wire U_dsdc_n575;
   wire U_dsdc_n574;
   wire U_dsdc_n573;
   wire U_dsdc_n572;
   wire U_dsdc_n571;
   wire U_dsdc_n570;
   wire U_dsdc_n569;
   wire U_dsdc_n568;
   wire U_dsdc_n567;
   wire U_dsdc_n566;
   wire U_dsdc_n565;
   wire U_dsdc_n564;
   wire U_dsdc_n563;
   wire U_dsdc_n562;
   wire U_dsdc_n561;
   wire U_dsdc_n560;
   wire U_dsdc_n559;
   wire U_dsdc_n558;
   wire U_dsdc_n557;
   wire U_dsdc_n556;
   wire U_dsdc_n555;
   wire U_dsdc_n553;
   wire U_dsdc_n552;
   wire U_dsdc_n551;
   wire U_dsdc_n550;
   wire U_dsdc_n549;
   wire U_dsdc_n548;
   wire U_dsdc_n547;
   wire U_dsdc_n546;
   wire U_dsdc_n545;
   wire U_dsdc_n544;
   wire U_dsdc_n543;
   wire U_dsdc_n542;
   wire U_dsdc_n541;
   wire U_dsdc_n540;
   wire U_dsdc_n539;
   wire U_dsdc_n538;
   wire U_dsdc_n537;
   wire U_dsdc_n536;
   wire U_dsdc_n535;
   wire U_dsdc_n534;
   wire U_dsdc_n533;
   wire U_dsdc_n532;
   wire U_dsdc_n531;
   wire U_dsdc_n530;
   wire U_dsdc_n529;
   wire U_dsdc_n528;
   wire U_dsdc_n527;
   wire U_dsdc_n526;
   wire U_dsdc_n525;
   wire U_dsdc_n524;
   wire U_dsdc_n523;
   wire U_dsdc_n522;
   wire U_dsdc_n519;
   wire U_dsdc_n517;
   wire U_dsdc_n516;
   wire U_dsdc_n515;
   wire U_dsdc_n514;
   wire U_dsdc_n513;
   wire U_dsdc_n512;
   wire U_dsdc_n511;
   wire U_dsdc_n510;
   wire U_dsdc_n509;
   wire U_dsdc_n508;
   wire U_dsdc_n507;
   wire U_dsdc_n504;
   wire U_dsdc_n503;
   wire U_dsdc_n502;
   wire U_dsdc_n501;
   wire U_dsdc_n500;
   wire U_dsdc_n499;
   wire U_dsdc_n498;
   wire U_dsdc_n497;
   wire U_dsdc_n496;
   wire U_dsdc_n495;
   wire U_dsdc_n494;
   wire U_dsdc_n493;
   wire U_dsdc_n492;
   wire U_dsdc_n491;
   wire U_dsdc_n488;
   wire U_dsdc_n487;
   wire U_dsdc_n486;
   wire U_dsdc_n485;
   wire U_dsdc_n484;
   wire U_dsdc_n483;
   wire U_dsdc_n482;
   wire U_dsdc_n481;
   wire U_dsdc_n480;
   wire U_dsdc_n479;
   wire U_dsdc_n478;
   wire U_dsdc_n477;
   wire U_dsdc_n476;
   wire U_dsdc_n474;
   wire U_dsdc_n473;
   wire U_dsdc_n468;
   wire U_dsdc_n467;
   wire U_dsdc_n465;
   wire U_dsdc_n464;
   wire U_dsdc_n463;
   wire U_dsdc_n462;
   wire U_dsdc_n461;
   wire U_dsdc_n460;
   wire U_dsdc_n459;
   wire U_dsdc_n458;
   wire U_dsdc_n457;
   wire U_dsdc_n456;
   wire U_dsdc_n455;
   wire U_dsdc_n454;
   wire U_dsdc_n453;
   wire U_dsdc_n452;
   wire U_dsdc_n451;
   wire U_dsdc_n450;
   wire U_dsdc_n449;
   wire U_dsdc_n448;
   wire U_dsdc_n447;
   wire U_dsdc_n442;
   wire U_dsdc_n441;
   wire U_dsdc_n440;
   wire U_dsdc_n439;
   wire U_dsdc_n438;
   wire U_dsdc_n437;
   wire U_dsdc_n436;
   wire U_dsdc_n435;
   wire U_dsdc_n434;
   wire U_dsdc_n433;
   wire U_dsdc_n432;
   wire U_dsdc_n430;
   wire U_dsdc_n429;
   wire U_dsdc_n428;
   wire U_dsdc_n427;
   wire U_dsdc_n426;
   wire U_dsdc_n425;
   wire U_dsdc_n424;
   wire U_dsdc_n422;
   wire U_dsdc_n421;
   wire U_dsdc_n420;
   wire U_dsdc_n419;
   wire U_dsdc_n402;
   wire U_dsdc_n401;
   wire U_dsdc_n400;
   wire U_dsdc_n399;
   wire U_dsdc_n398;
   wire U_dsdc_n397;
   wire U_dsdc_n396;
   wire U_dsdc_n395;
   wire U_dsdc_n385;
   wire U_dsdc_n384;
   wire U_dsdc_n383;
   wire U_dsdc_n382;
   wire U_dsdc_n365;
   wire U_dsdc_n364;
   wire U_dsdc_n363;
   wire U_dsdc_n362;
   wire U_dsdc_n361;
   wire U_dsdc_n360;
   wire U_dsdc_n359;
   wire U_dsdc_n358;
   wire U_dsdc_n357;
   wire U_dsdc_n356;
   wire U_dsdc_n355;
   wire U_dsdc_n354;
   wire U_dsdc_n353;
   wire U_dsdc_n352;
   wire U_dsdc_n351;
   wire U_dsdc_n350;
   wire U_dsdc_n349;
   wire U_dsdc_n347;
   wire U_dsdc_n346;
   wire U_dsdc_n345;
   wire U_dsdc_n344;
   wire U_dsdc_n343;
   wire U_dsdc_n342;
   wire U_dsdc_n341;
   wire U_dsdc_n340;
   wire U_dsdc_n339;
   wire U_dsdc_n338;
   wire U_dsdc_n337;
   wire U_dsdc_n336;
   wire U_dsdc_n335;
   wire U_dsdc_n334;
   wire U_dsdc_n333;
   wire U_dsdc_n332;
   wire U_dsdc_n331;
   wire U_dsdc_n330;
   wire U_dsdc_n328;
   wire U_dsdc_n327;
   wire U_dsdc_n326;
   wire U_dsdc_n325;
   wire U_dsdc_n318;
   wire U_dsdc_n314;
   wire U_dsdc_n312;
   wire U_dsdc_n309;
   wire U_dsdc_n308;
   wire U_dsdc_n306;
   wire U_dsdc_n305;
   wire U_dsdc_n304;
   wire U_dsdc_n303;
   wire U_dsdc_n302;
   wire U_dsdc_n301;
   wire U_dsdc_n299;
   wire U_dsdc_n298;
   wire U_dsdc_n292;
   wire U_dsdc_n284;
   wire U_dsdc_n239;
   wire U_dsdc_n208;
   wire U_dsdc_n207;
   wire U_dsdc_n206;
   wire U_dsdc_n205;
   wire U_dsdc_n204;
   wire U_dsdc_n203;
   wire U_dsdc_n202;
   wire U_dsdc_n201;
   wire U_dsdc_n200;
   wire U_dsdc_n199;
   wire U_dsdc_n198;
   wire U_dsdc_n197;
   wire U_dsdc_n196;
   wire U_dsdc_n195;
   wire U_dsdc_n194;
   wire U_dsdc_n193;
   wire U_dsdc_n192;
   wire U_dsdc_n191;
   wire U_dsdc_n190;
   wire U_dsdc_n189;
   wire U_dsdc_n188;
   wire U_dsdc_n187;
   wire U_dsdc_n186;
   wire U_dsdc_n185;
   wire U_dsdc_n184;
   wire U_dsdc_n183;
   wire U_dsdc_n182;
   wire U_dsdc_n181;
   wire U_dsdc_n180;
   wire U_dsdc_n179;
   wire U_dsdc_n178;
   wire U_dsdc_n177;
   wire U_dsdc_n176;
   wire U_dsdc_n174;
   wire U_dsdc_n173;
   wire U_dsdc_n172;
   wire U_dsdc_n171;
   wire U_dsdc_n170;
   wire U_dsdc_n169;
   wire U_dsdc_n168;
   wire U_dsdc_n167;
   wire U_dsdc_n166;
   wire U_dsdc_n165;
   wire U_dsdc_n164;
   wire U_dsdc_n163;
   wire U_dsdc_n162;
   wire U_dsdc_n159;
   wire U_dsdc_n158;
   wire U_dsdc_n157;
   wire U_dsdc_n156;
   wire U_dsdc_n155;
   wire U_dsdc_n154;
   wire U_dsdc_n153;
   wire U_dsdc_n152;
   wire U_dsdc_n151;
   wire U_dsdc_n150;
   wire U_dsdc_n149;
   wire U_dsdc_n148;
   wire U_dsdc_n147;
   wire U_dsdc_n145;
   wire U_dsdc_n144;
   wire U_dsdc_n143;
   wire U_dsdc_n142;
   wire U_dsdc_n141;
   wire U_dsdc_n140;
   wire U_dsdc_n139;
   wire U_dsdc_n137;
   wire U_dsdc_n134;
   wire U_dsdc_n133;
   wire U_dsdc_n131;
   wire U_dsdc_n130;
   wire U_dsdc_n129;
   wire U_dsdc_n128;
   wire U_dsdc_n126;
   wire U_dsdc_n125;
   wire U_dsdc_n124;
   wire U_dsdc_n123;
   wire U_dsdc_n121;
   wire U_dsdc_n120;
   wire U_dsdc_n109;
   wire U_dsdc_n108;
   wire U_dsdc_n107;
   wire U_dsdc_n106;
   wire U_dsdc_n105;
   wire U_dsdc_n101;
   wire U_dsdc_n100;
   wire U_dsdc_n99;
   wire U_dsdc_n98;
   wire U_dsdc_n92;
   wire U_dsdc_n90;
   wire U_dsdc_n89;
   wire U_dsdc_n88;
   wire U_dsdc_n87;
   wire U_dsdc_n86;
   wire U_dsdc_n84;
   wire U_dsdc_n82;
   wire U_dsdc_n81;
   wire U_dsdc_n80;
   wire U_dsdc_n75;
   wire U_dsdc_n74;
   wire U_dsdc_n73;
   wire U_dsdc_n72;
   wire U_dsdc_n71;
   wire U_dsdc_n70;
   wire U_dsdc_n69;
   wire U_dsdc_n68;
   wire U_dsdc_n67;
   wire U_dsdc_n66;
   wire U_dsdc_n65;
   wire U_dsdc_n63;
   wire U_dsdc_n62;
   wire U_dsdc_n60;
   wire U_dsdc_n59;
   wire U_dsdc_n58;
   wire U_dsdc_n53;
   wire U_dsdc_n52;
   wire U_dsdc_n51;
   wire U_dsdc_n48;
   wire U_dsdc_n47;
   wire U_dsdc_n46;
   wire U_dsdc_n45;
   wire U_dsdc_n44;
   wire U_dsdc_n43;
   wire U_dsdc_n42;
   wire U_dsdc_n41;
   wire U_dsdc_n40;
   wire U_dsdc_n39;
   wire U_dsdc_n36;
   wire U_dsdc_n35;
   wire U_dsdc_n34;
   wire U_dsdc_n33;
   wire U_dsdc_n30;
   wire U_dsdc_n29;
   wire U_dsdc_n28;
   wire U_dsdc_n27;
   wire U_dsdc_n26;
   wire U_dsdc_n25;
   wire U_dsdc_n24;
   wire U_dsdc_n23;
   wire U_dsdc_n22;
   wire U_dsdc_n18;
   wire U_dsdc_n17;
   wire U_dsdc_n16;
   wire U_dsdc_n15;
   wire U_dsdc_n14;
   wire U_dsdc_n12;
   wire U_dsdc_n11;
   wire U_dsdc_n10;
   wire U_dsdc_n9;
   wire U_dsdc_n8;
   wire U_dsdc_n7;
   wire U_dsdc_n6;
   wire U_dsdc_n5;
   wire U_dsdc_n4;
   wire U_dsdc_n3;
   wire U_dsdc_n2;
   wire U_dsdc_n1;
   wire U_dsdc_DP_OP_1642_126_2028_n1;
   wire U_dsdc_DP_OP_1642_126_2028_n2;
   wire U_dsdc_DP_OP_1642_126_2028_n3;
   wire U_dsdc_DP_OP_1642_126_2028_n4;
   wire U_dsdc_DP_OP_1642_126_2028_n5;
   wire U_dsdc_DP_OP_1642_126_2028_n6;
   wire U_dsdc_DP_OP_1642_126_2028_n7;
   wire U_dsdc_DP_OP_1642_126_2028_n8;
   wire U_dsdc_DP_OP_1642_126_2028_n9;
   wire U_dsdc_DP_OP_1642_126_2028_n11;
   wire U_dsdc_DP_OP_1642_126_2028_n12;
   wire U_dsdc_DP_OP_1642_126_2028_n13;
   wire U_dsdc_DP_OP_1642_126_2028_n14;
   wire U_dsdc_DP_OP_1642_126_2028_n15;
   wire U_dsdc_DP_OP_1642_126_2028_n19;
   wire U_dsdc_DP_OP_1642_126_2028_n20;
   wire U_dsdc_DP_OP_1642_126_2028_n21;
   wire U_dsdc_DP_OP_1642_126_2028_n23;
   wire U_dsdc_DP_OP_1642_126_2028_n24;
   wire U_dsdc_DP_OP_1642_126_2028_n25;
   wire U_dsdc_DP_OP_1642_126_2028_n26;
   wire U_dsdc_DP_OP_1642_126_2028_n27;
   wire U_dsdc_DP_OP_1642_126_2028_n28;
   wire U_dsdc_DP_OP_1642_126_2028_n30;
   wire U_dsdc_DP_OP_1642_126_2028_n31;
   wire U_dsdc_DP_OP_1642_126_2028_n34;
   wire U_dsdc_DP_OP_1642_126_2028_n35;
   wire U_dsdc_DP_OP_1642_126_2028_n36;
   wire U_dsdc_DP_OP_1642_126_2028_n37;
   wire U_dsdc_DP_OP_1642_126_2028_n38;
   wire U_dsdc_DP_OP_1642_126_2028_n39;
   wire U_dsdc_DP_OP_1642_126_2028_n40;
   wire U_dsdc_DP_OP_1642_126_2028_n42;
   wire U_dsdc_DP_OP_1642_126_2028_n43;
   wire U_dsdc_DP_OP_1642_126_2028_n44;
   wire U_dsdc_DP_OP_1642_126_2028_n45;
   wire U_dsdc_DP_OP_1642_126_2028_n46;
   wire U_dsdc_DP_OP_1642_126_2028_n47;
   wire U_dsdc_DP_OP_1642_126_2028_n48;
   wire U_dsdc_DP_OP_1642_126_2028_n49;
   wire U_dsdc_DP_OP_1642_126_2028_n50;
   wire U_dsdc_DP_OP_1642_126_2028_n51;
   wire U_dsdc_DP_OP_1642_126_2028_n52;
   wire U_dsdc_DP_OP_1642_126_2028_n58;
   wire U_dsdc_DP_OP_1642_126_2028_n59;
   wire U_dsdc_DP_OP_1642_126_2028_n60;
   wire U_dsdc_DP_OP_1642_126_2028_n61;
   wire U_dsdc_DP_OP_1642_126_2028_n62;
   wire U_dsdc_DP_OP_1642_126_2028_n85;
   wire U_dsdc_DP_OP_1642_126_2028_n86;
   wire U_dsdc_DP_OP_1642_126_2028_I6;
   wire U_dsdc_DP_OP_1642_126_2028_I5_0_;
   wire U_dsdc_DP_OP_1642_126_2028_I5_1_;
   wire U_dsdc_DP_OP_1642_126_2028_I5_2_;
   wire U_dsdc_DP_OP_1642_126_2028_I5_3_;
   wire U_dsdc_DP_OP_1642_126_2028_I5_4_;
   wire U_dsdc_DP_OP_1642_126_2028_I5_5_;
   wire U_dsdc_DP_OP_1642_126_2028_I4;
   wire U_dsdc_RSOP_1683_C2_CONTROL1;
   wire U_dsdc_n554;
   wire U_dsdc_n431;
   wire U_dsdc_n423;
   wire U_dsdc_n418;
   wire U_dsdc_n417;
   wire U_dsdc_n416;
   wire U_dsdc_n415;
   wire U_dsdc_n414;
   wire U_dsdc_n413;
   wire U_dsdc_n412;
   wire U_dsdc_n411;
   wire U_dsdc_n410;
   wire U_dsdc_n409;
   wire U_dsdc_n408;
   wire U_dsdc_n407;
   wire U_dsdc_n406;
   wire U_dsdc_n405;
   wire U_dsdc_n404;
   wire U_dsdc_n403;
   wire U_dsdc_n394;
   wire U_dsdc_n393;
   wire U_dsdc_n392;
   wire U_dsdc_n391;
   wire U_dsdc_n390;
   wire U_dsdc_n389;
   wire U_dsdc_n388;
   wire U_dsdc_n387;
   wire U_dsdc_n386;
   wire U_dsdc_n381;
   wire U_dsdc_n380;
   wire U_dsdc_n379;
   wire U_dsdc_n378;
   wire U_dsdc_n377;
   wire U_dsdc_n376;
   wire U_dsdc_n375;
   wire U_dsdc_n374;
   wire U_dsdc_n373;
   wire U_dsdc_n372;
   wire U_dsdc_n371;
   wire U_dsdc_n370;
   wire U_dsdc_n369;
   wire U_dsdc_n368;
   wire U_dsdc_n367;
   wire U_dsdc_n366;
   wire U_dsdc_n329;
   wire U_dsdc_n319;
   wire U_dsdc_n313;
   wire U_dsdc_n310;
   wire U_dsdc_n307;
   wire U_dsdc_n300;
   wire U_dsdc_n297;
   wire U_dsdc_n296;
   wire U_dsdc_n295;
   wire U_dsdc_n294;
   wire U_dsdc_n293;
   wire U_dsdc_n291;
   wire U_dsdc_n290;
   wire U_dsdc_n289;
   wire U_dsdc_n288;
   wire U_dsdc_n287;
   wire U_dsdc_n286;
   wire U_dsdc_n283;
   wire U_dsdc_n282;
   wire U_dsdc_n281;
   wire U_dsdc_n280;
   wire U_dsdc_n279;
   wire U_dsdc_n277;
   wire U_dsdc_n276;
   wire U_dsdc_n275;
   wire U_dsdc_n274;
   wire U_dsdc_n273;
   wire U_dsdc_n272;
   wire U_dsdc_n271;
   wire U_dsdc_n270;
   wire U_dsdc_n269;
   wire U_dsdc_n268;
   wire U_dsdc_n267;
   wire U_dsdc_n266;
   wire U_dsdc_n265;
   wire U_dsdc_n264;
   wire U_dsdc_n263;
   wire U_dsdc_n262;
   wire U_dsdc_n261;
   wire U_dsdc_n260;
   wire U_dsdc_n259;
   wire U_dsdc_n258;
   wire U_dsdc_n257;
   wire U_dsdc_n256;
   wire U_dsdc_n255;
   wire U_dsdc_n240;
   wire U_dsdc_n231;
   wire U_dsdc_n230;
   wire U_dsdc_n229;
   wire U_dsdc_n228;
   wire U_dsdc_n227;
   wire U_dsdc_n226;
   wire U_dsdc_n225;
   wire U_dsdc_n224;
   wire U_dsdc_n223;
   wire U_dsdc_n222;
   wire U_dsdc_n221;
   wire U_dsdc_n220;
   wire U_dsdc_n219;
   wire U_dsdc_n218;
   wire U_dsdc_n216;
   wire U_dsdc_n215;
   wire U_dsdc_n214;
   wire U_dsdc_n213;
   wire U_dsdc_n212;
   wire U_dsdc_n211;
   wire U_dsdc_n210;
   wire U_dsdc_n209;
   wire U_dsdc_add_x_2600_1_n8;
   wire U_dsdc_C880_DATA5_5;
   wire U_dsdc_C880_DATA5_3;
   wire U_dsdc_C880_DATA5_1;
   wire U_dsdc_bm_bank_age_0__0_;
   wire U_dsdc_bm_bank_age_0__1_;
   wire U_dsdc_bm_bank_age_0__2_;
   wire U_dsdc_bm_bank_age_0__3_;
   wire U_dsdc_bm_bank_age_0__4_;
   wire U_dsdc_bm_bank_age_1__0_;
   wire U_dsdc_bm_bank_age_1__1_;
   wire U_dsdc_bm_bank_age_1__2_;
   wire U_dsdc_bm_bank_age_1__3_;
   wire U_dsdc_bm_bank_age_1__4_;
   wire U_dsdc_bm_bank_age_2__0_;
   wire U_dsdc_bm_bank_age_2__1_;
   wire U_dsdc_bm_bank_age_2__2_;
   wire U_dsdc_bm_bank_age_2__3_;
   wire U_dsdc_bm_bank_age_2__4_;
   wire U_dsdc_bm_bank_age_3__0_;
   wire U_dsdc_bm_bank_age_3__1_;
   wire U_dsdc_bm_bank_age_3__2_;
   wire U_dsdc_bm_bank_age_3__3_;
   wire U_dsdc_bm_bank_age_3__4_;
   wire U_dsdc_N4496;
   wire U_dsdc_N4492;
   wire U_dsdc_N4491;
   wire U_dsdc_N4490;
   wire U_dsdc_N4489;
   wire U_dsdc_N4488;
   wire U_dsdc_N4487;
   wire U_dsdc_N4486;
   wire U_dsdc_N4485;
   wire U_dsdc_N4484;
   wire U_dsdc_N4483;
   wire U_dsdc_N4482;
   wire U_dsdc_N4481;
   wire U_dsdc_N4480;
   wire U_dsdc_N4479;
   wire U_dsdc_N4478;
   wire U_dsdc_N4477;
   wire U_dsdc_N4476;
   wire U_dsdc_N4475;
   wire U_dsdc_N4474;
   wire U_dsdc_N4473;
   wire U_dsdc_N4463;
   wire U_dsdc_N4462;
   wire U_dsdc_N4461;
   wire U_dsdc_N4460;
   wire U_dsdc_N4449;
   wire U_dsdc_N4445;
   wire U_dsdc_N4444;
   wire U_dsdc_N4443;
   wire U_dsdc_N4442;
   wire U_dsdc_N4441;
   wire U_dsdc_N4440;
   wire U_dsdc_N4439;
   wire U_dsdc_N4438;
   wire U_dsdc_N4437;
   wire U_dsdc_N4436;
   wire U_dsdc_N4435;
   wire U_dsdc_N4434;
   wire U_dsdc_N4433;
   wire U_dsdc_N4432;
   wire U_dsdc_N4431;
   wire U_dsdc_N4430;
   wire U_dsdc_N4429;
   wire U_dsdc_N4428;
   wire U_dsdc_N4427;
   wire U_dsdc_N4426;
   wire U_dsdc_N4416;
   wire U_dsdc_N4415;
   wire U_dsdc_N4414;
   wire U_dsdc_N4413;
   wire U_dsdc_N4402;
   wire U_dsdc_N4398;
   wire U_dsdc_N4397;
   wire U_dsdc_N4396;
   wire U_dsdc_N4395;
   wire U_dsdc_N4394;
   wire U_dsdc_N4393;
   wire U_dsdc_N4392;
   wire U_dsdc_N4391;
   wire U_dsdc_N4390;
   wire U_dsdc_N4389;
   wire U_dsdc_N4388;
   wire U_dsdc_N4387;
   wire U_dsdc_N4386;
   wire U_dsdc_N4385;
   wire U_dsdc_N4384;
   wire U_dsdc_N4383;
   wire U_dsdc_N4382;
   wire U_dsdc_N4381;
   wire U_dsdc_N4380;
   wire U_dsdc_N4379;
   wire U_dsdc_N4369;
   wire U_dsdc_N4368;
   wire U_dsdc_N4367;
   wire U_dsdc_N4366;
   wire U_dsdc_N4355;
   wire U_dsdc_N4351;
   wire U_dsdc_N4350;
   wire U_dsdc_N4349;
   wire U_dsdc_N4348;
   wire U_dsdc_N4347;
   wire U_dsdc_N4346;
   wire U_dsdc_N4345;
   wire U_dsdc_N4344;
   wire U_dsdc_N4343;
   wire U_dsdc_N4342;
   wire U_dsdc_N4341;
   wire U_dsdc_N4340;
   wire U_dsdc_N4339;
   wire U_dsdc_N4338;
   wire U_dsdc_N4337;
   wire U_dsdc_N4336;
   wire U_dsdc_N4335;
   wire U_dsdc_N4334;
   wire U_dsdc_N4333;
   wire U_dsdc_N4332;
   wire U_dsdc_N4322;
   wire U_dsdc_N4321;
   wire U_dsdc_N4320;
   wire U_dsdc_N4319;
   wire U_dsdc_N4284;
   wire U_dsdc_N4283;
   wire U_dsdc_N4282;
   wire U_dsdc_N4281;
   wire U_dsdc_bm_ras_cnt_0__0_;
   wire U_dsdc_bm_ras_cnt_0__1_;
   wire U_dsdc_bm_ras_cnt_0__2_;
   wire U_dsdc_bm_ras_cnt_0__3_;
   wire U_dsdc_bm_ras_cnt_1__0_;
   wire U_dsdc_bm_ras_cnt_1__1_;
   wire U_dsdc_bm_ras_cnt_1__2_;
   wire U_dsdc_bm_ras_cnt_1__3_;
   wire U_dsdc_bm_ras_cnt_2__0_;
   wire U_dsdc_bm_ras_cnt_2__1_;
   wire U_dsdc_bm_ras_cnt_2__2_;
   wire U_dsdc_bm_ras_cnt_2__3_;
   wire U_dsdc_bm_ras_cnt_3__0_;
   wire U_dsdc_bm_ras_cnt_3__1_;
   wire U_dsdc_bm_ras_cnt_3__2_;
   wire U_dsdc_bm_ras_cnt_3__3_;
   wire U_dsdc_bm_rc_cnt_0__0_;
   wire U_dsdc_bm_rc_cnt_0__1_;
   wire U_dsdc_bm_rc_cnt_0__2_;
   wire U_dsdc_bm_rc_cnt_0__3_;
   wire U_dsdc_bm_rc_cnt_1__0_;
   wire U_dsdc_bm_rc_cnt_1__1_;
   wire U_dsdc_bm_rc_cnt_1__2_;
   wire U_dsdc_bm_rc_cnt_1__3_;
   wire U_dsdc_bm_rc_cnt_2__0_;
   wire U_dsdc_bm_rc_cnt_2__1_;
   wire U_dsdc_bm_rc_cnt_2__2_;
   wire U_dsdc_bm_rc_cnt_2__3_;
   wire U_dsdc_bm_rc_cnt_3__0_;
   wire U_dsdc_bm_rc_cnt_3__1_;
   wire U_dsdc_bm_rc_cnt_3__2_;
   wire U_dsdc_bm_rc_cnt_3__3_;
   wire U_dsdc_bm_row_addr_0__0_;
   wire U_dsdc_bm_row_addr_0__1_;
   wire U_dsdc_bm_row_addr_0__2_;
   wire U_dsdc_bm_row_addr_0__3_;
   wire U_dsdc_bm_row_addr_0__4_;
   wire U_dsdc_bm_row_addr_0__5_;
   wire U_dsdc_bm_row_addr_0__6_;
   wire U_dsdc_bm_row_addr_0__7_;
   wire U_dsdc_bm_row_addr_0__8_;
   wire U_dsdc_bm_row_addr_0__9_;
   wire U_dsdc_bm_row_addr_0__10_;
   wire U_dsdc_bm_row_addr_0__11_;
   wire U_dsdc_bm_row_addr_0__12_;
   wire U_dsdc_bm_row_addr_0__13_;
   wire U_dsdc_bm_row_addr_0__14_;
   wire U_dsdc_bm_row_addr_0__15_;
   wire U_dsdc_bm_row_addr_1__0_;
   wire U_dsdc_bm_row_addr_1__1_;
   wire U_dsdc_bm_row_addr_1__2_;
   wire U_dsdc_bm_row_addr_1__3_;
   wire U_dsdc_bm_row_addr_1__4_;
   wire U_dsdc_bm_row_addr_1__5_;
   wire U_dsdc_bm_row_addr_1__6_;
   wire U_dsdc_bm_row_addr_1__7_;
   wire U_dsdc_bm_row_addr_1__8_;
   wire U_dsdc_bm_row_addr_1__9_;
   wire U_dsdc_bm_row_addr_1__10_;
   wire U_dsdc_bm_row_addr_1__11_;
   wire U_dsdc_bm_row_addr_1__12_;
   wire U_dsdc_bm_row_addr_1__13_;
   wire U_dsdc_bm_row_addr_1__14_;
   wire U_dsdc_bm_row_addr_1__15_;
   wire U_dsdc_bm_row_addr_2__0_;
   wire U_dsdc_bm_row_addr_2__1_;
   wire U_dsdc_bm_row_addr_2__2_;
   wire U_dsdc_bm_row_addr_2__3_;
   wire U_dsdc_bm_row_addr_2__4_;
   wire U_dsdc_bm_row_addr_2__5_;
   wire U_dsdc_bm_row_addr_2__6_;
   wire U_dsdc_bm_row_addr_2__7_;
   wire U_dsdc_bm_row_addr_2__8_;
   wire U_dsdc_bm_row_addr_2__9_;
   wire U_dsdc_bm_row_addr_2__10_;
   wire U_dsdc_bm_row_addr_2__11_;
   wire U_dsdc_bm_row_addr_2__12_;
   wire U_dsdc_bm_row_addr_2__13_;
   wire U_dsdc_bm_row_addr_2__14_;
   wire U_dsdc_bm_row_addr_2__15_;
   wire U_dsdc_bm_row_addr_3__0_;
   wire U_dsdc_bm_row_addr_3__1_;
   wire U_dsdc_bm_row_addr_3__2_;
   wire U_dsdc_bm_row_addr_3__3_;
   wire U_dsdc_bm_row_addr_3__4_;
   wire U_dsdc_bm_row_addr_3__5_;
   wire U_dsdc_bm_row_addr_3__6_;
   wire U_dsdc_bm_row_addr_3__7_;
   wire U_dsdc_bm_row_addr_3__8_;
   wire U_dsdc_bm_row_addr_3__9_;
   wire U_dsdc_bm_row_addr_3__10_;
   wire U_dsdc_bm_row_addr_3__11_;
   wire U_dsdc_bm_row_addr_3__12_;
   wire U_dsdc_bm_row_addr_3__13_;
   wire U_dsdc_bm_row_addr_3__14_;
   wire U_dsdc_bm_row_addr_3__15_;
   wire U_dsdc_N4253;
   wire U_dsdc_N4252;
   wire U_dsdc_N4250;
   wire U_dsdc_N4248;
   wire U_dsdc_N4246;
   wire U_dsdc_N4244;
   wire U_dsdc_N4242;
   wire U_dsdc_N4241;
   wire U_dsdc_N4240;
   wire U_dsdc_N4239;
   wire U_dsdc_N4229;
   wire U_dsdc_N4228;
   wire U_dsdc_t_xp_cnt_0_;
   wire U_dsdc_t_xp_cnt_1_;
   wire U_dsdc_N4174;
   wire U_dsdc_N4141;
   wire U_dsdc_N4140;
   wire U_dsdc_N4139;
   wire U_dsdc_N4129;
   wire U_dsdc_N4128;
   wire U_dsdc_N4127;
   wire U_dsdc_N2002;
   wire U_dsdc_N1991;
   wire U_dsdc_N1990;
   wire U_dsdc_N1989;
   wire U_dsdc_N1988;
   wire U_dsdc_N1987;
   wire U_dsdc_N1767;
   wire U_dsdc_N1766;
   wire U_dsdc_N1765;
   wire U_dsdc_N1764;
   wire U_dsdc_N1763;
   wire U_dsdc_N1762;
   wire U_dsdc_rcd_cnt_0_;
   wire U_dsdc_rcd_cnt_2_;
   wire U_dsdc_bm_num_open_bank_0_;
   wire U_dsdc_bm_num_open_bank_1_;
   wire U_dsdc_bm_num_open_bank_2_;
   wire U_dsdc_bm_num_open_bank_3_;
   wire U_dsdc_bm_num_open_bank_4_;
   wire U_dsdc_cas_latency_cnt_0_;
   wire U_dsdc_cas_latency_cnt_1_;
   wire U_dsdc_cas_latency_cnt_2_;
   wire U_dsdc_cas_latency_cnt_3_;
   wire U_dsdc_oldest_bank_0_;
   wire U_dsdc_oldest_bank_1_;
   wire U_dsdc_bm_ras_cnt_max_0_;
   wire U_dsdc_bm_ras_cnt_max_1_;
   wire U_dsdc_bm_ras_cnt_max_2_;
   wire U_dsdc_bm_ras_cnt_max_3_;
   wire U_dsdc_bm_bank_status_0_;
   wire U_dsdc_bm_bank_status_1_;
   wire U_dsdc_bm_bank_status_2_;
   wire U_dsdc_bm_bank_status_3_;
   wire U_dsdc_init_cnt_0_;
   wire U_dsdc_init_cnt_1_;
   wire U_dsdc_init_cnt_2_;
   wire U_dsdc_init_cnt_3_;
   wire U_dsdc_init_cnt_4_;
   wire U_dsdc_init_cnt_5_;
   wire U_dsdc_init_cnt_6_;
   wire U_dsdc_init_cnt_7_;
   wire U_dsdc_init_cnt_8_;
   wire U_dsdc_init_cnt_9_;
   wire U_dsdc_init_cnt_10_;
   wire U_dsdc_init_cnt_11_;
   wire U_dsdc_init_cnt_12_;
   wire U_dsdc_init_cnt_13_;
   wire U_dsdc_init_cnt_14_;
   wire U_dsdc_init_cnt_15_;
   wire U_dsdc_xsr_cnt_0_;
   wire U_dsdc_xsr_cnt_1_;
   wire U_dsdc_xsr_cnt_2_;
   wire U_dsdc_xsr_cnt_3_;
   wire U_dsdc_xsr_cnt_4_;
   wire U_dsdc_xsr_cnt_5_;
   wire U_dsdc_xsr_cnt_7_;
   wire U_dsdc_xsr_cnt_8_;
   wire U_dsdc_mrd_cnt_0_;
   wire U_dsdc_mrd_cnt_1_;
   wire U_dsdc_close_bank_addr_0_;
   wire U_dsdc_close_bank_addr_1_;
   wire U_dsdc_bm_close_bank_0_;
   wire U_dsdc_bm_close_bank_1_;
   wire U_dsdc_bm_close_bank_2_;
   wire U_dsdc_bm_close_bank_3_;
   wire U_dsdc_write_start_nxt;
   wire U_dsdc_wrapped_pop_flag_nxt;
   wire U_dsdc_cas_latency_1_;
   wire U_dsdc_cas_latency_2_;
   wire U_dsdc_N430;
   wire U_dsdc_auto_ref_en_nxt;
   wire U_dsdc_N429;
   wire U_dsdc_r_bm_close_all;
   wire U_dsdc_r_close_bank_addr_0_;
   wire U_dsdc_r_close_bank_addr_1_;
   wire U_dsdc_r_bm_close_bank_0_;
   wire U_dsdc_r_bm_close_bank_1_;
   wire U_dsdc_r_bm_close_bank_2_;
   wire U_dsdc_r_bm_close_bank_3_;
   wire U_dsdc_data_flag;
   wire U_dsdc_delta_delay_0_;
   wire U_dsdc_delta_delay_1_;
   wire U_dsdc_delta_delay_2_;
   wire U_dsdc_wrapped_pop_flag;
   wire U_dsdc_early_term_flag;
   wire U_dsdc_i_col_addr_1_;
   wire U_dsdc_r_cas_latency_0_;
   wire U_dsdc_r_cas_latency_1_;
   wire U_dsdc_r_cas_latency_2_;
   wire U_dsdc_r_cas_latency_3_;
   wire U_dsdc_r_wrapped_burst;
   wire U_dsdc_r_burst_size_0_;
   wire U_dsdc_r_burst_size_1_;
   wire U_dsdc_r_burst_size_2_;
   wire U_dsdc_r_burst_size_3_;
   wire U_dsdc_r_burst_size_4_;
   wire U_dsdc_r_burst_size_5_;
   wire U_dsdc_r_rw;
   wire U_dsdc_r_col_addr_1_;
   wire U_dsdc_r_row_addr_0_;
   wire U_dsdc_r_row_addr_1_;
   wire U_dsdc_r_row_addr_2_;
   wire U_dsdc_r_row_addr_3_;
   wire U_dsdc_r_row_addr_4_;
   wire U_dsdc_r_row_addr_5_;
   wire U_dsdc_r_row_addr_6_;
   wire U_dsdc_r_row_addr_7_;
   wire U_dsdc_r_row_addr_8_;
   wire U_dsdc_r_row_addr_9_;
   wire U_dsdc_r_row_addr_10_;
   wire U_dsdc_r_row_addr_11_;
   wire U_dsdc_r_row_addr_12_;
   wire U_dsdc_r_row_addr_13_;
   wire U_dsdc_r_row_addr_14_;
   wire U_dsdc_r_row_addr_15_;
   wire U_dsdc_r_chip_slct_0_;
   wire U_dsdc_data_cnt_0_;
   wire U_dsdc_data_cnt_1_;
   wire U_dsdc_data_cnt_2_;
   wire U_dsdc_data_cnt_3_;
   wire U_dsdc_data_cnt_4_;
   wire U_dsdc_data_cnt_5_;
   wire U_dsdc_cas_cnt_1_;
   wire U_dsdc_cas_cnt_2_;
   wire U_dsdc_cas_cnt_3_;
   wire U_dsdc_cas_cnt_4_;
   wire U_dsdc_cas_cnt_5_;
   wire U_dsdc_row_cnt_0_;
   wire U_dsdc_row_cnt_1_;
   wire U_dsdc_row_cnt_2_;
   wire U_dsdc_row_cnt_3_;
   wire U_dsdc_row_cnt_4_;
   wire U_dsdc_row_cnt_5_;
   wire U_dsdc_row_cnt_6_;
   wire U_dsdc_row_cnt_7_;
   wire U_dsdc_row_cnt_8_;
   wire U_dsdc_row_cnt_9_;
   wire U_dsdc_row_cnt_10_;
   wire U_dsdc_row_cnt_11_;
   wire U_dsdc_row_cnt_12_;
   wire U_dsdc_row_cnt_13_;
   wire U_dsdc_row_cnt_14_;
   wire U_dsdc_row_cnt_15_;
   wire U_dsdc_num_init_ref_cnt_0_;
   wire U_dsdc_num_init_ref_cnt_1_;
   wire U_dsdc_num_init_ref_cnt_2_;
   wire U_dsdc_num_init_ref_cnt_3_;
   wire U_dsdc_wtr_cnt_0_;
   wire U_dsdc_wtr_cnt_2_;
   wire U_dsdc_wr_cnt_0_;
   wire U_dsdc_wr_cnt_2_;
   wire U_dsdc_term_cnt_0_;
   wire U_dsdc_term_cnt_1_;
   wire U_dsdc_term_cnt_2_;
   wire U_dsdc_term_cnt_3_;
   wire U_dsdc_term_cnt_4_;
   wire U_dsdc_rp_cnt2_2_;
   wire U_dsdc_rp_cnt1_0_;
   wire U_dsdc_rp_cnt1_1_;
   wire U_dsdc_rp_cnt1_2_;
   wire U_dsdc_rcar_cnt2_0_;
   wire U_dsdc_rcar_cnt2_1_;
   wire U_dsdc_rcar_cnt2_2_;
   wire U_dsdc_rcar_cnt2_3_;
   wire U_dsdc_rcar_cnt1_0_;
   wire U_dsdc_rcar_cnt1_1_;
   wire U_dsdc_rcar_cnt1_2_;
   wire U_dsdc_rcar_cnt1_3_;
   wire U_dsdc_operation_cs_0_;
   wire U_dsdc_operation_cs_1_;
   wire U_dsdc_operation_cs_2_;
   wire U_dsdc_operation_cs_3_;
   wire U_dsdc_access_cs_0_;
   wire U_dsdc_access_cs_1_;
   wire U_dsdc_access_cs_2_;
   wire U_dsdc_access_cs_3_;
   wire U_dsdc_access_cs_4_;
   wire U_dsdc_n2097;
   wire U_dsdc_n2096;
   wire U_dsdc_n2095;
   wire U_dsdc_n2094;
   wire U_dsdc_n2093;
   wire U_cr_n550;
   wire U_cr_n549;
   wire U_cr_n548;
   wire U_cr_n547;
   wire U_cr_n546;
   wire U_cr_n545;
   wire U_cr_n544;
   wire U_cr_n543;
   wire U_cr_n542;
   wire U_cr_n541;
   wire U_cr_n540;
   wire U_cr_n539;
   wire U_cr_n538;
   wire U_cr_n537;
   wire U_cr_n536;
   wire U_cr_n535;
   wire U_cr_n534;
   wire U_cr_n533;
   wire U_cr_n532;
   wire U_cr_n531;
   wire U_cr_n530;
   wire U_cr_n529;
   wire U_cr_n528;
   wire U_cr_n527;
   wire U_cr_n526;
   wire U_cr_n525;
   wire U_cr_n524;
   wire U_cr_n523;
   wire U_cr_n522;
   wire U_cr_n521;
   wire U_cr_n520;
   wire U_cr_n519;
   wire U_cr_n518;
   wire U_cr_n517;
   wire U_cr_n516;
   wire U_cr_n515;
   wire U_cr_n514;
   wire U_cr_n513;
   wire U_cr_n512;
   wire U_cr_n511;
   wire U_cr_n510;
   wire U_cr_n509;
   wire U_cr_n508;
   wire U_cr_n507;
   wire U_cr_n506;
   wire U_cr_n505;
   wire U_cr_n504;
   wire U_cr_n503;
   wire U_cr_n502;
   wire U_cr_n501;
   wire U_cr_n500;
   wire U_cr_n499;
   wire U_cr_n498;
   wire U_cr_n497;
   wire U_cr_n496;
   wire U_cr_n495;
   wire U_cr_n494;
   wire U_cr_n493;
   wire U_cr_n492;
   wire U_cr_n491;
   wire U_cr_n490;
   wire U_cr_n489;
   wire U_cr_n488;
   wire U_cr_n487;
   wire U_cr_n486;
   wire U_cr_n485;
   wire U_cr_n484;
   wire U_cr_n483;
   wire U_cr_n482;
   wire U_cr_n481;
   wire U_cr_n480;
   wire U_cr_n479;
   wire U_cr_n478;
   wire U_cr_n477;
   wire U_cr_n476;
   wire U_cr_n475;
   wire U_cr_n474;
   wire U_cr_n473;
   wire U_cr_n472;
   wire U_cr_n471;
   wire U_cr_n470;
   wire U_cr_n469;
   wire U_cr_n468;
   wire U_cr_n467;
   wire U_cr_n466;
   wire U_cr_n465;
   wire U_cr_n464;
   wire U_cr_n463;
   wire U_cr_n462;
   wire U_cr_n461;
   wire U_cr_n460;
   wire U_cr_n459;
   wire U_cr_n458;
   wire U_cr_n457;
   wire U_cr_n456;
   wire U_cr_n455;
   wire U_cr_n454;
   wire U_cr_n453;
   wire U_cr_n452;
   wire U_cr_n451;
   wire U_cr_n450;
   wire U_cr_n449;
   wire U_cr_n448;
   wire U_cr_n447;
   wire U_cr_n446;
   wire U_cr_n445;
   wire U_cr_n444;
   wire U_cr_n443;
   wire U_cr_n442;
   wire U_cr_n441;
   wire U_cr_n440;
   wire U_cr_n439;
   wire U_cr_n438;
   wire U_cr_n437;
   wire U_cr_n436;
   wire U_cr_n435;
   wire U_cr_n434;
   wire U_cr_n433;
   wire U_cr_n432;
   wire U_cr_n431;
   wire U_cr_n430;
   wire U_cr_n429;
   wire U_cr_n428;
   wire U_cr_n427;
   wire U_cr_n426;
   wire U_cr_n425;
   wire U_cr_n424;
   wire U_cr_n423;
   wire U_cr_n422;
   wire U_cr_n421;
   wire U_cr_n420;
   wire U_cr_n419;
   wire U_cr_n418;
   wire U_cr_n417;
   wire U_cr_n416;
   wire U_cr_n415;
   wire U_cr_n414;
   wire U_cr_n413;
   wire U_cr_n412;
   wire U_cr_n411;
   wire U_cr_n410;
   wire U_cr_n409;
   wire U_cr_n408;
   wire U_cr_n407;
   wire U_cr_n406;
   wire U_cr_n405;
   wire U_cr_n404;
   wire U_cr_n403;
   wire U_cr_n402;
   wire U_cr_n401;
   wire U_cr_n400;
   wire U_cr_n399;
   wire U_cr_n398;
   wire U_cr_n397;
   wire U_cr_n396;
   wire U_cr_n395;
   wire U_cr_n394;
   wire U_cr_n393;
   wire U_cr_n392;
   wire U_cr_n391;
   wire U_cr_n390;
   wire U_cr_n389;
   wire U_cr_n388;
   wire U_cr_n387;
   wire U_cr_n386;
   wire U_cr_n385;
   wire U_cr_n384;
   wire U_cr_n383;
   wire U_cr_n382;
   wire U_cr_n381;
   wire U_cr_n380;
   wire U_cr_n379;
   wire U_cr_n378;
   wire U_cr_n377;
   wire U_cr_n376;
   wire U_cr_n375;
   wire U_cr_n374;
   wire U_cr_n373;
   wire U_cr_n372;
   wire U_cr_n371;
   wire U_cr_n370;
   wire U_cr_n369;
   wire U_cr_n368;
   wire U_cr_n367;
   wire U_cr_n366;
   wire U_cr_n365;
   wire U_cr_n364;
   wire U_cr_n363;
   wire U_cr_n362;
   wire U_cr_n361;
   wire U_cr_n360;
   wire U_cr_n359;
   wire U_cr_n358;
   wire U_cr_n357;
   wire U_cr_n356;
   wire U_cr_n355;
   wire U_cr_n354;
   wire U_cr_n353;
   wire U_cr_n352;
   wire U_cr_n351;
   wire U_cr_n350;
   wire U_cr_n349;
   wire U_cr_n348;
   wire U_cr_n347;
   wire U_cr_n346;
   wire U_cr_n345;
   wire U_cr_n344;
   wire U_cr_n343;
   wire U_cr_n342;
   wire U_cr_n341;
   wire U_cr_n340;
   wire U_cr_n339;
   wire U_cr_n338;
   wire U_cr_n337;
   wire U_cr_n336;
   wire U_cr_n335;
   wire U_cr_n334;
   wire U_cr_n333;
   wire U_cr_n332;
   wire U_cr_n331;
   wire U_cr_n330;
   wire U_cr_n329;
   wire U_cr_n328;
   wire U_cr_n327;
   wire U_cr_n326;
   wire U_cr_n325;
   wire U_cr_n324;
   wire U_cr_n323;
   wire U_cr_n322;
   wire U_cr_n321;
   wire U_cr_n320;
   wire U_cr_n319;
   wire U_cr_n318;
   wire U_cr_n317;
   wire U_cr_n316;
   wire U_cr_n315;
   wire U_cr_n314;
   wire U_cr_n313;
   wire U_cr_n312;
   wire U_cr_n311;
   wire U_cr_n310;
   wire U_cr_n309;
   wire U_cr_n308;
   wire U_cr_n307;
   wire U_cr_n306;
   wire U_cr_n305;
   wire U_cr_n304;
   wire U_cr_n303;
   wire U_cr_n302;
   wire U_cr_n301;
   wire U_cr_n300;
   wire U_cr_n299;
   wire U_cr_n298;
   wire U_cr_n297;
   wire U_cr_n296;
   wire U_cr_n295;
   wire U_cr_n294;
   wire U_cr_n293;
   wire U_cr_n292;
   wire U_cr_n291;
   wire U_cr_n290;
   wire U_cr_n289;
   wire U_cr_n288;
   wire U_cr_n287;
   wire U_cr_n286;
   wire U_cr_n285;
   wire U_cr_n284;
   wire U_cr_n283;
   wire U_cr_n282;
   wire U_cr_n281;
   wire U_cr_n280;
   wire U_cr_n279;
   wire U_cr_n278;
   wire U_cr_n277;
   wire U_cr_n276;
   wire U_cr_n275;
   wire U_cr_n274;
   wire U_cr_n273;
   wire U_cr_n272;
   wire U_cr_n271;
   wire U_cr_n270;
   wire U_cr_n269;
   wire U_cr_n268;
   wire U_cr_n267;
   wire U_cr_n266;
   wire U_cr_n265;
   wire U_cr_n264;
   wire U_cr_n263;
   wire U_cr_n262;
   wire U_cr_n261;
   wire U_cr_n260;
   wire U_cr_n259;
   wire U_cr_n258;
   wire U_cr_n257;
   wire U_cr_n256;
   wire U_cr_n255;
   wire U_cr_n254;
   wire U_cr_n253;
   wire U_cr_n252;
   wire U_cr_n251;
   wire U_cr_n250;
   wire U_cr_n249;
   wire U_cr_n248;
   wire U_cr_n247;
   wire U_cr_n246;
   wire U_cr_n245;
   wire U_cr_n244;
   wire U_cr_n243;
   wire U_cr_n242;
   wire U_cr_n241;
   wire U_cr_n240;
   wire U_cr_n239;
   wire U_cr_n238;
   wire U_cr_n237;
   wire U_cr_n236;
   wire U_cr_n235;
   wire U_cr_n234;
   wire U_cr_n233;
   wire U_cr_n232;
   wire U_cr_n231;
   wire U_cr_n230;
   wire U_cr_n229;
   wire U_cr_n228;
   wire U_cr_n227;
   wire U_cr_n226;
   wire U_cr_n225;
   wire U_cr_n224;
   wire U_cr_n223;
   wire U_cr_n222;
   wire U_cr_n221;
   wire U_cr_n220;
   wire U_cr_n219;
   wire U_cr_n218;
   wire U_cr_n217;
   wire U_cr_n216;
   wire U_cr_n215;
   wire U_cr_n214;
   wire U_cr_n213;
   wire U_cr_n212;
   wire U_cr_n211;
   wire U_cr_n210;
   wire U_cr_n209;
   wire U_cr_n208;
   wire U_cr_n207;
   wire U_cr_n206;
   wire U_cr_n205;
   wire U_cr_n204;
   wire U_cr_n203;
   wire U_cr_n202;
   wire U_cr_n201;
   wire U_cr_n200;
   wire U_cr_n199;
   wire U_cr_n198;
   wire U_cr_n197;
   wire U_cr_n196;
   wire U_cr_n195;
   wire U_cr_n194;
   wire U_cr_n193;
   wire U_cr_n192;
   wire U_cr_n191;
   wire U_cr_n190;
   wire U_cr_n189;
   wire U_cr_n188;
   wire U_cr_n187;
   wire U_cr_n186;
   wire U_cr_n185;
   wire U_cr_n184;
   wire U_cr_n182;
   wire U_cr_n181;
   wire U_cr_n180;
   wire U_cr_n179;
   wire U_cr_n178;
   wire U_cr_n177;
   wire U_cr_n176;
   wire U_cr_n175;
   wire U_cr_n174;
   wire U_cr_n171;
   wire U_cr_n170;
   wire U_cr_n169;
   wire U_cr_n168;
   wire U_cr_n167;
   wire U_cr_n166;
   wire U_cr_n165;
   wire U_cr_n164;
   wire U_cr_n163;
   wire U_cr_n162;
   wire U_cr_n161;
   wire U_cr_n160;
   wire U_cr_n159;
   wire U_cr_n158;
   wire U_cr_n157;
   wire U_cr_n156;
   wire U_cr_n155;
   wire U_cr_n154;
   wire U_cr_n153;
   wire U_cr_n152;
   wire U_cr_n151;
   wire U_cr_n150;
   wire U_cr_n149;
   wire U_cr_n148;
   wire U_cr_n147;
   wire U_cr_n146;
   wire U_cr_n145;
   wire U_cr_n144;
   wire U_cr_n143;
   wire U_cr_n142;
   wire U_cr_n141;
   wire U_cr_n140;
   wire U_cr_n139;
   wire U_cr_n138;
   wire U_cr_n137;
   wire U_cr_n136;
   wire U_cr_n135;
   wire U_cr_n134;
   wire U_cr_n133;
   wire U_cr_n132;
   wire U_cr_n131;
   wire U_cr_n130;
   wire U_cr_n129;
   wire U_cr_n128;
   wire U_cr_n127;
   wire U_cr_n126;
   wire U_cr_n125;
   wire U_cr_n124;
   wire U_cr_n123;
   wire U_cr_n122;
   wire U_cr_n121;
   wire U_cr_n120;
   wire U_cr_n119;
   wire U_cr_n118;
   wire U_cr_n117;
   wire U_cr_n116;
   wire U_cr_n115;
   wire U_cr_n114;
   wire U_cr_n113;
   wire U_cr_n112;
   wire U_cr_n111;
   wire U_cr_n110;
   wire U_cr_n109;
   wire U_cr_n108;
   wire U_cr_n107;
   wire U_cr_n106;
   wire U_cr_n105;
   wire U_cr_n104;
   wire U_cr_n103;
   wire U_cr_n102;
   wire U_cr_n101;
   wire U_cr_n100;
   wire U_cr_n97;
   wire U_cr_n72;
   wire U_cr_n71;
   wire U_cr_n70;
   wire U_cr_n69;
   wire U_cr_n68;
   wire U_cr_n67;
   wire U_cr_n66;
   wire U_cr_n65;
   wire U_cr_n64;
   wire U_cr_n63;
   wire U_cr_n61;
   wire U_cr_n60;
   wire U_cr_n59;
   wire U_cr_n58;
   wire U_cr_n57;
   wire U_cr_n56;
   wire U_cr_n55;
   wire U_cr_n54;
   wire U_cr_n53;
   wire U_cr_n52;
   wire U_cr_n51;
   wire U_cr_n50;
   wire U_cr_n49;
   wire U_cr_n48;
   wire U_cr_n47;
   wire U_cr_n46;
   wire U_cr_n45;
   wire U_cr_n44;
   wire U_cr_n43;
   wire U_cr_n42;
   wire U_cr_n41;
   wire U_cr_n40;
   wire U_cr_n39;
   wire U_cr_n38;
   wire U_cr_n37;
   wire U_cr_n36;
   wire U_cr_n35;
   wire U_cr_n34;
   wire U_cr_n33;
   wire U_cr_n32;
   wire U_cr_n31;
   wire U_cr_n30;
   wire U_cr_n29;
   wire U_cr_n28;
   wire U_cr_n27;
   wire U_cr_n26;
   wire U_cr_n25;
   wire U_cr_n24;
   wire U_cr_n23;
   wire U_cr_n22;
   wire U_cr_n21;
   wire U_cr_n20;
   wire U_cr_n19;
   wire U_cr_n18;
   wire U_cr_n17;
   wire U_cr_n16;
   wire U_cr_n13;
   wire U_cr_n12;
   wire U_cr_n11;
   wire U_cr_n10;
   wire U_cr_n9;
   wire U_cr_n8;
   wire U_cr_n7;
   wire U_cr_n6;
   wire U_cr_n5;
   wire U_cr_n4;
   wire U_cr_n3;
   wire U_cr_n2;
   wire U_cr_n1;
   wire U_cr_n99;
   wire U_cr_n98;
   wire U_cr_n96;
   wire U_cr_n95;
   wire U_cr_n94;
   wire U_cr_n93;
   wire U_cr_n92;
   wire U_cr_n91;
   wire U_cr_n90;
   wire U_cr_n89;
   wire U_cr_n88;
   wire U_cr_n87;
   wire U_cr_n86;
   wire U_cr_n85;
   wire U_cr_n84;
   wire U_cr_n83;
   wire U_cr_n82;
   wire U_cr_n81;
   wire U_cr_n80;
   wire U_cr_n79;
   wire U_cr_n78;
   wire U_cr_n77;
   wire U_cr_n76;
   wire U_cr_n75;
   wire U_cr_n74;
   wire U_cr_n73;
   wire U_cr_cr_cs_0_;
   wire U_cr_cr_cs_1_;
   wire U_cr_cr_cs_2_;
   wire U_cr_s_sda_d;
   wire U_cr_s_sda_d1;
   wire U_cr_N745;
   wire U_cr_N740;
   wire U_cr_N739;
   wire U_cr_N738;
   wire U_cr_N737;
   wire U_cr_N736;
   wire U_cr_N735;
   wire U_cr_N734;
   wire U_cr_N733;
   wire U_cr_N700;
   wire U_cr_N699;
   wire U_cr_N698;
   wire U_cr_N697;
   wire U_cr_N696;
   wire U_cr_N695;
   wire U_cr_N694;
   wire U_cr_N693;
   wire U_cr_N692;
   wire U_cr_N691;
   wire U_cr_N690;
   wire U_cr_N689;
   wire U_cr_N688;
   wire U_cr_N655;
   wire U_cr_N654;
   wire U_cr_N653;
   wire U_cr_N652;
   wire U_cr_N651;
   wire U_cr_N650;
   wire U_cr_N649;
   wire U_cr_N648;
   wire U_cr_N647;
   wire U_cr_N646;
   wire U_cr_N645;
   wire U_cr_N644;
   wire U_cr_N643;
   wire U_cr_N642;
   wire U_cr_N641;
   wire U_cr_N640;
   wire U_cr_N639;
   wire U_cr_N638;
   wire U_cr_N637;
   wire U_cr_N636;
   wire U_cr_N635;
   wire U_cr_N634;
   wire U_cr_N577;
   wire U_cr_N576;
   wire U_cr_N574;
   wire U_cr_N573;
   wire U_cr_N572;
   wire U_cr_N571;
   wire U_cr_N567;
   wire U_cr_N566;
   wire U_cr_N565;
   wire U_cr_N564;
   wire U_cr_N563;
   wire U_cr_N562;
   wire U_cr_N561;
   wire U_cr_N560;
   wire U_cr_N559;
   wire U_cr_N558;
   wire U_cr_N557;
   wire U_cr_N556;
   wire U_cr_N555;
   wire U_cr_N554;
   wire U_cr_N553;
   wire U_cr_N552;
   wire U_cr_N551;
   wire U_cr_N550;
   wire U_cr_N479;
   wire U_cr_N478;
   wire U_cr_N477;
   wire U_cr_N476;
   wire U_cr_N475;
   wire U_cr_N474;
   wire U_cr_N473;
   wire U_cr_N472;
   wire U_cr_N471;
   wire U_cr_N470;
   wire U_cr_N469;
   wire U_cr_N468;
   wire U_cr_N467;
   wire U_cr_N466;
   wire U_cr_N465;
   wire U_cr_N464;
   wire U_cr_N420;
   wire U_cr_N419;
   wire U_cr_N418;
   wire U_cr_N417;
   wire U_cr_N416;
   wire U_cr_N415;
   wire U_cr_N414;
   wire U_cr_N413;
   wire U_cr_N412;
   wire U_cr_N411;
   wire U_cr_N410;
   wire U_cr_N409;
   wire U_cr_N408;
   wire U_cr_N407;
   wire U_cr_N406;
   wire U_cr_N405;
   wire U_cr_N404;
   wire U_cr_N403;
   wire U_cr_N402;
   wire U_cr_N401;
   wire U_cr_N400;
   wire U_cr_N399;
   wire U_cr_N398;
   wire U_cr_N397;
   wire U_cr_N396;
   wire U_cr_N395;
   wire U_cr_N394;
   wire U_cr_N393;
   wire U_cr_N392;
   wire U_cr_N391;
   wire U_cr_N390;
   wire U_cr_N389;
   wire U_cr_N315;
   wire U_cr_N313;
   wire U_cr_N312;
   wire U_cr_N311;
   wire U_cr_N310;
   wire U_cr_N308;
   wire U_cr_N307;
   wire U_cr_N306;
   wire U_cr_N305;
   wire U_cr_N304;
   wire U_cr_N303;
   wire U_cr_N302;
   wire U_cr_N301;
   wire U_cr_N300;
   wire U_cr_N299;
   wire U_cr_N298;
   wire U_cr_sctlr_default_11;
   wire U_cr_stmg0r_0_;
   wire U_cr_stmg0r_1_;
   wire U_cr_stmg0r_26;
   wire U_cr_sctlr_12_;
   wire U_cr_sctlr_13_;
   wire U_cr_sctlr_14_;
   wire U_cr_sctlr_15_;
   wire U_cr_sctlr_16_;
   wire U_cr_n572;
   wire U_cr_n571;
   wire U_cr_n570;
   wire U_cr_n569;
   wire U_cr_n568;
   wire U_cr_n567;
   wire U_cr_n566;
   wire U_cr_n565;
   wire U_cr_n564;
   wire U_cr_n563;
   wire U_cr_n562;
   wire U_cr_n561;
   wire U_cr_n560;
   wire U_cr_n559;
   wire U_cr_n558;
   wire U_cr_n557;
   wire U_cr_n556;
   wire U_cr_n555;
   wire U_cr_n554;
   wire U_cr_n553;
   wire U_cr_n552;
   wire U_cr_n551;
   wire U_addrdec_n311;
   wire U_addrdec_n310;
   wire U_addrdec_n309;
   wire U_addrdec_n303;
   wire U_addrdec_n302;
   wire U_addrdec_n301;
   wire U_addrdec_n300;
   wire U_addrdec_n299;
   wire U_addrdec_n298;
   wire U_addrdec_n297;
   wire U_addrdec_n296;
   wire U_addrdec_n295;
   wire U_addrdec_n294;
   wire U_addrdec_n293;
   wire U_addrdec_n292;
   wire U_addrdec_n291;
   wire U_addrdec_n290;
   wire U_addrdec_n287;
   wire U_addrdec_n286;
   wire U_addrdec_n285;
   wire U_addrdec_n284;
   wire U_addrdec_n283;
   wire U_addrdec_n282;
   wire U_addrdec_n281;
   wire U_addrdec_n280;
   wire U_addrdec_n278;
   wire U_addrdec_n277;
   wire U_addrdec_n276;
   wire U_addrdec_n275;
   wire U_addrdec_n274;
   wire U_addrdec_n273;
   wire U_addrdec_n272;
   wire U_addrdec_n271;
   wire U_addrdec_n270;
   wire U_addrdec_n269;
   wire U_addrdec_n268;
   wire U_addrdec_n267;
   wire U_addrdec_n266;
   wire U_addrdec_n265;
   wire U_addrdec_n264;
   wire U_addrdec_n263;
   wire U_addrdec_n262;
   wire U_addrdec_n261;
   wire U_addrdec_n260;
   wire U_addrdec_n259;
   wire U_addrdec_n258;
   wire U_addrdec_n257;
   wire U_addrdec_n256;
   wire U_addrdec_n255;
   wire U_addrdec_n254;
   wire U_addrdec_n253;
   wire U_addrdec_n252;
   wire U_addrdec_n251;
   wire U_addrdec_n250;
   wire U_addrdec_n249;
   wire U_addrdec_n248;
   wire U_addrdec_n247;
   wire U_addrdec_n246;
   wire U_addrdec_n245;
   wire U_addrdec_n244;
   wire U_addrdec_n243;
   wire U_addrdec_n242;
   wire U_addrdec_n241;
   wire U_addrdec_n240;
   wire U_addrdec_n239;
   wire U_addrdec_n238;
   wire U_addrdec_n237;
   wire U_addrdec_n236;
   wire U_addrdec_n235;
   wire U_addrdec_n234;
   wire U_addrdec_n233;
   wire U_addrdec_n232;
   wire U_addrdec_n231;
   wire U_addrdec_n230;
   wire U_addrdec_n229;
   wire U_addrdec_n228;
   wire U_addrdec_n227;
   wire U_addrdec_n226;
   wire U_addrdec_n225;
   wire U_addrdec_n224;
   wire U_addrdec_n223;
   wire U_addrdec_n222;
   wire U_addrdec_n221;
   wire U_addrdec_n220;
   wire U_addrdec_n219;
   wire U_addrdec_n218;
   wire U_addrdec_n217;
   wire U_addrdec_n216;
   wire U_addrdec_n215;
   wire U_addrdec_n214;
   wire U_addrdec_n213;
   wire U_addrdec_n212;
   wire U_addrdec_n211;
   wire U_addrdec_n210;
   wire U_addrdec_n209;
   wire U_addrdec_n208;
   wire U_addrdec_n207;
   wire U_addrdec_n206;
   wire U_addrdec_n205;
   wire U_addrdec_n204;
   wire U_addrdec_n203;
   wire U_addrdec_n202;
   wire U_addrdec_n201;
   wire U_addrdec_n200;
   wire U_addrdec_n199;
   wire U_addrdec_n198;
   wire U_addrdec_n197;
   wire U_addrdec_n196;
   wire U_addrdec_n195;
   wire U_addrdec_n194;
   wire U_addrdec_n193;
   wire U_addrdec_n192;
   wire U_addrdec_n191;
   wire U_addrdec_n190;
   wire U_addrdec_n189;
   wire U_addrdec_n188;
   wire U_addrdec_n187;
   wire U_addrdec_n186;
   wire U_addrdec_n185;
   wire U_addrdec_n184;
   wire U_addrdec_n183;
   wire U_addrdec_n182;
   wire U_addrdec_n181;
   wire U_addrdec_n180;
   wire U_addrdec_n179;
   wire U_addrdec_n178;
   wire U_addrdec_n177;
   wire U_addrdec_n176;
   wire U_addrdec_n175;
   wire U_addrdec_n174;
   wire U_addrdec_n173;
   wire U_addrdec_n172;
   wire U_addrdec_n171;
   wire U_addrdec_n170;
   wire U_addrdec_n169;
   wire U_addrdec_n168;
   wire U_addrdec_n167;
   wire U_addrdec_n166;
   wire U_addrdec_n165;
   wire U_addrdec_n164;
   wire U_addrdec_n163;
   wire U_addrdec_n162;
   wire U_addrdec_n161;
   wire U_addrdec_n160;
   wire U_addrdec_n159;
   wire U_addrdec_n158;
   wire U_addrdec_n156;
   wire U_addrdec_n155;
   wire U_addrdec_n154;
   wire U_addrdec_n153;
   wire U_addrdec_n152;
   wire U_addrdec_n151;
   wire U_addrdec_n150;
   wire U_addrdec_n149;
   wire U_addrdec_n148;
   wire U_addrdec_n147;
   wire U_addrdec_n145;
   wire U_addrdec_n144;
   wire U_addrdec_n143;
   wire U_addrdec_n142;
   wire U_addrdec_n141;
   wire U_addrdec_n140;
   wire U_addrdec_n139;
   wire U_addrdec_n138;
   wire U_addrdec_n137;
   wire U_addrdec_n136;
   wire U_addrdec_n135;
   wire U_addrdec_n134;
   wire U_addrdec_n133;
   wire U_addrdec_n132;
   wire U_addrdec_n131;
   wire U_addrdec_n130;
   wire U_addrdec_n129;
   wire U_addrdec_n128;
   wire U_addrdec_n127;
   wire U_addrdec_n126;
   wire U_addrdec_n125;
   wire U_addrdec_n124;
   wire U_addrdec_n123;
   wire U_addrdec_n122;
   wire U_addrdec_n121;
   wire U_addrdec_n120;
   wire U_addrdec_n119;
   wire U_addrdec_n118;
   wire U_addrdec_n117;
   wire U_addrdec_n116;
   wire U_addrdec_n115;
   wire U_addrdec_n114;
   wire U_addrdec_n113;
   wire U_addrdec_n112;
   wire U_addrdec_n111;
   wire U_addrdec_n110;
   wire U_addrdec_n109;
   wire U_addrdec_n108;
   wire U_addrdec_n107;
   wire U_addrdec_n106;
   wire U_addrdec_n105;
   wire U_addrdec_n104;
   wire U_addrdec_n103;
   wire U_addrdec_n102;
   wire U_addrdec_n101;
   wire U_addrdec_n100;
   wire U_addrdec_n99;
   wire U_addrdec_n98;
   wire U_addrdec_n97;
   wire U_addrdec_n96;
   wire U_addrdec_n95;
   wire U_addrdec_n94;
   wire U_addrdec_n93;
   wire U_addrdec_n92;
   wire U_addrdec_n91;
   wire U_addrdec_n90;
   wire U_addrdec_n88;
   wire U_addrdec_n87;
   wire U_addrdec_n86;
   wire U_addrdec_n85;
   wire U_addrdec_n84;
   wire U_addrdec_n83;
   wire U_addrdec_n82;
   wire U_addrdec_n81;
   wire U_addrdec_n80;
   wire U_addrdec_n79;
   wire U_addrdec_n78;
   wire U_addrdec_n77;
   wire U_addrdec_n76;
   wire U_addrdec_n75;
   wire U_addrdec_n74;
   wire U_addrdec_n73;
   wire U_addrdec_n71;
   wire U_addrdec_n70;
   wire U_addrdec_n67;
   wire U_addrdec_n66;
   wire U_addrdec_n65;
   wire U_addrdec_n64;
   wire U_addrdec_n63;
   wire U_addrdec_n62;
   wire U_addrdec_n61;
   wire U_addrdec_n60;
   wire U_addrdec_n59;
   wire U_addrdec_n57;
   wire U_addrdec_n56;
   wire U_addrdec_n54;
   wire U_addrdec_n53;
   wire U_addrdec_n44;
   wire U_addrdec_n43;
   wire U_addrdec_n42;
   wire U_addrdec_n41;
   wire U_addrdec_n40;
   wire U_addrdec_n39;
   wire U_addrdec_n38;
   wire U_addrdec_n37;
   wire U_addrdec_n36;
   wire U_addrdec_n35;
   wire U_addrdec_n34;
   wire U_addrdec_n32;
   wire U_addrdec_n30;
   wire U_addrdec_n28;
   wire U_addrdec_n27;
   wire U_addrdec_n26;
   wire U_addrdec_n25;
   wire U_addrdec_n24;
   wire U_addrdec_n23;
   wire U_addrdec_n22;
   wire U_addrdec_n21;
   wire U_addrdec_n20;
   wire U_addrdec_n18;
   wire U_addrdec_n17;
   wire U_addrdec_n16;
   wire U_addrdec_n15;
   wire U_addrdec_n14;
   wire U_addrdec_n13;
   wire U_addrdec_n11;
   wire U_addrdec_n10;
   wire U_addrdec_n9;
   wire U_addrdec_n7;
   wire U_addrdec_n5;
   wire U_addrdec_n4;
   wire U_addrdec_n3;
   wire U_addrdec_n2;
   wire U_addrdec_n1;
   wire U_addrdec_n348;
   wire U_addrdec_n347;
   wire U_addrdec_n346;
   wire U_addrdec_n345;
   wire U_addrdec_n58;
   wire U_addrdec_N133;
   wire U_addrdec_N131;
   wire U_addrdec_N130;
   wire U_addrdec_N129;
   wire U_addrdec_N119;
   wire U_addrdec_N111;
   wire U_addrdec_N110;
   wire U_addrdec_N109;
   wire U_addrdec_N108;
   wire U_addrdec_N107;
   wire U_addrdec_bank_addr_mask_1_;
   wire U_addrdec_bcawp_0_;
   wire U_addrdec_bcawp_1_;
   wire U_addrdec_bcawp_2_;
   wire U_addrdec_bcawp_3_;
   wire U_addrdec_bcawp_4_;
   wire U_addrdec_flash_select_0_;
   wire U_addrdec_sram_select_0_;
   wire U_addrdec_rom_select_0_;
   wire U_refctl_n127;
   wire U_refctl_n126;
   wire U_refctl_n124;
   wire U_refctl_n123;
   wire U_refctl_n122;
   wire U_refctl_n121;
   wire U_refctl_n120;
   wire U_refctl_n119;
   wire U_refctl_n118;
   wire U_refctl_n117;
   wire U_refctl_n116;
   wire U_refctl_n115;
   wire U_refctl_n114;
   wire U_refctl_n113;
   wire U_refctl_n112;
   wire U_refctl_n111;
   wire U_refctl_n110;
   wire U_refctl_n109;
   wire U_refctl_n108;
   wire U_refctl_n107;
   wire U_refctl_n106;
   wire U_refctl_n105;
   wire U_refctl_n104;
   wire U_refctl_n103;
   wire U_refctl_n102;
   wire U_refctl_n101;
   wire U_refctl_n100;
   wire U_refctl_n99;
   wire U_refctl_n98;
   wire U_refctl_n97;
   wire U_refctl_n96;
   wire U_refctl_n95;
   wire U_refctl_n94;
   wire U_refctl_n93;
   wire U_refctl_n92;
   wire U_refctl_n91;
   wire U_refctl_n90;
   wire U_refctl_n89;
   wire U_refctl_n88;
   wire U_refctl_n87;
   wire U_refctl_n86;
   wire U_refctl_n85;
   wire U_refctl_n84;
   wire U_refctl_n83;
   wire U_refctl_n82;
   wire U_refctl_n81;
   wire U_refctl_n80;
   wire U_refctl_n79;
   wire U_refctl_n78;
   wire U_refctl_n77;
   wire U_refctl_n76;
   wire U_refctl_n75;
   wire U_refctl_n74;
   wire U_refctl_n73;
   wire U_refctl_n66;
   wire U_refctl_n65;
   wire U_refctl_n64;
   wire U_refctl_n63;
   wire U_refctl_n62;
   wire U_refctl_n61;
   wire U_refctl_n60;
   wire U_refctl_n59;
   wire U_refctl_n58;
   wire U_refctl_n57;
   wire U_refctl_n56;
   wire U_refctl_n55;
   wire U_refctl_n54;
   wire U_refctl_n53;
   wire U_refctl_n52;
   wire U_refctl_n51;
   wire U_refctl_n50;
   wire U_refctl_n49;
   wire U_refctl_n48;
   wire U_refctl_n47;
   wire U_refctl_n46;
   wire U_refctl_n45;
   wire U_refctl_n44;
   wire U_refctl_n43;
   wire U_refctl_n42;
   wire U_refctl_n41;
   wire U_refctl_n40;
   wire U_refctl_n39;
   wire U_refctl_n38;
   wire U_refctl_n37;
   wire U_refctl_n36;
   wire U_refctl_n35;
   wire U_refctl_n34;
   wire U_refctl_n33;
   wire U_refctl_n32;
   wire U_refctl_n30;
   wire U_refctl_n29;
   wire U_refctl_n28;
   wire U_refctl_n27;
   wire U_refctl_n25;
   wire U_refctl_n23;
   wire U_refctl_n22;
   wire U_refctl_n21;
   wire U_refctl_n20;
   wire U_refctl_n19;
   wire U_refctl_n18;
   wire U_refctl_n17;
   wire U_refctl_n16;
   wire U_refctl_n15;
   wire U_refctl_n14;
   wire U_refctl_n12;
   wire U_refctl_n11;
   wire U_refctl_n10;
   wire U_refctl_n9;
   wire U_refctl_n8;
   wire U_refctl_n7;
   wire U_refctl_n6;
   wire U_refctl_n5;
   wire U_refctl_n4;
   wire U_refctl_n3;
   wire U_refctl_n2;
   wire U_refctl_n1;
   wire U_refctl_N31;
   wire U_refctl_N30;
   wire U_refctl_N29;
   wire U_refctl_N28;
   wire U_refctl_N27;
   wire U_refctl_N26;
   wire U_refctl_N25;
   wire U_refctl_N24;
   wire U_refctl_N23;
   wire U_refctl_N22;
   wire U_refctl_N21;
   wire U_refctl_N20;
   wire U_refctl_N19;
   wire U_refctl_N18;
   wire U_refctl_N17;
   wire U_refctl_N16;
   wire U_refctl_next_state_0_;
   wire U_refctl_ref_req_next;
   wire U_refctl_count_next_0_;
   wire U_refctl_count_next_1_;
   wire U_refctl_count_next_2_;
   wire U_refctl_count_next_3_;
   wire U_refctl_count_next_4_;
   wire U_refctl_count_next_5_;
   wire U_refctl_count_next_7_;
   wire U_refctl_count_next_9_;
   wire U_refctl_count_next_11_;
   wire U_refctl_count_next_13_;
   wire U_refctl_count_next_14_;
   wire U_refctl_count_next_15_;
   wire U_refctl_count_0_;
   wire U_refctl_count_1_;
   wire U_refctl_count_2_;
   wire U_refctl_count_3_;
   wire U_refctl_count_4_;
   wire U_refctl_count_5_;
   wire U_refctl_count_6_;
   wire U_refctl_count_7_;
   wire U_refctl_count_8_;
   wire U_refctl_count_9_;
   wire U_refctl_count_10_;
   wire U_refctl_count_11_;
   wire U_refctl_count_12_;
   wire U_refctl_count_13_;
   wire U_refctl_count_14_;
   wire U_refctl_count_15_;
   wire U_refctl_current_state_0_;
   wire U_refctl_current_state_1_;
   wire U_dmc_n70;
   wire U_dmc_n69;
   wire U_dmc_n68;
   wire U_dmc_n67;
   wire U_dmc_n66;
   wire U_dmc_n65;
   wire U_dmc_n64;
   wire U_dmc_n63;
   wire U_dmc_n62;
   wire U_dmc_n61;
   wire U_dmc_n60;
   wire U_dmc_n59;
   wire U_dmc_n58;
   wire U_dmc_n55;
   wire U_dmc_n54;
   wire U_dmc_n53;
   wire U_dmc_n52;
   wire U_dmc_n51;
   wire U_dmc_n50;
   wire U_dmc_n49;
   wire U_dmc_n48;
   wire U_dmc_n47;
   wire U_dmc_n46;
   wire U_dmc_n45;
   wire U_dmc_n44;
   wire U_dmc_n43;
   wire U_dmc_n42;
   wire U_dmc_n41;
   wire U_dmc_n40;
   wire U_dmc_n39;
   wire U_dmc_n35;
   wire U_dmc_n34;
   wire U_dmc_n33;
   wire U_dmc_n32;
   wire U_dmc_n31;
   wire U_dmc_n30;
   wire U_dmc_n29;
   wire U_dmc_n28;
   wire U_dmc_n27;
   wire U_dmc_n26;
   wire U_dmc_n25;
   wire U_dmc_n24;
   wire U_dmc_n23;
   wire U_dmc_n22;
   wire U_dmc_n21;
   wire U_dmc_n20;
   wire U_dmc_n19;
   wire U_dmc_n18;
   wire U_dmc_n16;
   wire U_dmc_n15;
   wire U_dmc_n11;
   wire U_dmc_n10;
   wire U_dmc_n8;
   wire U_dmc_n7;
   wire U_dmc_n6;
   wire U_dmc_n5;
   wire U_dmc_n4;
   wire U_dmc_n3;
   wire U_dmc_n2;
   wire U_dmc_n1;
   wire U_dmc_n14;
   wire U_dmc_n13;
   wire U_dmc_n12;
   wire U_dmc_N24;
   wire U_dmc_N23;
   wire U_dmc_terminate;
   wire U_dmc_data_cnt_0_;
   wire U_dmc_data_cnt_1_;
   wire U_dmc_data_cnt_2_;
   wire U_dmc_data_cnt_3_;
   wire U_dmc_data_cnt_4_;
   wire U_dmc_data_cnt_5_;
   wire U_dmc_dmc_cs_0_;
   wire U_dmc_dmc_cs_1_;
   wire U_dmc_dmc_cs_2_;
   wire U_dsdc_U_minmax1_dwbb_n34;
   wire U_dsdc_U_minmax1_dwbb_n33;
   wire U_dsdc_U_minmax1_dwbb_n32;
   wire U_dsdc_U_minmax1_dwbb_n31;
   wire U_dsdc_U_minmax1_dwbb_n30;
   wire U_dsdc_U_minmax1_dwbb_n29;
   wire U_dsdc_U_minmax1_dwbb_n26;
   wire U_dsdc_U_minmax1_dwbb_n24;
   wire U_dsdc_U_minmax1_dwbb_n22;
   wire U_dsdc_U_minmax1_dwbb_n21;
   wire U_dsdc_U_minmax1_dwbb_n20;
   wire U_dsdc_U_minmax1_dwbb_n19;
   wire U_dsdc_U_minmax1_dwbb_n15;
   wire U_dsdc_U_minmax1_dwbb_n12;
   wire U_dsdc_U_minmax1_dwbb_n11;
   wire U_dsdc_U_minmax1_dwbb_n9;
   wire U_dsdc_U_minmax1_dwbb_n6;
   wire U_dsdc_U_minmax1_dwbb_n5;
   wire U_dsdc_U_minmax1_dwbb_n4;
   wire U_dsdc_U_minmax1_dwbb_n2;
   wire U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_GT_4_;
   wire U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_PI_1_;
   wire U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_0_;
   wire U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_1_;
   wire U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_;
   wire U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire [23:26] n;
   wire [31:0] miu_rd_data_reg;
   wire [31:0] cr_reg_data_out;
   wire [3:0] pre_dqm;
   wire [3:0] ad_data_mask;
   wire [3:0] cr_row_addr_width;
   wire [4:0] cr_num_open_banks;
   wire [12:0] cr_exn_mode_value;
   wire [3:0] cr_t_ras_min;
   wire [2:0] cr_t_rcd;
   wire [2:0] cr_t_rp;
   wire [3:1] cr_t_rc;
   wire [1:0] cr_t_wr;
   wire [1:0] cr_t_wtr;
   wire [3:0] cr_t_rcar;
   wire [8:0] cr_t_xsr;
   wire [15:0] cr_t_init;
   wire [3:0] cr_num_init_ref;
   wire [3:0] ad_cr_data_mask;
   wire [1:0] cr_bank_addr_width;
   wire [7:5] cr_block_size1;
   wire [15:0] cr_t_ref;
   wire [15:2] U_dsdc_num_row;
   wire [14:4] U_dsdc_i_col_addr_nxt;
   wire [5:0] U_dsdc_cas_cnt_nxt;
   wire [2:0] U_dsdc_num_init_ref_cnt_nxt;
   wire [4:0] U_dsdc_term_cnt_nxt;
   wire [2:0] U_dsdc_wtr_cnt_nxt;
   wire [2:0] U_dsdc_wr_cnt_nxt;
   wire [2:0] U_dsdc_rp_cnt2_nxt;
   wire [2:0] U_dsdc_rp_cnt1_nxt;
   wire [3:0] U_dsdc_rcar_cnt2_nxt;
   wire [3:0] U_dsdc_rcar_cnt1_nxt;
   wire [15:13] U_dsdc_s_addr_nxt_a;
   wire [3:0] U_dsdc_r_bm_open_bank;
   wire [3:0] U_dsdc_r_data_mask;
   wire [2088:2092] U_dsdc_n;
   wire [1:0] U_ddrwr_ddr_dqm;
   wire [15:0] U_ddrwr_ddr_wr_data;
   wire [1:0] U_ddrwr_i2_dqs;
   wire [31:24] U_cr_srefr;
   wire [15:11] U_addrdec_row_addr_mask;
   wire [5:0] U_dmc_data_cnt_nxt;

   BUF_X8 FE_PHC5253_U_cr_N551 (.Z(FE_PHN5253_U_cr_N551), 
	.A(FE_PHN1504_U_cr_N551));
   CLKBUF_X1 FE_PHC5237_U_cr_n455 (.Z(FE_PHN5237_U_cr_n455), 
	.A(U_cr_n455));
   BUF_X32 FE_PHC5234_U_cr_N551 (.Z(FE_PHN5234_U_cr_N551), 
	.A(FE_PHN5253_U_cr_N551));
   BUF_X1 FE_PHC5176_U_dsdc_n1637 (.Z(FE_PHN5176_U_dsdc_n1637), 
	.A(FE_PHN4625_U_dsdc_n1637));
   CLKBUF_X1 FE_PHC5174_U_dsdc_n1436 (.Z(FE_PHN5174_U_dsdc_n1436), 
	.A(FE_PHN4623_U_dsdc_n1436));
   CLKBUF_X1 FE_PHC5171_n27 (.Z(FE_PHN5171_n27), 
	.A(FE_PHN2432_n27));
   CLKBUF_X1 FE_PHC5144_U_dsdc_n226 (.Z(FE_PHN5144_U_dsdc_n226), 
	.A(U_dsdc_n226));
   CLKBUF_X1 FE_PHC5142_U_dsdc_n378 (.Z(FE_PHN5142_U_dsdc_n378), 
	.A(FE_PHN3165_U_dsdc_n378));
   CLKBUF_X1 FE_PHC5112_U_cr_N556 (.Z(FE_PHN5112_U_cr_N556), 
	.A(FE_PHN4204_U_cr_N556));
   BUF_X1 FE_PHC5110_U_cr_N398 (.Z(FE_PHN5110_U_cr_N398), 
	.A(U_cr_N398));
   CLKBUF_X1 FE_PHC5102_U_addrdec_N133 (.Z(FE_PHN5102_U_addrdec_N133), 
	.A(FE_PHN1594_U_addrdec_N133));
   CLKBUF_X1 FE_PHC5064_s_read_pipe_0_ (.Z(FE_PHN5064_s_read_pipe_0_), 
	.A(FE_PHN4152_s_read_pipe_0_));
   CLKBUF_X1 FE_PHC5056_U_dsdc_n376 (.Z(FE_PHN5056_U_dsdc_n376), 
	.A(FE_PHN3044_U_dsdc_n376));
   BUF_X1 FE_PHC5047_U_dsdc_n228 (.Z(FE_PHN5047_U_dsdc_n228), 
	.A(FE_PHN3234_U_dsdc_n228));
   CLKBUF_X1 FE_PHC5042_U_dsdc_N4228 (.Z(FE_PHN5042_U_dsdc_N4228), 
	.A(FE_PHN3183_U_dsdc_N4228));
   CLKBUF_X1 FE_PHC5012_U_dsdc_n371 (.Z(FE_PHN5012_U_dsdc_n371), 
	.A(FE_PHN3170_U_dsdc_n371));
   CLKBUF_X1 FE_PHC5011_U_cr_N559 (.Z(FE_PHN5011_U_cr_N559), 
	.A(FE_PHN3867_U_cr_N559));
   CLKBUF_X1 FE_PHC4966_U_cr_n65 (.Z(FE_PHN4966_U_cr_n65), 
	.A(FE_PHN3229_U_cr_n65));
   CLKBUF_X1 FE_PHC4962_U_dsdc_n230 (.Z(FE_PHN4962_U_dsdc_n230), 
	.A(FE_PHN3239_U_dsdc_n230));
   BUF_X1 FE_PHC4952_U_cr_n108 (.Z(FE_PHN4952_U_cr_n108), 
	.A(FE_PHN4013_U_cr_n108));
   CLKBUF_X1 FE_PHC4938_U_dmc_n12 (.Z(FE_PHN4938_U_dmc_n12), 
	.A(U_dmc_n12));
   CLKBUF_X1 FE_PHC4934_U_refctl_count_next_1_ (.Z(FE_PHN4934_U_refctl_count_next_1_), 
	.A(FE_PHN3305_U_refctl_count_next_1_));
   CLKBUF_X1 FE_PHC4922_U_cr_N564 (.Z(FE_PHN4922_U_cr_N564), 
	.A(U_cr_N564));
   CLKBUF_X1 FE_PHC4915_U_cr_n51 (.Z(FE_PHN4915_U_cr_n51), 
	.A(FE_PHN3968_U_cr_n51));
   CLKBUF_X1 FE_PHC4914_U_cr_n59 (.Z(FE_PHN4914_U_cr_n59), 
	.A(U_cr_n59));
   BUF_X1 FE_PHC4913_U_cr_N404 (.Z(FE_PHN4913_U_cr_N404), 
	.A(FE_PHN3479_U_cr_N404));
   CLKBUF_X1 FE_PHC4894_U_cr_n48 (.Z(FE_PHN4894_U_cr_n48), 
	.A(FE_PHN3938_U_cr_n48));
   CLKBUF_X1 FE_PHC4893_U_cr_N473 (.Z(FE_PHN4893_U_cr_N473), 
	.A(FE_PHN3816_U_cr_N473));
   CLKBUF_X1 FE_PHC4878_U_dsdc_n366 (.Z(FE_PHN4878_U_dsdc_n366), 
	.A(FE_PHN3167_U_dsdc_n366));
   BUF_X1 FE_PHC4871_U_cr_n46 (.Z(FE_PHN4871_U_cr_n46), 
	.A(FE_PHN4045_U_cr_n46));
   CLKBUF_X1 FE_PHC4855_U_cr_n49 (.Z(FE_PHN4855_U_cr_n49), 
	.A(FE_PHN4006_U_cr_n49));
   CLKBUF_X1 FE_PHC4851_U_cr_N691 (.Z(FE_PHN4851_U_cr_N691), 
	.A(FE_PHN3830_U_cr_N691));
   CLKBUF_X1 FE_PHC4849_U_cr_N395 (.Z(FE_PHN4849_U_cr_N395), 
	.A(U_cr_N395));
   CLKBUF_X1 FE_PHC4845_U_cr_n47 (.Z(FE_PHN4845_U_cr_n47), 
	.A(FE_PHN3889_U_cr_n47));
   CLKBUF_X1 FE_PHC4842_U_cr_N636 (.Z(FE_PHN4842_U_cr_N636), 
	.A(FE_PHN3810_U_cr_N636));
   CLKBUF_X1 FE_PHC4841_U_cr_N313 (.Z(FE_PHN4841_U_cr_N313), 
	.A(FE_PHN3223_U_cr_N313));
   CLKBUF_X1 FE_PHC4818_U_cr_N469 (.Z(FE_PHN4818_U_cr_N469), 
	.A(FE_PHN3786_U_cr_N469));
   CLKBUF_X1 FE_PHC4805_U_cr_N468 (.Z(FE_PHN4805_U_cr_N468), 
	.A(FE_PHN3781_U_cr_N468));
   CLKBUF_X1 FE_PHC4798_U_cr_n50 (.Z(FE_PHN4798_U_cr_n50), 
	.A(FE_PHN3876_U_cr_n50));
   CLKBUF_X1 FE_PHC4792_U_cr_N635 (.Z(FE_PHN4792_U_cr_N635), 
	.A(FE_PHN3771_U_cr_N635));
   CLKBUF_X1 FE_PHC4787_U_cr_N736 (.Z(FE_PHN4787_U_cr_N736), 
	.A(FE_PHN3776_U_cr_N736));
   CLKBUF_X1 FE_PHC4785_U_dsdc_N4229 (.Z(FE_PHN4785_U_dsdc_N4229), 
	.A(FE_PHN3288_U_dsdc_N4229));
   CLKBUF_X1 FE_PHC4777_U_dsdc_n214 (.Z(FE_PHN4777_U_dsdc_n214), 
	.A(FE_PHN2971_U_dsdc_n214));
   CLKBUF_X1 FE_PHC4776_U_cr_N558 (.Z(FE_PHN4776_U_cr_N558), 
	.A(FE_PHN3745_U_cr_N558));
   CLKBUF_X1 FE_PHC4775_U_cr_N476 (.Z(FE_PHN4775_U_cr_N476), 
	.A(FE_PHN3739_U_cr_N476));
   CLKBUF_X1 FE_PHC4763_U_cr_N479 (.Z(FE_PHN4763_U_cr_N479), 
	.A(FE_PHN3707_U_cr_N479));
   CLKBUF_X1 FE_PHC4760_U_cr_N397 (.Z(FE_PHN4760_U_cr_N397), 
	.A(FE_PHN3800_U_cr_N397));
   CLKBUF_X1 FE_PHC4759_U_cr_N745 (.Z(FE_PHN4759_U_cr_N745), 
	.A(FE_PHN3686_U_cr_N745));
   CLKBUF_X1 FE_PHC4736_U_cr_N403 (.Z(FE_PHN4736_U_cr_N403), 
	.A(FE_PHN3051_U_cr_N403));
   BUF_X32 FE_PHC4728_U_cr_N551 (.Z(FE_PHN4728_U_cr_N551), 
	.A(FE_PHN5234_U_cr_N551));
   CLKBUF_X2 FE_PHC4727_U_refctl_ref_req_next (.Z(FE_PHN4727_U_refctl_ref_req_next), 
	.A(FE_PHN3049_U_refctl_ref_req_next));
   CLKBUF_X1 FE_PHC4718_U_dsdc_n389 (.Z(FE_PHN4718_U_dsdc_n389), 
	.A(FE_PHN3298_U_dsdc_n389));
   CLKBUF_X1 FE_PHC4717_U_dsdc_n268 (.Z(FE_PHN4717_U_dsdc_n268), 
	.A(U_dsdc_n268));
   CLKBUF_X1 FE_PHC4716_U_dsdc_n261 (.Z(FE_PHN4716_U_dsdc_n261), 
	.A(U_dsdc_n261));
   CLKBUF_X1 FE_PHC4715_U_dsdc_n276 (.Z(FE_PHN4715_U_dsdc_n276), 
	.A(U_dsdc_n276));
   BUF_X1 FE_PHC4714_cr_t_xsr_1_ (.Z(FE_PHN4714_cr_t_xsr_1_), 
	.A(FE_PHN3292_cr_t_xsr_1_));
   CLKBUF_X1 FE_PHC4713_U_dmc_data_cnt_nxt_5_ (.Z(FE_PHN4713_U_dmc_data_cnt_nxt_5_), 
	.A(FE_PHN3291_U_dmc_data_cnt_nxt_5_));
   BUF_X1 FE_PHC4678_U_dsdc_N4428 (.Z(FE_PHN4678_U_dsdc_N4428), 
	.A(FE_PHN1097_U_dsdc_N4428));
   BUF_X1 FE_PHC4676_U_dsdc_N4381 (.Z(FE_PHN4676_U_dsdc_N4381), 
	.A(FE_PHN1096_U_dsdc_N4381));
   CLKBUF_X1 FE_PHC4645_U_cr_N302 (.Z(FE_PHN4645_U_cr_N302), 
	.A(FE_PHN3052_U_cr_N302));
   CLKBUF_X1 FE_PHC4627_U_cr_N405 (.Z(FE_PHN4627_U_cr_N405), 
	.A(FE_PHN2964_U_cr_N405));
   BUF_X8 FE_PHC4625_U_dsdc_n1637 (.Z(FE_PHN4625_U_dsdc_n1637), 
	.A(FE_PHN2910_U_dsdc_n1637));
   BUF_X8 FE_PHC4623_U_dsdc_n1436 (.Z(FE_PHN4623_U_dsdc_n1436), 
	.A(FE_PHN672_U_dsdc_n1436));
   BUF_X32 FE_PHC4620_U_cr_s_sda_d (.Z(FE_PHN4620_U_cr_s_sda_d), 
	.A(U_cr_s_sda_d));
   BUF_X32 FE_PHC4618_U_cr_n20 (.Z(FE_PHN4618_U_cr_n20), 
	.A(U_cr_n20));
   BUF_X32 FE_PHC4617_U_cr_n18 (.Z(FE_PHN4617_U_cr_n18), 
	.A(FE_PHN2051_U_cr_n18));
   CLKBUF_X1 FE_PHC4616_n27 (.Z(FE_PHN4616_n27), 
	.A(n27));
   CLKBUF_X1 FE_PHC4614_U_dsdc_n409 (.Z(FE_PHN4614_U_dsdc_n409), 
	.A(U_dsdc_n409));
   CLKBUF_X1 FE_PHC4613_U_dsdc_n386 (.Z(FE_PHN4613_U_dsdc_n386), 
	.A(U_dsdc_n386));
   CLKBUF_X1 FE_PHC4612_U_cr_n285 (.Z(FE_PHN4612_U_cr_n285), 
	.A(U_cr_n285));
   CLKBUF_X1 FE_PHC4610_U_dsdc_rcar_cnt1_nxt_0_ (.Z(FE_PHN4610_U_dsdc_rcar_cnt1_nxt_0_), 
	.A(U_dsdc_rcar_cnt1_nxt[0]));
   CLKBUF_X1 FE_PHC4609_U_cr_N301 (.Z(FE_PHN4609_U_cr_N301), 
	.A(U_cr_N301));
   CLKBUF_X1 FE_PHC4606_U_dsdc_N4347 (.Z(FE_PHN4606_U_dsdc_N4347), 
	.A(U_dsdc_N4347));
   CLKBUF_X1 FE_PHC4605_U_dsdc_N4339 (.Z(FE_PHN4605_U_dsdc_N4339), 
	.A(U_dsdc_N4339));
   CLKBUF_X1 FE_PHC4604_U_dsdc_N4341 (.Z(FE_PHN4604_U_dsdc_N4341), 
	.A(U_dsdc_N4341));
   CLKBUF_X1 FE_PHC4603_U_dsdc_n295 (.Z(FE_PHN4603_U_dsdc_n295), 
	.A(U_dsdc_n295));
   CLKBUF_X1 FE_PHC4600_U_dsdc_n393 (.Z(FE_PHN4600_U_dsdc_n393), 
	.A(U_dsdc_n393));
   CLKBUF_X1 FE_PHC4599_U_dsdc_n221 (.Z(FE_PHN4599_U_dsdc_n221), 
	.A(U_dsdc_n221));
   CLKBUF_X1 FE_PHC4598_U_dsdc_N4345 (.Z(FE_PHN4598_U_dsdc_N4345), 
	.A(U_dsdc_N4345));
   CLKBUF_X1 FE_PHC4594_U_cr_N409 (.Z(FE_PHN4594_U_cr_N409), 
	.A(U_cr_N409));
   CLKBUF_X1 FE_PHC4593_U_dsdc_N4337 (.Z(FE_PHN4593_U_dsdc_N4337), 
	.A(U_dsdc_N4337));
   CLKBUF_X1 FE_PHC4592_U_dsdc_n390 (.Z(FE_PHN4592_U_dsdc_n390), 
	.A(U_dsdc_n390));
   CLKBUF_X1 FE_PHC4591_U_dsdc_N4349 (.Z(FE_PHN4591_U_dsdc_N4349), 
	.A(U_dsdc_N4349));
   CLKBUF_X1 FE_PHC4589_U_cr_n286 (.Z(FE_PHN4589_U_cr_n286), 
	.A(U_cr_n286));
   CLKBUF_X1 FE_PHC4587_U_dsdc_N4140 (.Z(FE_PHN4587_U_dsdc_N4140), 
	.A(U_dsdc_N4140));
   CLKBUF_X1 FE_PHC4582_U_dsdc_n294 (.Z(FE_PHN4582_U_dsdc_n294), 
	.A(U_dsdc_n294));
   CLKBUF_X1 FE_PHC4581_U_dsdc_N4492 (.Z(FE_PHN4581_U_dsdc_N4492), 
	.A(U_dsdc_N4492));
   CLKBUF_X1 FE_PHC4578_U_dsdc_N4343 (.Z(FE_PHN4578_U_dsdc_N4343), 
	.A(U_dsdc_N4343));
   CLKBUF_X1 FE_PHC4574_U_cr_N563 (.Z(FE_PHN4574_U_cr_N563), 
	.A(U_cr_N563));
   CLKBUF_X1 FE_PHC4568_U_cr_N553 (.Z(FE_PHN4568_U_cr_N553), 
	.A(U_cr_N553));
   CLKBUF_X1 FE_PHC4558_U_dsdc_N4384 (.Z(FE_PHN4558_U_dsdc_N4384), 
	.A(U_dsdc_N4384));
   CLKBUF_X1 FE_PHC4551_U_dsdc_N4389 (.Z(FE_PHN4551_U_dsdc_N4389), 
	.A(U_dsdc_N4389));
   CLKBUF_X1 FE_PHC4547_U_dsdc_N4440 (.Z(FE_PHN4547_U_dsdc_N4440), 
	.A(U_dsdc_N4440));
   CLKBUF_X1 FE_PHC4546_U_dsdc_N4434 (.Z(FE_PHN4546_U_dsdc_N4434), 
	.A(U_dsdc_N4434));
   CLKBUF_X1 FE_PHC4543_U_refctl_count_next_0_ (.Z(FE_PHN4543_U_refctl_count_next_0_), 
	.A(U_refctl_count_next_0_));
   CLKBUF_X1 FE_PHC4542_U_dsdc_N4351 (.Z(FE_PHN4542_U_dsdc_N4351), 
	.A(U_dsdc_N4351));
   CLKBUF_X1 FE_PHC4537_U_dsdc_N4340 (.Z(FE_PHN4537_U_dsdc_N4340), 
	.A(U_dsdc_N4340));
   CLKBUF_X1 FE_PHC4530_U_dsdc_N4397 (.Z(FE_PHN4530_U_dsdc_N4397), 
	.A(U_dsdc_N4397));
   CLKBUF_X1 FE_PHC4528_U_dsdc_N4477 (.Z(FE_PHN4528_U_dsdc_N4477), 
	.A(U_dsdc_N4477));
   CLKBUF_X1 FE_PHC4527_U_dsdc_N4388 (.Z(FE_PHN4527_U_dsdc_N4388), 
	.A(U_dsdc_N4388));
   CLKBUF_X1 FE_PHC4522_U_dsdc_n300 (.Z(FE_PHN4522_U_dsdc_n300), 
	.A(U_dsdc_n300));
   CLKBUF_X1 FE_PHC4521_U_dsdc_N4436 (.Z(FE_PHN4521_U_dsdc_N4436), 
	.A(U_dsdc_N4436));
   CLKBUF_X1 FE_PHC4520_U_dsdc_N4433 (.Z(FE_PHN4520_U_dsdc_N4433), 
	.A(U_dsdc_N4433));
   CLKBUF_X1 FE_PHC4519_U_dsdc_N4336 (.Z(FE_PHN4519_U_dsdc_N4336), 
	.A(U_dsdc_N4336));
   CLKBUF_X1 FE_PHC4513_U_dsdc_N4383 (.Z(FE_PHN4513_U_dsdc_N4383), 
	.A(U_dsdc_N4383));
   CLKBUF_X1 FE_PHC4507_U_dsdc_N4444 (.Z(FE_PHN4507_U_dsdc_N4444), 
	.A(U_dsdc_N4444));
   CLKBUF_X1 FE_PHC4503_U_dsdc_N4473 (.Z(FE_PHN4503_U_dsdc_N4473), 
	.A(U_dsdc_N4473));
   CLKBUF_X1 FE_PHC4502_U_dsdc_N4442 (.Z(FE_PHN4502_U_dsdc_N4442), 
	.A(U_dsdc_N4442));
   CLKBUF_X1 FE_PHC4501_U_dsdc_N4431 (.Z(FE_PHN4501_U_dsdc_N4431), 
	.A(U_dsdc_N4431));
   CLKBUF_X1 FE_PHC4498_U_dsdc_N4481 (.Z(FE_PHN4498_U_dsdc_N4481), 
	.A(U_dsdc_N4481));
   CLKBUF_X1 FE_PHC4497_U_dsdc_wrapped_pop_flag_nxt (.Z(FE_PHN4497_U_dsdc_wrapped_pop_flag_nxt), 
	.A(U_dsdc_wrapped_pop_flag_nxt));
   CLKBUF_X1 FE_PHC4491_U_dsdc_N4491 (.Z(FE_PHN4491_U_dsdc_N4491), 
	.A(U_dsdc_N4491));
   CLKBUF_X1 FE_PHC4489_U_dsdc_N4430 (.Z(FE_PHN4489_U_dsdc_N4430), 
	.A(U_dsdc_N4430));
   CLKBUF_X1 FE_PHC4483_U_cr_N638 (.Z(FE_PHN4483_U_cr_N638), 
	.A(U_cr_N638));
   CLKBUF_X1 FE_PHC4480_U_dsdc_N4441 (.Z(FE_PHN4480_U_dsdc_N4441), 
	.A(U_dsdc_N4441));
   CLKBUF_X1 FE_PHC4473_U_dsdc_N4482 (.Z(FE_PHN4473_U_dsdc_N4482), 
	.A(U_dsdc_N4482));
   CLKBUF_X1 FE_PHC4470_U_cr_N646 (.Z(FE_PHN4470_U_cr_N646), 
	.A(U_cr_N646));
   CLKBUF_X1 FE_PHC4469_U_dsdc_N4439 (.Z(FE_PHN4469_U_dsdc_N4439), 
	.A(U_dsdc_N4439));
   CLKBUF_X1 FE_PHC4465_U_dsdc_N4488 (.Z(FE_PHN4465_U_dsdc_N4488), 
	.A(U_dsdc_N4488));
   CLKBUF_X1 FE_PHC4464_U_cr_n19 (.Z(FE_PHN4464_U_cr_n19), 
	.A(U_cr_n19));
   CLKBUF_X1 FE_PHC4461_U_dsdc_N4350 (.Z(FE_PHN4461_U_dsdc_N4350), 
	.A(U_dsdc_N4350));
   CLKBUF_X1 FE_PHC4455_U_dsdc_N4395 (.Z(FE_PHN4455_U_dsdc_N4395), 
	.A(U_dsdc_N4395));
   CLKBUF_X1 FE_PHC4445_U_dsdc_N4479 (.Z(FE_PHN4445_U_dsdc_N4479), 
	.A(U_dsdc_N4479));
   CLKBUF_X1 FE_PHC4443_U_dsdc_N4435 (.Z(FE_PHN4443_U_dsdc_N4435), 
	.A(U_dsdc_N4435));
   CLKBUF_X1 FE_PHC4442_U_dsdc_N4438 (.Z(FE_PHN4442_U_dsdc_N4438), 
	.A(U_dsdc_N4438));
   CLKBUF_X1 FE_PHC4435_U_dsdc_N4478 (.Z(FE_PHN4435_U_dsdc_N4478), 
	.A(U_dsdc_N4478));
   CLKBUF_X1 FE_PHC4434_U_dsdc_N4398 (.Z(FE_PHN4434_U_dsdc_N4398), 
	.A(U_dsdc_N4398));
   CLKBUF_X1 FE_PHC4429_U_cr_N644 (.Z(FE_PHN4429_U_cr_N644), 
	.A(U_cr_N644));
   CLKBUF_X1 FE_PHC4428_U_cr_N692 (.Z(FE_PHN4428_U_cr_N692), 
	.A(U_cr_N692));
   CLKBUF_X1 FE_PHC4424_U_dsdc_N4342 (.Z(FE_PHN4424_U_dsdc_N4342), 
	.A(U_dsdc_N4342));
   CLKBUF_X1 FE_PHC4423_U_dsdc_N4487 (.Z(FE_PHN4423_U_dsdc_N4487), 
	.A(U_dsdc_N4487));
   CLKBUF_X1 FE_PHC4415_U_dsdc_N4391 (.Z(FE_PHN4415_U_dsdc_N4391), 
	.A(U_dsdc_N4391));
   CLKBUF_X1 FE_PHC4414_U_dsdc_N4386 (.Z(FE_PHN4414_U_dsdc_N4386), 
	.A(U_dsdc_N4386));
   CLKBUF_X1 FE_PHC4410_U_refctl_count_next_4_ (.Z(FE_PHN4410_U_refctl_count_next_4_), 
	.A(U_refctl_count_next_4_));
   CLKBUF_X1 FE_PHC4409_U_cr_N305 (.Z(FE_PHN4409_U_cr_N305), 
	.A(U_cr_N305));
   CLKBUF_X1 FE_PHC4408_U_dsdc_N4390 (.Z(FE_PHN4408_U_dsdc_N4390), 
	.A(U_dsdc_N4390));
   CLKBUF_X1 FE_PHC4398_U_cr_N303 (.Z(FE_PHN4398_U_cr_N303), 
	.A(U_cr_N303));
   CLKBUF_X1 FE_PHC4397_U_dsdc_n279 (.Z(FE_PHN4397_U_dsdc_n279), 
	.A(U_dsdc_n279));
   CLKBUF_X1 FE_PHC4395_U_dsdc_wtr_cnt_nxt_0_ (.Z(FE_PHN4395_U_dsdc_wtr_cnt_nxt_0_), 
	.A(U_dsdc_wtr_cnt_nxt[0]));
   CLKBUF_X1 FE_PHC4391_U_dsdc_n209 (.Z(FE_PHN4391_U_dsdc_n209), 
	.A(U_dsdc_n209));
   CLKBUF_X1 FE_PHC4390_U_dsdc_N4483 (.Z(FE_PHN4390_U_dsdc_N4483), 
	.A(U_dsdc_N4483));
   CLKBUF_X1 FE_PHC4389_U_dsdc_N4392 (.Z(FE_PHN4389_U_dsdc_N4392), 
	.A(U_dsdc_N4392));
   CLKBUF_X1 FE_PHC4388_U_dsdc_N4394 (.Z(FE_PHN4388_U_dsdc_N4394), 
	.A(U_dsdc_N4394));
   CLKBUF_X1 FE_PHC4381_U_dsdc_N4489 (.Z(FE_PHN4381_U_dsdc_N4489), 
	.A(U_dsdc_N4489));
   CLKBUF_X1 FE_PHC4365_U_dsdc_N4485 (.Z(FE_PHN4365_U_dsdc_N4485), 
	.A(U_dsdc_N4485));
   CLKBUF_X1 FE_PHC4360_U_cr_N640 (.Z(FE_PHN4360_U_cr_N640), 
	.A(U_cr_N640));
   CLKBUF_X1 FE_PHC4359_U_dsdc_N4445 (.Z(FE_PHN4359_U_dsdc_N4445), 
	.A(U_dsdc_N4445));
   CLKBUF_X1 FE_PHC4354_U_dsdc_N4385 (.Z(FE_PHN4354_U_dsdc_N4385), 
	.A(U_dsdc_N4385));
   CLKBUF_X1 FE_PHC4353_U_dsdc_N4338 (.Z(FE_PHN4353_U_dsdc_N4338), 
	.A(U_dsdc_N4338));
   CLKBUF_X1 FE_PHC4349_U_dsdc_N4480 (.Z(FE_PHN4349_U_dsdc_N4480), 
	.A(U_dsdc_N4480));
   CLKBUF_X1 FE_PHC4345_U_dsdc_N4486 (.Z(FE_PHN4345_U_dsdc_N4486), 
	.A(U_dsdc_N4486));
   CLKBUF_X1 FE_PHC4344_U_dsdc_N4344 (.Z(FE_PHN4344_U_dsdc_N4344), 
	.A(U_dsdc_N4344));
   CLKBUF_X1 FE_PHC4342_U_dsdc_N4393 (.Z(FE_PHN4342_U_dsdc_N4393), 
	.A(U_dsdc_N4393));
   CLKBUF_X1 FE_PHC4339_U_dsdc_N4437 (.Z(FE_PHN4339_U_dsdc_N4437), 
	.A(U_dsdc_N4437));
   CLKBUF_X1 FE_PHC4328_U_dsdc_N4443 (.Z(FE_PHN4328_U_dsdc_N4443), 
	.A(U_dsdc_N4443));
   CLKBUF_X1 FE_PHC4323_U_dsdc_N4346 (.Z(FE_PHN4323_U_dsdc_N4346), 
	.A(U_dsdc_N4346));
   CLKBUF_X1 FE_PHC4315_U_dsdc_N4348 (.Z(FE_PHN4315_U_dsdc_N4348), 
	.A(U_dsdc_N4348));
   CLKBUF_X1 FE_PHC4308_U_dsdc_n213 (.Z(FE_PHN4308_U_dsdc_n213), 
	.A(U_dsdc_n213));
   CLKBUF_X1 FE_PHC4307_U_dsdc_N4396 (.Z(FE_PHN4307_U_dsdc_N4396), 
	.A(U_dsdc_N4396));
   CLKBUF_X1 FE_PHC4306_U_dsdc_N4490 (.Z(FE_PHN4306_U_dsdc_N4490), 
	.A(U_dsdc_N4490));
   CLKBUF_X1 FE_PHC4304_U_dsdc_N4484 (.Z(FE_PHN4304_U_dsdc_N4484), 
	.A(U_dsdc_N4484));
   CLKBUF_X1 FE_PHC4293_U_dsdc_n293 (.Z(FE_PHN4293_U_dsdc_n293), 
	.A(U_dsdc_n293));
   CLKBUF_X1 FE_PHC4286_U_dsdc_N4432 (.Z(FE_PHN4286_U_dsdc_N4432), 
	.A(U_dsdc_N4432));
   CLKBUF_X1 FE_PHC4277_U_dsdc_N4387 (.Z(FE_PHN4277_U_dsdc_N4387), 
	.A(U_dsdc_N4387));
   CLKBUF_X1 FE_PHC4265_U_cr_n29 (.Z(FE_PHN4265_U_cr_n29), 
	.A(U_cr_n29));
   CLKBUF_X1 FE_PHC4246_U_dsdc_n356 (.Z(FE_PHN4246_U_dsdc_n356), 
	.A(U_dsdc_n356));
   CLKBUF_X1 FE_PHC4204_U_cr_N556 (.Z(FE_PHN4204_U_cr_N556), 
	.A(U_cr_N556));
   CLKBUF_X1 FE_PHC4152_s_read_pipe_0_ (.Z(FE_PHN4152_s_read_pipe_0_), 
	.A(s_read_pipe[0]));
   BUF_X8 FE_PHC4110_U_cr_n53 (.Z(FE_PHN4110_U_cr_n53), 
	.A(U_cr_n53));
   BUF_X8 FE_PHC4075_U_dsdc_n185 (.Z(FE_PHN4075_U_dsdc_n185), 
	.A(U_dsdc_n185));
   CLKBUF_X1 FE_PHC4045_U_cr_n46 (.Z(FE_PHN4045_U_cr_n46), 
	.A(U_cr_n46));
   BUF_X8 FE_PHC4029_U_cr_N306 (.Z(FE_PHN4029_U_cr_N306), 
	.A(U_cr_N306));
   CLKBUF_X1 FE_PHC4013_U_cr_n108 (.Z(FE_PHN4013_U_cr_n108), 
	.A(U_cr_n108));
   CLKBUF_X1 FE_PHC4006_U_cr_n49 (.Z(FE_PHN4006_U_cr_n49), 
	.A(U_cr_n49));
   BUF_X8 FE_PHC3988_U_cr_n60 (.Z(FE_PHN3988_U_cr_n60), 
	.A(U_cr_n60));
   CLKBUF_X1 FE_PHC3968_U_cr_n51 (.Z(FE_PHN3968_U_cr_n51), 
	.A(U_cr_n51));
   BUF_X8 FE_PHC3951_U_dsdc_N4139 (.Z(FE_PHN3951_U_dsdc_N4139), 
	.A(U_dsdc_N4139));
   CLKBUF_X1 FE_PHC3938_U_cr_n48 (.Z(FE_PHN3938_U_cr_n48), 
	.A(U_cr_n48));
   CLKBUF_X1 FE_PHC3889_U_cr_n47 (.Z(FE_PHN3889_U_cr_n47), 
	.A(U_cr_n47));
   CLKBUF_X1 FE_PHC3876_U_cr_n50 (.Z(FE_PHN3876_U_cr_n50), 
	.A(U_cr_n50));
   BUF_X8 FE_PHC3870_U_dmc_n12 (.Z(FE_PHN3870_U_dmc_n12), 
	.A(FE_PHN4938_U_dmc_n12));
   BUF_X8 FE_PHC3867_U_cr_N559 (.Z(FE_PHN3867_U_cr_N559), 
	.A(U_cr_N559));
   BUF_X16 FE_PHC3844_U_cr_N472 (.Z(FE_PHN3844_U_cr_N472), 
	.A(U_cr_N472));
   BUF_X16 FE_PHC3833_U_cr_N642 (.Z(FE_PHN3833_U_cr_N642), 
	.A(U_cr_N642));
   BUF_X16 FE_PHC3831_U_cr_N696 (.Z(FE_PHN3831_U_cr_N696), 
	.A(U_cr_N696));
   BUF_X8 FE_PHC3830_U_cr_N691 (.Z(FE_PHN3830_U_cr_N691), 
	.A(U_cr_N691));
   BUF_X16 FE_PHC3826_U_cr_n83 (.Z(FE_PHN3826_U_cr_n83), 
	.A(U_cr_n83));
   BUF_X8 FE_PHC3816_U_cr_N473 (.Z(FE_PHN3816_U_cr_N473), 
	.A(U_cr_N473));
   BUF_X8 FE_PHC3810_U_cr_N636 (.Z(FE_PHN3810_U_cr_N636), 
	.A(U_cr_N636));
   BUF_X8 FE_PHC3800_U_cr_N397 (.Z(FE_PHN3800_U_cr_N397), 
	.A(U_cr_N397));
   BUF_X8 FE_PHC3786_U_cr_N469 (.Z(FE_PHN3786_U_cr_N469), 
	.A(U_cr_N469));
   BUF_X8 FE_PHC3781_U_cr_N468 (.Z(FE_PHN3781_U_cr_N468), 
	.A(U_cr_N468));
   BUF_X16 FE_PHC3777_U_cr_N697 (.Z(FE_PHN3777_U_cr_N697), 
	.A(U_cr_N697));
   BUF_X8 FE_PHC3776_U_cr_N736 (.Z(FE_PHN3776_U_cr_N736), 
	.A(U_cr_N736));
   BUF_X8 FE_PHC3771_U_cr_N635 (.Z(FE_PHN3771_U_cr_N635), 
	.A(U_cr_N635));
   BUF_X16 FE_PHC3768_U_cr_N637 (.Z(FE_PHN3768_U_cr_N637), 
	.A(U_cr_N637));
   BUF_X16 FE_PHC3766_U_cr_N402 (.Z(FE_PHN3766_U_cr_N402), 
	.A(U_cr_N402));
   BUF_X16 FE_PHC3760_U_cr_N471 (.Z(FE_PHN3760_U_cr_N471), 
	.A(U_cr_N471));
   BUF_X16 FE_PHC3759_U_cr_N394 (.Z(FE_PHN3759_U_cr_N394), 
	.A(U_cr_N394));
   BUF_X16 FE_PHC3758_U_cr_N560 (.Z(FE_PHN3758_U_cr_N560), 
	.A(U_cr_N560));
   BUF_X16 FE_PHC3757_U_cr_n82 (.Z(FE_PHN3757_U_cr_n82), 
	.A(U_cr_n82));
   BUF_X16 FE_PHC3751_U_cr_N478 (.Z(FE_PHN3751_U_cr_N478), 
	.A(U_cr_N478));
   BUF_X8 FE_PHC3745_U_cr_N558 (.Z(FE_PHN3745_U_cr_N558), 
	.A(U_cr_N558));
   BUF_X8 FE_PHC3739_U_cr_N476 (.Z(FE_PHN3739_U_cr_N476), 
	.A(U_cr_N476));
   BUF_X16 FE_PHC3738_U_cr_N474 (.Z(FE_PHN3738_U_cr_N474), 
	.A(U_cr_N474));
   BUF_X16 FE_PHC3737_U_cr_N737 (.Z(FE_PHN3737_U_cr_N737), 
	.A(U_cr_N737));
   BUF_X16 FE_PHC3736_U_cr_N645 (.Z(FE_PHN3736_U_cr_N645), 
	.A(U_cr_N645));
   BUF_X16 FE_PHC3724_U_cr_N396 (.Z(FE_PHN3724_U_cr_N396), 
	.A(U_cr_N396));
   BUF_X16 FE_PHC3722_U_cr_N699 (.Z(FE_PHN3722_U_cr_N699), 
	.A(U_cr_N699));
   BUF_X16 FE_PHC3714_U_cr_N694 (.Z(FE_PHN3714_U_cr_N694), 
	.A(U_cr_N694));
   BUF_X16 FE_PHC3713_U_cr_N299 (.Z(FE_PHN3713_U_cr_N299), 
	.A(U_cr_N299));
   BUF_X16 FE_PHC3712_U_cr_N555 (.Z(FE_PHN3712_U_cr_N555), 
	.A(U_cr_N555));
   BUF_X8 FE_PHC3707_U_cr_N479 (.Z(FE_PHN3707_U_cr_N479), 
	.A(U_cr_N479));
   BUF_X16 FE_PHC3704_U_cr_n90 (.Z(FE_PHN3704_U_cr_n90), 
	.A(U_cr_n90));
   BUF_X16 FE_PHC3702_U_cr_N695 (.Z(FE_PHN3702_U_cr_N695), 
	.A(U_cr_N695));
   BUF_X16 FE_PHC3698_U_cr_N740 (.Z(FE_PHN3698_U_cr_N740), 
	.A(U_cr_N740));
   BUF_X16 FE_PHC3697_U_cr_n89 (.Z(FE_PHN3697_U_cr_n89), 
	.A(U_cr_n89));
   BUF_X16 FE_PHC3692_U_cr_N298 (.Z(FE_PHN3692_U_cr_N298), 
	.A(U_cr_N298));
   BUF_X16 FE_PHC3687_U_cr_n91 (.Z(FE_PHN3687_U_cr_n91), 
	.A(U_cr_n91));
   BUF_X8 FE_PHC3686_U_cr_N745 (.Z(FE_PHN3686_U_cr_N745), 
	.A(U_cr_N745));
   BUF_X16 FE_PHC3684_U_cr_N643 (.Z(FE_PHN3684_U_cr_N643), 
	.A(U_cr_N643));
   BUF_X16 FE_PHC3683_U_cr_N310 (.Z(FE_PHN3683_U_cr_N310), 
	.A(U_cr_N310));
   BUF_X16 FE_PHC3680_U_cr_N693 (.Z(FE_PHN3680_U_cr_N693), 
	.A(U_cr_N693));
   BUF_X16 FE_PHC3672_U_cr_n88 (.Z(FE_PHN3672_U_cr_n88), 
	.A(U_cr_n88));
   BUF_X16 FE_PHC3669_U_cr_N477 (.Z(FE_PHN3669_U_cr_N477), 
	.A(U_cr_N477));
   BUF_X16 FE_PHC3666_U_cr_N700 (.Z(FE_PHN3666_U_cr_N700), 
	.A(U_cr_N700));
   BUF_X16 FE_PHC3665_U_cr_N470 (.Z(FE_PHN3665_U_cr_N470), 
	.A(U_cr_N470));
   BUF_X16 FE_PHC3660_U_cr_N647 (.Z(FE_PHN3660_U_cr_N647), 
	.A(U_cr_N647));
   BUF_X16 FE_PHC3659_U_cr_N639 (.Z(FE_PHN3659_U_cr_N639), 
	.A(U_cr_N639));
   BUF_X16 FE_PHC3657_U_cr_N698 (.Z(FE_PHN3657_U_cr_N698), 
	.A(U_cr_N698));
   BUF_X16 FE_PHC3651_U_cr_N554 (.Z(FE_PHN3651_U_cr_N554), 
	.A(U_cr_N554));
   BUF_X16 FE_PHC3645_U_cr_N738 (.Z(FE_PHN3645_U_cr_N738), 
	.A(U_cr_N738));
   BUF_X16 FE_PHC3643_U_cr_N641 (.Z(FE_PHN3643_U_cr_N641), 
	.A(U_cr_N641));
   BUF_X16 FE_PHC3640_U_cr_N475 (.Z(FE_PHN3640_U_cr_N475), 
	.A(U_cr_N475));
   BUF_X16 FE_PHC3638_U_cr_N739 (.Z(FE_PHN3638_U_cr_N739), 
	.A(U_cr_N739));
   BUF_X16 FE_PHC3628_U_cr_n92 (.Z(FE_PHN3628_U_cr_n92), 
	.A(U_cr_n92));
   BUF_X16 FE_PHC3619_U_cr_n94 (.Z(FE_PHN3619_U_cr_n94), 
	.A(U_cr_n94));
   BUF_X16 FE_PHC3614_U_cr_N550 (.Z(FE_PHN3614_U_cr_N550), 
	.A(U_cr_N550));
   BUF_X16 FE_PHC3613_U_dsdc_n405 (.Z(FE_PHN3613_U_dsdc_n405), 
	.A(U_dsdc_n405));
   BUF_X32 FE_PHC3607_U_refctl_count_next_2_ (.Z(FE_PHN3607_U_refctl_count_next_2_), 
	.A(FE_PHN1140_U_refctl_count_next_2_));
   BUF_X16 FE_PHC3600_U_cr_n59 (.Z(FE_PHN3600_U_cr_n59), 
	.A(FE_PHN4914_U_cr_n59));
   BUF_X16 FE_PHC3588_U_cr_n149 (.Z(FE_PHN3588_U_cr_n149), 
	.A(U_cr_n149));
   BUF_X32 FE_PHC3579_U_cr_N467 (.Z(FE_PHN3579_U_cr_N467), 
	.A(U_cr_N467));
   BUF_X32 FE_PHC3575_U_cr_N401 (.Z(FE_PHN3575_U_cr_N401), 
	.A(U_cr_N401));
   BUF_X32 FE_PHC3549_U_cr_n165 (.Z(FE_PHN3549_U_cr_n165), 
	.A(U_cr_n165));
   BUF_X32 FE_PHC3515_U_cr_N551 (.Z(FE_PHN3515_U_cr_N551), 
	.A(FE_PHN4728_U_cr_N551));
   CLKBUF_X1 FE_PHC3514_U_cr_n148 (.Z(FE_PHN3514_U_cr_n148), 
	.A(U_cr_n148));
   CLKBUF_X1 FE_PHC3513_U_dsdc_bm_ras_cnt_3__0_ (.Z(FE_PHN3513_U_dsdc_bm_ras_cnt_3__0_), 
	.A(U_dsdc_bm_ras_cnt_3__0_));
   CLKBUF_X1 FE_PHC3511_U_dsdc_bm_ras_cnt_0__0_ (.Z(FE_PHN3511_U_dsdc_bm_ras_cnt_0__0_), 
	.A(U_dsdc_bm_ras_cnt_0__0_));
   CLKBUF_X1 FE_PHC3510_U_dsdc_bm_ras_cnt_2__0_ (.Z(FE_PHN3510_U_dsdc_bm_ras_cnt_2__0_), 
	.A(U_dsdc_bm_ras_cnt_2__0_));
   CLKBUF_X1 FE_PHC3509_U_dsdc_bm_rc_cnt_2__0_ (.Z(FE_PHN3509_U_dsdc_bm_rc_cnt_2__0_), 
	.A(U_dsdc_bm_rc_cnt_2__0_));
   CLKBUF_X1 FE_PHC3508_U_dsdc_bm_rc_cnt_1__0_ (.Z(FE_PHN3508_U_dsdc_bm_rc_cnt_1__0_), 
	.A(U_dsdc_bm_rc_cnt_1__0_));
   CLKBUF_X1 FE_PHC3507_U_dsdc_bm_ras_cnt_1__0_ (.Z(FE_PHN3507_U_dsdc_bm_ras_cnt_1__0_), 
	.A(U_dsdc_bm_ras_cnt_1__0_));
   CLKBUF_X1 FE_PHC3505_U_cr_n45 (.Z(FE_PHN3505_U_cr_n45), 
	.A(U_cr_n45));
   CLKBUF_X1 FE_PHC3503_U_dsdc_rp_cnt1_nxt_0_ (.Z(FE_PHN3503_U_dsdc_rp_cnt1_nxt_0_), 
	.A(U_dsdc_rp_cnt1_nxt[0]));
   BUF_X8 FE_PHC3485_U_cr_n77 (.Z(FE_PHN3485_U_cr_n77), 
	.A(U_cr_n77));
   CLKBUF_X1 FE_PHC3480_U_cr_n80 (.Z(FE_PHN3480_U_cr_n80), 
	.A(U_cr_n80));
   CLKBUF_X1 FE_PHC3479_U_cr_N404 (.Z(FE_PHN3479_U_cr_N404), 
	.A(U_cr_N404));
   BUF_X16 FE_PHC3476_U_cr_n75 (.Z(FE_PHN3476_U_cr_n75), 
	.A(U_cr_n75));
   BUF_X32 FE_PHC3475_U_cr_n74 (.Z(FE_PHN3475_U_cr_n74), 
	.A(U_cr_n74));
   BUF_X32 FE_PHC3473_U_dsdc_n2095 (.Z(FE_PHN3473_U_dsdc_n2095), 
	.A(FE_PHN772_U_dsdc_n2095));
   CLKBUF_X1 FE_PHC3467_U_dsdc_n1924 (.Z(FE_PHN3467_U_dsdc_n1924), 
	.A(U_dsdc_n1924));
   CLKBUF_X1 FE_PHC3464_U_dsdc_n319 (.Z(FE_PHN3464_U_dsdc_n319), 
	.A(U_dsdc_n319));
   BUF_X1 FE_PHC3463_U_dsdc_n1594 (.Z(FE_PHN3463_U_dsdc_n1594), 
	.A(U_dsdc_n1594));
   BUF_X1 FE_PHC3461_U_dsdc_n394 (.Z(FE_PHN3461_U_dsdc_n394), 
	.A(U_dsdc_n394));
   CLKBUF_X1 FE_PHC3456_U_cr_N690 (.Z(FE_PHN3456_U_cr_N690), 
	.A(U_cr_N690));
   CLKBUF_X1 FE_PHC3454_U_dmc_n40 (.Z(FE_PHN3454_U_dmc_n40), 
	.A(U_dmc_n40));
   CLKBUF_X1 FE_PHC3452_U_dsdc_n410 (.Z(FE_PHN3452_U_dsdc_n410), 
	.A(U_dsdc_n410));
   CLKBUF_X1 FE_PHC3450_U_dsdc_wtr_cnt_nxt_1_ (.Z(FE_PHN3450_U_dsdc_wtr_cnt_nxt_1_), 
	.A(U_dsdc_wtr_cnt_nxt[1]));
   CLKBUF_X1 FE_PHC3449_U_refctl_next_state_0_ (.Z(FE_PHN3449_U_refctl_next_state_0_), 
	.A(U_refctl_next_state_0_));
   CLKBUF_X1 FE_PHC3446_U_dsdc_n269 (.Z(FE_PHN3446_U_dsdc_n269), 
	.A(U_dsdc_n269));
   CLKBUF_X1 FE_PHC3445_U_dsdc_n391 (.Z(FE_PHN3445_U_dsdc_n391), 
	.A(U_dsdc_n391));
   CLKBUF_X1 FE_PHC3443_U_dsdc_n282 (.Z(FE_PHN3443_U_dsdc_n282), 
	.A(U_dsdc_n282));
   CLKBUF_X1 FE_PHC3442_U_dsdc_n240 (.Z(FE_PHN3442_U_dsdc_n240), 
	.A(U_dsdc_n240));
   CLKBUF_X1 FE_PHC3440_U_dsdc_n265 (.Z(FE_PHN3440_U_dsdc_n265), 
	.A(U_dsdc_n265));
   CLKBUF_X1 FE_PHC3432_U_dsdc_n296 (.Z(FE_PHN3432_U_dsdc_n296), 
	.A(U_dsdc_n296));
   CLKBUF_X1 FE_PHC3431_U_dsdc_n256 (.Z(FE_PHN3431_U_dsdc_n256), 
	.A(U_dsdc_n256));
   CLKBUF_X1 FE_PHC3427_U_dsdc_rp_cnt2_nxt_2_ (.Z(FE_PHN3427_U_dsdc_rp_cnt2_nxt_2_), 
	.A(U_dsdc_rp_cnt2_nxt[2]));
   CLKBUF_X1 FE_PHC3415_U_dsdc_n266 (.Z(FE_PHN3415_U_dsdc_n266), 
	.A(U_dsdc_n266));
   CLKBUF_X1 FE_PHC3407_U_dsdc_n267 (.Z(FE_PHN3407_U_dsdc_n267), 
	.A(U_dsdc_n267));
   CLKBUF_X1 FE_PHC3399_U_dsdc_n412 (.Z(FE_PHN3399_U_dsdc_n412), 
	.A(U_dsdc_n412));
   CLKBUF_X1 FE_PHC3389_U_cr_N734 (.Z(FE_PHN3389_U_cr_N734), 
	.A(U_cr_N734));
   CLKBUF_X1 FE_PHC3379_U_cr_N733 (.Z(FE_PHN3379_U_cr_N733), 
	.A(U_cr_N733));
   CLKBUF_X1 FE_PHC3378_U_cr_N735 (.Z(FE_PHN3378_U_cr_N735), 
	.A(U_cr_N735));
   CLKBUF_X1 FE_PHC3373_U_addrdec_n347 (.Z(FE_PHN3373_U_addrdec_n347), 
	.A(FE_PHN2427_U_addrdec_n347));
   CLKBUF_X1 FE_PHC3371_U_dsdc_n1231 (.Z(FE_PHN3371_U_dsdc_n1231), 
	.A(U_dsdc_n1231));
   CLKBUF_X1 FE_PHC3370_U_dsdc_n271 (.Z(FE_PHN3370_U_dsdc_n271), 
	.A(U_dsdc_n271));
   CLKBUF_X1 FE_PHC3355_U_dsdc_n406 (.Z(FE_PHN3355_U_dsdc_n406), 
	.A(U_dsdc_n406));
   CLKBUF_X1 FE_PHC3352_U_cr_n87 (.Z(FE_PHN3352_U_cr_n87), 
	.A(U_cr_n87));
   CLKBUF_X1 FE_PHC3349_U_cr_n86 (.Z(FE_PHN3349_U_cr_n86), 
	.A(U_cr_n86));
   CLKBUF_X1 FE_PHC3346_U_dsdc_n277 (.Z(FE_PHN3346_U_dsdc_n277), 
	.A(U_dsdc_n277));
   CLKBUF_X1 FE_PHC3345_U_dmc_n13 (.Z(FE_PHN3345_U_dmc_n13), 
	.A(FE_PHN866_U_dmc_n13));
   CLKBUF_X1 FE_PHC3343_U_refctl_count_next_3_ (.Z(FE_PHN3343_U_refctl_count_next_3_), 
	.A(U_refctl_count_next_3_));
   CLKBUF_X1 FE_PHC3337_U_dsdc_N4429 (.Z(FE_PHN3337_U_dsdc_N4429), 
	.A(U_dsdc_N4429));
   CLKBUF_X1 FE_PHC3328_U_dsdc_N4476 (.Z(FE_PHN3328_U_dsdc_N4476), 
	.A(U_dsdc_N4476));
   CLKBUF_X1 FE_PHC3327_U_dsdc_wr_cnt_nxt_0_ (.Z(FE_PHN3327_U_dsdc_wr_cnt_nxt_0_), 
	.A(U_dsdc_wr_cnt_nxt[0]));
   CLKBUF_X1 FE_PHC3326_U_refctl_count_next_15_ (.Z(FE_PHN3326_U_refctl_count_next_15_), 
	.A(U_refctl_count_next_15_));
   CLKBUF_X1 FE_PHC3325_U_dsdc_n262 (.Z(FE_PHN3325_U_dsdc_n262), 
	.A(U_dsdc_n262));
   CLKBUF_X1 FE_PHC3324_U_dsdc_num_init_ref_cnt_nxt_1_ (.Z(FE_PHN3324_U_dsdc_num_init_ref_cnt_nxt_1_), 
	.A(U_dsdc_num_init_ref_cnt_nxt[1]));
   CLKBUF_X1 FE_PHC3322_U_dsdc_n270 (.Z(FE_PHN3322_U_dsdc_n270), 
	.A(U_dsdc_n270));
   CLKBUF_X1 FE_PHC3321_U_dsdc_n263 (.Z(FE_PHN3321_U_dsdc_n263), 
	.A(U_dsdc_n263));
   CLKBUF_X1 FE_PHC3320_U_dsdc_n222 (.Z(FE_PHN3320_U_dsdc_n222), 
	.A(U_dsdc_n222));
   CLKBUF_X1 FE_PHC3319_U_dsdc_n255 (.Z(FE_PHN3319_U_dsdc_n255), 
	.A(U_dsdc_n255));
   CLKBUF_X1 FE_PHC3318_U_dsdc_n264 (.Z(FE_PHN3318_U_dsdc_n264), 
	.A(U_dsdc_n264));
   CLKBUF_X1 FE_PHC3317_U_dsdc_n259 (.Z(FE_PHN3317_U_dsdc_n259), 
	.A(U_dsdc_n259));
   CLKBUF_X1 FE_PHC3316_U_dsdc_n260 (.Z(FE_PHN3316_U_dsdc_n260), 
	.A(U_dsdc_n260));
   CLKBUF_X1 FE_PHC3315_U_dsdc_n211 (.Z(FE_PHN3315_U_dsdc_n211), 
	.A(U_dsdc_n211));
   CLKBUF_X1 FE_PHC3314_U_dsdc_n261 (.Z(FE_PHN3314_U_dsdc_n261), 
	.A(FE_PHN4716_U_dsdc_n261));
   CLKBUF_X1 FE_PHC3313_U_dsdc_rp_cnt1_0_ (.Z(FE_PHN3313_U_dsdc_rp_cnt1_0_), 
	.A(U_dsdc_rp_cnt1_0_));
   CLKBUF_X1 FE_PHC3312_U_dsdc_n257 (.Z(FE_PHN3312_U_dsdc_n257), 
	.A(U_dsdc_n257));
   CLKBUF_X1 FE_PHC3311_U_dsdc_n268 (.Z(FE_PHN3311_U_dsdc_n268), 
	.A(FE_PHN4717_U_dsdc_n268));
   BUF_X8 FE_PHC3309_U_dsdc_cas_latency_cnt_2_ (.Z(FE_PHN3309_U_dsdc_cas_latency_cnt_2_), 
	.A(U_dsdc_cas_latency_cnt_2_));
   CLKBUF_X1 FE_PHC3305_U_refctl_count_next_1_ (.Z(FE_PHN3305_U_refctl_count_next_1_), 
	.A(U_refctl_count_next_1_));
   BUF_X8 FE_PHC3299_U_dsdc_n274 (.Z(FE_PHN3299_U_dsdc_n274), 
	.A(U_dsdc_n274));
   BUF_X8 FE_PHC3298_U_dsdc_n389 (.Z(FE_PHN3298_U_dsdc_n389), 
	.A(U_dsdc_n389));
   BUF_X8 FE_PHC3297_U_dsdc_n283 (.Z(FE_PHN3297_U_dsdc_n283), 
	.A(U_dsdc_n283));
   BUF_X8 FE_PHC3293_U_dsdc_n276 (.Z(FE_PHN3293_U_dsdc_n276), 
	.A(FE_PHN4715_U_dsdc_n276));
   BUF_X8 FE_PHC3292_cr_t_xsr_1_ (.Z(FE_PHN3292_cr_t_xsr_1_), 
	.A(cr_t_xsr[1]));
   BUF_X8 FE_PHC3291_U_dmc_data_cnt_nxt_5_ (.Z(FE_PHN3291_U_dmc_data_cnt_nxt_5_), 
	.A(FE_PHN1211_U_dmc_data_cnt_nxt_5_));
   BUF_X16 FE_PHC3289_U_dsdc_n275 (.Z(FE_PHN3289_U_dsdc_n275), 
	.A(U_dsdc_n275));
   BUF_X8 FE_PHC3288_U_dsdc_N4229 (.Z(FE_PHN3288_U_dsdc_N4229), 
	.A(U_dsdc_N4229));
   BUF_X16 FE_PHC3287_U_cr_N576 (.Z(FE_PHN3287_U_cr_N576), 
	.A(FE_PHN1640_U_cr_N576));
   BUF_X16 FE_PHC3286_U_cr_n85 (.Z(FE_PHN3286_U_cr_n85), 
	.A(U_cr_n85));
   BUF_X16 FE_PHC3283_cr_reg_data_out_24_ (.Z(FE_PHN3283_cr_reg_data_out_24_), 
	.A(cr_reg_data_out[24]));
   CLKBUF_X1 FE_PHC3268_U_dsdc_init_cnt_10_ (.Z(FE_PHN3268_U_dsdc_init_cnt_10_), 
	.A(U_dsdc_init_cnt_10_));
   CLKBUF_X1 FE_PHC3260_U_dsdc_n1212 (.Z(FE_PHN3260_U_dsdc_n1212), 
	.A(U_dsdc_n1212));
   CLKBUF_X1 FE_PHC3259_U_dsdc_n1205 (.Z(FE_PHN3259_U_dsdc_n1205), 
	.A(U_dsdc_n1205));
   CLKBUF_X1 FE_PHC3258_U_dsdc_n1184 (.Z(FE_PHN3258_U_dsdc_n1184), 
	.A(U_dsdc_n1184));
   CLKBUF_X1 FE_PHC3256_U_dsdc_n1198 (.Z(FE_PHN3256_U_dsdc_n1198), 
	.A(U_dsdc_n1198));
   CLKBUF_X1 FE_PHC3255_U_dsdc_n1241 (.Z(FE_PHN3255_U_dsdc_n1241), 
	.A(U_dsdc_n1241));
   CLKBUF_X1 FE_PHC3252_U_dsdc_n1191 (.Z(FE_PHN3252_U_dsdc_n1191), 
	.A(U_dsdc_n1191));
   CLKBUF_X1 FE_PHC3250_U_cr_N311 (.Z(FE_PHN3250_U_cr_N311), 
	.A(U_cr_N311));
   CLKBUF_X1 FE_PHC3249_U_cr_N312 (.Z(FE_PHN3249_U_cr_N312), 
	.A(U_cr_N312));
   CLKBUF_X1 FE_PHC3247_U_dsdc_n1177 (.Z(FE_PHN3247_U_dsdc_n1177), 
	.A(U_dsdc_n1177));
   CLKBUF_X1 FE_PHC3245_U_dsdc_N4462 (.Z(FE_PHN3245_U_dsdc_N4462), 
	.A(FE_PHN1059_U_dsdc_N4462));
   CLKBUF_X1 FE_PHC3244_U_dsdc_n227 (.Z(FE_PHN3244_U_dsdc_n227), 
	.A(U_dsdc_n227));
   CLKBUF_X1 FE_PHC3242_U_dsdc_N4332 (.Z(FE_PHN3242_U_dsdc_N4332), 
	.A(U_dsdc_N4332));
   CLKBUF_X1 FE_PHC3241_U_dsdc_n212 (.Z(FE_PHN3241_U_dsdc_n212), 
	.A(U_dsdc_n212));
   CLKBUF_X1 FE_PHC3240_cr_t_rcar_2_ (.Z(FE_PHN3240_cr_t_rcar_2_), 
	.A(cr_t_rcar[2]));
   CLKBUF_X1 FE_PHC3239_U_dsdc_n230 (.Z(FE_PHN3239_U_dsdc_n230), 
	.A(U_dsdc_n230));
   CLKBUF_X1 FE_PHC3238_U_dsdc_rp_cnt1_nxt_1_ (.Z(FE_PHN3238_U_dsdc_rp_cnt1_nxt_1_), 
	.A(U_dsdc_rp_cnt1_nxt[1]));
   CLKBUF_X1 FE_PHC3237_U_cr_N562 (.Z(FE_PHN3237_U_cr_N562), 
	.A(U_cr_N562));
   CLKBUF_X1 FE_PHC3235_U_dsdc_n201 (.Z(FE_PHN3235_U_dsdc_n201), 
	.A(U_dsdc_n201));
   BUF_X8 FE_PHC3234_U_dsdc_n228 (.Z(FE_PHN3234_U_dsdc_n228), 
	.A(U_dsdc_n228));
   BUF_X8 FE_PHC3233_U_dsdc_n377 (.Z(FE_PHN3233_U_dsdc_n377), 
	.A(U_dsdc_n377));
   BUF_X8 FE_PHC3232_U_dsdc_n370 (.Z(FE_PHN3232_U_dsdc_n370), 
	.A(U_dsdc_n370));
   BUF_X8 FE_PHC3231_U_dsdc_n379 (.Z(FE_PHN3231_U_dsdc_n379), 
	.A(U_dsdc_n379));
   CLKBUF_X1 FE_PHC3230_U_cr_n81 (.Z(FE_PHN3230_U_cr_n81), 
	.A(U_cr_n81));
   BUF_X8 FE_PHC3229_U_cr_n65 (.Z(FE_PHN3229_U_cr_n65), 
	.A(U_cr_n65));
   BUF_X8 FE_PHC3228_U_dsdc_n368 (.Z(FE_PHN3228_U_dsdc_n368), 
	.A(U_dsdc_n368));
   BUF_X8 FE_PHC3227_U_dsdc_n372 (.Z(FE_PHN3227_U_dsdc_n372), 
	.A(U_dsdc_n372));
   BUF_X16 FE_PHC3224_U_cr_N410 (.Z(FE_PHN3224_U_cr_N410), 
	.A(U_cr_N410));
   BUF_X8 FE_PHC3223_U_cr_N313 (.Z(FE_PHN3223_U_cr_N313), 
	.A(U_cr_N313));
   BUF_X16 FE_PHC3222_U_dsdc_n375 (.Z(FE_PHN3222_U_dsdc_n375), 
	.A(U_dsdc_n375));
   BUF_X8 FE_PHC3221_U_dsdc_n381 (.Z(FE_PHN3221_U_dsdc_n381), 
	.A(U_dsdc_n381));
   BUF_X16 FE_PHC3220_U_cr_N408 (.Z(FE_PHN3220_U_cr_N408), 
	.A(FE_PHN1524_U_cr_N408));
   BUF_X16 FE_PHC3216_U_dsdc_n373 (.Z(FE_PHN3216_U_dsdc_n373), 
	.A(U_dsdc_n373));
   BUF_X16 FE_PHC3215_U_cr_n76 (.Z(FE_PHN3215_U_cr_n76), 
	.A(U_cr_n76));
   BUF_X32 FE_PHC3212_U_cr_n93 (.Z(FE_PHN3212_U_cr_n93), 
	.A(U_cr_n93));
   BUF_X32 FE_PHC3208_U_dsdc_n2096 (.Z(FE_PHN3208_U_dsdc_n2096), 
	.A(U_dsdc_n2096));
   CLKBUF_X1 FE_PHC3197_U_dmc_n59 (.Z(FE_PHN3197_U_dmc_n59), 
	.A(U_dmc_n59));
   CLKBUF_X1 FE_PHC3196_U_cr_n99 (.Z(FE_PHN3196_U_cr_n99), 
	.A(U_cr_n99));
   CLKBUF_X1 FE_PHC3195_U_dsdc_n417 (.Z(FE_PHN3195_U_dsdc_n417), 
	.A(U_dsdc_n417));
   CLKBUF_X1 FE_PHC3194_U_dsdc_cas_cnt_nxt_3_ (.Z(FE_PHN3194_U_dsdc_cas_cnt_nxt_3_), 
	.A(U_dsdc_cas_cnt_nxt[3]));
   CLKBUF_X1 FE_PHC3193_U_dmc_n1 (.Z(FE_PHN3193_U_dmc_n1), 
	.A(FE_PHN1597_U_dmc_n1));
   CLKBUF_X1 FE_PHC3192_U_cr_n128 (.Z(FE_PHN3192_U_cr_n128), 
	.A(U_cr_n128));
   CLKBUF_X1 FE_PHC3191_U_dsdc_n388 (.Z(FE_PHN3191_U_dsdc_n388), 
	.A(U_dsdc_n388));
   CLKBUF_X1 FE_PHC3189_U_dsdc_N4334 (.Z(FE_PHN3189_U_dsdc_N4334), 
	.A(FE_PHN1098_U_dsdc_N4334));
   CLKBUF_X1 FE_PHC3188_U_addrdec_N119 (.Z(FE_PHN3188_U_addrdec_N119), 
	.A(U_addrdec_N119));
   CLKBUF_X1 FE_PHC3187_U_dsdc_rcar_cnt1_nxt_3_ (.Z(FE_PHN3187_U_dsdc_rcar_cnt1_nxt_3_), 
	.A(U_dsdc_rcar_cnt1_nxt[3]));
   CLKBUF_X1 FE_PHC3186_U_dsdc_num_init_ref_cnt_nxt_0_ (.Z(FE_PHN3186_U_dsdc_num_init_ref_cnt_nxt_0_), 
	.A(U_dsdc_num_init_ref_cnt_nxt[0]));
   CLKBUF_X1 FE_PHC3185_U_cr_n73 (.Z(FE_PHN3185_U_cr_n73), 
	.A(U_cr_n73));
   CLKBUF_X1 FE_PHC3183_U_dsdc_N4228 (.Z(FE_PHN3183_U_dsdc_N4228), 
	.A(U_dsdc_N4228));
   CLKBUF_X1 FE_PHC3182_U_dsdc_N4368 (.Z(FE_PHN3182_U_dsdc_N4368), 
	.A(FE_PHN1055_U_dsdc_N4368));
   BUF_X8 FE_PHC3170_U_dsdc_n371 (.Z(FE_PHN3170_U_dsdc_n371), 
	.A(U_dsdc_n371));
   BUF_X16 FE_PHC3169_U_dsdc_n367 (.Z(FE_PHN3169_U_dsdc_n367), 
	.A(U_dsdc_n367));
   BUF_X16 FE_PHC3168_U_dsdc_n380 (.Z(FE_PHN3168_U_dsdc_n380), 
	.A(U_dsdc_n380));
   BUF_X8 FE_PHC3167_U_dsdc_n366 (.Z(FE_PHN3167_U_dsdc_n366), 
	.A(U_dsdc_n366));
   BUF_X16 FE_PHC3166_U_dsdc_n374 (.Z(FE_PHN3166_U_dsdc_n374), 
	.A(U_dsdc_n374));
   BUF_X8 FE_PHC3165_U_dsdc_n378 (.Z(FE_PHN3165_U_dsdc_n378), 
	.A(U_dsdc_n378));
   CLKBUF_X1 FE_PHC3164_U_addrdec_N130 (.Z(FE_PHN3164_U_addrdec_N130), 
	.A(U_addrdec_N130));
   BUF_X16 FE_PHC3162_U_dsdc_n369 (.Z(FE_PHN3162_U_dsdc_n369), 
	.A(U_dsdc_n369));
   BUF_X32 FE_PHC3160_U_dsdc_n423 (.Z(FE_PHN3160_U_dsdc_n423), 
	.A(U_dsdc_n423));
   BUF_X32 FE_PHC3156_U_dsdc_n281 (.Z(FE_PHN3156_U_dsdc_n281), 
	.A(U_dsdc_n281));
   CLKBUF_X1 FE_PHC3127_U_dsdc_n414 (.Z(FE_PHN3127_U_dsdc_n414), 
	.A(FE_PHN1029_U_dsdc_n414));
   CLKBUF_X1 FE_PHC3126_cr_block_size1_6_ (.Z(FE_PHN3126_cr_block_size1_6_), 
	.A(cr_block_size1[6]));
   CLKBUF_X1 FE_PHC3123_U_dsdc_n407 (.Z(FE_PHN3123_U_dsdc_n407), 
	.A(FE_PHN1220_U_dsdc_n407));
   CLKBUF_X1 FE_PHC3119_U_dsdc_n411 (.Z(FE_PHN3119_U_dsdc_n411), 
	.A(FE_PHN1214_U_dsdc_n411));
   CLKBUF_X1 FE_PHC3115_U_dsdc_n297 (.Z(FE_PHN3115_U_dsdc_n297), 
	.A(U_dsdc_n297));
   CLKBUF_X1 FE_PHC3113_U_cr_n63 (.Z(FE_PHN3113_U_cr_n63), 
	.A(U_cr_n63));
   CLKBUF_X1 FE_PHC3112_U_dsdc_n415 (.Z(FE_PHN3112_U_dsdc_n415), 
	.A(FE_PHN968_U_dsdc_n415));
   CLKBUF_X1 FE_PHC3111_cr_s_data_width_early_0_ (.Z(FE_PHN3111_cr_s_data_width_early_0_), 
	.A(cr_s_data_width_early_0_));
   CLKBUF_X1 FE_PHC3110_U_dsdc_num_init_ref_cnt_nxt_2_ (.Z(FE_PHN3110_U_dsdc_num_init_ref_cnt_nxt_2_), 
	.A(U_dsdc_num_init_ref_cnt_nxt[2]));
   CLKBUF_X1 FE_PHC3109_U_dsdc_N4415 (.Z(FE_PHN3109_U_dsdc_N4415), 
	.A(FE_PHN1057_U_dsdc_N4415));
   CLKBUF_X1 FE_PHC3108_U_dsdc_N4321 (.Z(FE_PHN3108_U_dsdc_N4321), 
	.A(FE_PHN1060_U_dsdc_N4321));
   CLKBUF_X1 FE_PHC3107_U_cr_n44 (.Z(FE_PHN3107_U_cr_n44), 
	.A(U_cr_n44));
   BUF_X16 FE_PHC3106_U_cr_n43 (.Z(FE_PHN3106_U_cr_n43), 
	.A(U_cr_n43));
   BUF_X16 FE_PHC3105_U_dsdc_n_2090_ (.Z(FE_PHN3105_U_dsdc_n_2090_), 
	.A(FE_PHN934_U_dsdc_n_2090_));
   BUF_X16 FE_PHC3104_U_dsdc_N4174 (.Z(FE_PHN3104_U_dsdc_N4174), 
	.A(U_dsdc_N4174));
   CLKBUF_X1 FE_PHC3087_U_dsdc_cas_cnt_nxt_2_ (.Z(FE_PHN3087_U_dsdc_cas_cnt_nxt_2_), 
	.A(U_dsdc_cas_cnt_nxt[2]));
   CLKBUF_X1 FE_PHC3086_U_dsdc_n1275 (.Z(FE_PHN3086_U_dsdc_n1275), 
	.A(U_dsdc_n1275));
   CLKBUF_X1 FE_PHC3085_U_dsdc_rp_cnt2_nxt_0_ (.Z(FE_PHN3085_U_dsdc_rp_cnt2_nxt_0_), 
	.A(U_dsdc_rp_cnt2_nxt[0]));
   CLKBUF_X1 FE_PHC3083_U_dsdc_n280 (.Z(FE_PHN3083_U_dsdc_n280), 
	.A(U_dsdc_n280));
   CLKBUF_X1 FE_PHC3082_U_dsdc_n418 (.Z(FE_PHN3082_U_dsdc_n418), 
	.A(U_dsdc_n418));
   CLKBUF_X1 FE_PHC3081_U_dsdc_n416 (.Z(FE_PHN3081_U_dsdc_n416), 
	.A(FE_PHN966_U_dsdc_n416));
   CLKBUF_X1 FE_PHC3080_U_dsdc_n431 (.Z(FE_PHN3080_U_dsdc_n431), 
	.A(U_dsdc_n431));
   CLKBUF_X1 FE_PHC3079_U_dsdc_rcar_cnt2_nxt_3_ (.Z(FE_PHN3079_U_dsdc_rcar_cnt2_nxt_3_), 
	.A(U_dsdc_rcar_cnt2_nxt[3]));
   CLKBUF_X1 FE_PHC3077_U_dsdc_n460 (.Z(FE_PHN3077_U_dsdc_n460), 
	.A(U_dsdc_n460));
   CLKBUF_X1 FE_PHC3075_cr_push_n (.Z(FE_PHN3075_cr_push_n), 
	.A(cr_push_n));
   CLKBUF_X2 FE_PHC3054_cr_row_addr_width_2_ (.Z(FE_PHN3054_cr_row_addr_width_2_), 
	.A(cr_row_addr_width[2]));
   BUF_X16 FE_PHC3053_U_dsdc_n231 (.Z(FE_PHN3053_U_dsdc_n231), 
	.A(FE_PHN961_U_dsdc_n231));
   CLKBUF_X1 FE_PHC3052_U_cr_N302 (.Z(FE_PHN3052_U_cr_N302), 
	.A(U_cr_N302));
   CLKBUF_X1 FE_PHC3051_U_cr_N403 (.Z(FE_PHN3051_U_cr_N403), 
	.A(U_cr_N403));
   BUF_X16 FE_PHC3049_U_refctl_ref_req_next (.Z(FE_PHN3049_U_refctl_ref_req_next), 
	.A(FE_PHN1251_U_refctl_ref_req_next));
   CLKBUF_X1 FE_PHC3047_U_dsdc_wr_cnt_nxt_2_ (.Z(FE_PHN3047_U_dsdc_wr_cnt_nxt_2_), 
	.A(U_dsdc_wr_cnt_nxt[2]));
   CLKBUF_X1 FE_PHC3046_ctl_sd_in_sf_mode (.Z(FE_PHN3046_ctl_sd_in_sf_mode), 
	.A(FE_PHN1224_ctl_sd_in_sf_mode));
   CLKBUF_X1 FE_PHC3045_U_dsdc_rp_cnt1_nxt_2_ (.Z(FE_PHN3045_U_dsdc_rp_cnt1_nxt_2_), 
	.A(U_dsdc_rp_cnt1_nxt[2]));
   BUF_X8 FE_PHC3044_U_dsdc_n376 (.Z(FE_PHN3044_U_dsdc_n376), 
	.A(U_dsdc_n376));
   BUF_X32 FE_PHC3043_U_cr_N413 (.Z(FE_PHN3043_U_cr_N413), 
	.A(U_cr_N413));
   CLKBUF_X1 FE_PHC3041_cr_t_init_0_ (.Z(FE_PHN3041_cr_t_init_0_), 
	.A(cr_t_init[0]));
   CLKBUF_X1 FE_PHC3034_U_dsdc_N4381 (.Z(FE_PHN3034_U_dsdc_N4381), 
	.A(FE_PHN4676_U_dsdc_N4381));
   CLKBUF_X1 FE_PHC3033_U_dsdc_N4428 (.Z(FE_PHN3033_U_dsdc_N4428), 
	.A(FE_PHN4678_U_dsdc_N4428));
   BUF_X32 FE_PHC3031_n4 (.Z(FE_PHN3031_n4), 
	.A(n4));
   BUF_X32 FE_PHC3030_n6 (.Z(FE_PHN3030_n6), 
	.A(n6));
   BUF_X32 FE_PHC3029_n5 (.Z(FE_PHN3029_n5), 
	.A(n5));
   BUF_X32 FE_PHC3028_U_dsdc_term_cnt_nxt_4_ (.Z(FE_PHN3028_U_dsdc_term_cnt_nxt_4_), 
	.A(U_dsdc_term_cnt_nxt[4]));
   BUF_X8 FE_PHC3013_U_dsdc_N4475 (.Z(FE_PHN3013_U_dsdc_N4475), 
	.A(FE_PHN1061_U_dsdc_N4475));
   CLKBUF_X1 FE_PHC3012_U_cr_n147 (.Z(FE_PHN3012_U_cr_n147), 
	.A(U_cr_n147));
   BUF_X32 FE_PHC3011_U_dsdc_term_cnt_nxt_2_ (.Z(FE_PHN3011_U_dsdc_term_cnt_nxt_2_), 
	.A(U_dsdc_term_cnt_nxt[2]));
   CLKBUF_X1 FE_PHC2978_U_dsdc_N4141 (.Z(FE_PHN2978_U_dsdc_N4141), 
	.A(FE_PHN1058_U_dsdc_N4141));
   BUF_X32 FE_PHC2977_U_cr_N315 (.Z(FE_PHN2977_U_cr_N315), 
	.A(FE_PHN932_U_cr_N315));
   BUF_X32 FE_PHC2975_U_dsdc_n216 (.Z(FE_PHN2975_U_dsdc_n216), 
	.A(U_dsdc_n216));
   BUF_X8 FE_PHC2971_U_dsdc_n214 (.Z(FE_PHN2971_U_dsdc_n214), 
	.A(U_dsdc_n214));
   CLKBUF_X1 FE_PHC2964_U_cr_N405 (.Z(FE_PHN2964_U_cr_N405), 
	.A(U_cr_N405));
   BUF_X32 FE_PHC2941_U_dsdc_term_cnt_nxt_0_ (.Z(FE_PHN2941_U_dsdc_term_cnt_nxt_0_), 
	.A(U_dsdc_term_cnt_nxt[0]));
   BUF_X32 FE_PHC2929_cr_reg_data_out_15_ (.Z(FE_PHN2929_cr_reg_data_out_15_), 
	.A(FE_PHN694_cr_reg_data_out_15_));
   BUF_X32 FE_PHC2915_U_cr_N566 (.Z(FE_PHN2915_U_cr_N566), 
	.A(U_cr_N566));
   BUF_X32 FE_PHC2910_U_dsdc_n1637 (.Z(FE_PHN2910_U_dsdc_n1637), 
	.A(U_dsdc_n1637));
   CLKBUF_X1 FE_PHC2909_U_dsdc_n1436 (.Z(FE_PHN2909_U_dsdc_n1436), 
	.A(FE_PHN5174_U_dsdc_n1436));
   BUF_X32 FE_PHC2905_U_cr_s_sda_d (.Z(FE_PHN2905_U_cr_s_sda_d), 
	.A(FE_PHN4620_U_cr_s_sda_d));
   BUF_X32 FE_PHC2455_U_cr_n20 (.Z(FE_PHN2455_U_cr_n20), 
	.A(FE_PHN4618_U_cr_n20));
   BUF_X32 FE_PHC2432_n27 (.Z(FE_PHN2432_n27), 
	.A(FE_PHN4616_n27));
   CLKBUF_X1 FE_PHC2431_U_addrdec_N129 (.Z(FE_PHN2431_U_addrdec_N129), 
	.A(U_addrdec_N129));
   BUF_X8 FE_PHC2427_U_addrdec_n347 (.Z(FE_PHN2427_U_addrdec_n347), 
	.A(U_addrdec_n347));
   BUF_X32 FE_PHC2425_U_dsdc_N4341 (.Z(FE_PHN2425_U_dsdc_N4341), 
	.A(FE_PHN4604_U_dsdc_N4341));
   BUF_X32 FE_PHC2424_U_dsdc_N4347 (.Z(FE_PHN2424_U_dsdc_N4347), 
	.A(FE_PHN4606_U_dsdc_N4347));
   BUF_X32 FE_PHC2423_U_dsdc_N4345 (.Z(FE_PHN2423_U_dsdc_N4345), 
	.A(FE_PHN4598_U_dsdc_N4345));
   BUF_X32 FE_PHC2422_U_addrdec_n348 (.Z(FE_PHN2422_U_addrdec_n348), 
	.A(U_addrdec_n348));
   BUF_X32 FE_PHC2419_U_dsdc_N4343 (.Z(FE_PHN2419_U_dsdc_N4343), 
	.A(FE_PHN4578_U_dsdc_N4343));
   BUF_X32 FE_PHC2418_U_dsdc_N4440 (.Z(FE_PHN2418_U_dsdc_N4440), 
	.A(FE_PHN4547_U_dsdc_N4440));
   BUF_X32 FE_PHC2417_U_dsdc_N4477 (.Z(FE_PHN2417_U_dsdc_N4477), 
	.A(FE_PHN4528_U_dsdc_N4477));
   BUF_X32 FE_PHC2416_U_dsdc_N4492 (.Z(FE_PHN2416_U_dsdc_N4492), 
	.A(FE_PHN4581_U_dsdc_N4492));
   BUF_X32 FE_PHC2414_U_dsdc_N4389 (.Z(FE_PHN2414_U_dsdc_N4389), 
	.A(FE_PHN4551_U_dsdc_N4389));
   BUF_X32 FE_PHC2413_U_dsdc_N4397 (.Z(FE_PHN2413_U_dsdc_N4397), 
	.A(FE_PHN4530_U_dsdc_N4397));
   BUF_X32 FE_PHC2411_U_dsdc_N4430 (.Z(FE_PHN2411_U_dsdc_N4430), 
	.A(FE_PHN4489_U_dsdc_N4430));
   BUF_X32 FE_PHC2410_U_dsdc_N4336 (.Z(FE_PHN2410_U_dsdc_N4336), 
	.A(FE_PHN4519_U_dsdc_N4336));
   BUF_X32 FE_PHC2409_U_dsdc_N4491 (.Z(FE_PHN2409_U_dsdc_N4491), 
	.A(FE_PHN4491_U_dsdc_N4491));
   BUF_X32 FE_PHC2408_U_dsdc_N4351 (.Z(FE_PHN2408_U_dsdc_N4351), 
	.A(FE_PHN4542_U_dsdc_N4351));
   BUF_X32 FE_PHC2407_U_dsdc_N4433 (.Z(FE_PHN2407_U_dsdc_N4433), 
	.A(FE_PHN4520_U_dsdc_N4433));
   BUF_X32 FE_PHC2406_U_dsdc_N4444 (.Z(FE_PHN2406_U_dsdc_N4444), 
	.A(FE_PHN4507_U_dsdc_N4444));
   BUF_X32 FE_PHC2405_U_dsdc_N4438 (.Z(FE_PHN2405_U_dsdc_N4438), 
	.A(FE_PHN4442_U_dsdc_N4438));
   BUF_X32 FE_PHC2404_U_dsdc_N4388 (.Z(FE_PHN2404_U_dsdc_N4388), 
	.A(FE_PHN4527_U_dsdc_N4388));
   BUF_X32 FE_PHC2402_U_dsdc_N4483 (.Z(FE_PHN2402_U_dsdc_N4483), 
	.A(FE_PHN4390_U_dsdc_N4483));
   BUF_X32 FE_PHC2401_U_dsdc_N4342 (.Z(FE_PHN2401_U_dsdc_N4342), 
	.A(FE_PHN4424_U_dsdc_N4342));
   BUF_X32 FE_PHC2400_U_dsdc_N4488 (.Z(FE_PHN2400_U_dsdc_N4488), 
	.A(FE_PHN4465_U_dsdc_N4488));
   BUF_X32 FE_PHC2399_U_dsdc_N4384 (.Z(FE_PHN2399_U_dsdc_N4384), 
	.A(FE_PHN4558_U_dsdc_N4384));
   BUF_X32 FE_PHC2398_U_dsdc_N4391 (.Z(FE_PHN2398_U_dsdc_N4391), 
	.A(FE_PHN4415_U_dsdc_N4391));
   BUF_X32 FE_PHC2397_U_dsdc_N4480 (.Z(FE_PHN2397_U_dsdc_N4480), 
	.A(FE_PHN4349_U_dsdc_N4480));
   BUF_X32 FE_PHC2396_U_dsdc_N4386 (.Z(FE_PHN2396_U_dsdc_N4386), 
	.A(FE_PHN4414_U_dsdc_N4386));
   BUF_X32 FE_PHC2395_U_dsdc_N4395 (.Z(FE_PHN2395_U_dsdc_N4395), 
	.A(FE_PHN4455_U_dsdc_N4395));
   BUF_X32 FE_PHC2394_U_dsdc_N4390 (.Z(FE_PHN2394_U_dsdc_N4390), 
	.A(FE_PHN4408_U_dsdc_N4390));
   BUF_X32 FE_PHC2393_U_dsdc_N4478 (.Z(FE_PHN2393_U_dsdc_N4478), 
	.A(FE_PHN4435_U_dsdc_N4478));
   BUF_X32 FE_PHC2392_U_dsdc_N4392 (.Z(FE_PHN2392_U_dsdc_N4392), 
	.A(FE_PHN4389_U_dsdc_N4392));
   BUF_X32 FE_PHC2391_U_dsdc_N4385 (.Z(FE_PHN2391_U_dsdc_N4385), 
	.A(FE_PHN4354_U_dsdc_N4385));
   BUF_X32 FE_PHC2390_U_dsdc_N4437 (.Z(FE_PHN2390_U_dsdc_N4437), 
	.A(FE_PHN4339_U_dsdc_N4437));
   BUF_X32 FE_PHC2389_U_dsdc_N4432 (.Z(FE_PHN2389_U_dsdc_N4432), 
	.A(FE_PHN4286_U_dsdc_N4432));
   BUF_X32 FE_PHC2388_U_dsdc_N4338 (.Z(FE_PHN2388_U_dsdc_N4338), 
	.A(FE_PHN4353_U_dsdc_N4338));
   BUF_X32 FE_PHC2387_U_dsdc_N4486 (.Z(FE_PHN2387_U_dsdc_N4486), 
	.A(FE_PHN4345_U_dsdc_N4486));
   BUF_X32 FE_PHC2386_U_dsdc_N4396 (.Z(FE_PHN2386_U_dsdc_N4396), 
	.A(FE_PHN4307_U_dsdc_N4396));
   BUF_X32 FE_PHC2384_U_dsdc_N4393 (.Z(FE_PHN2384_U_dsdc_N4393), 
	.A(FE_PHN4342_U_dsdc_N4393));
   BUF_X32 FE_PHC2383_U_dsdc_N4443 (.Z(FE_PHN2383_U_dsdc_N4443), 
	.A(FE_PHN4328_U_dsdc_N4443));
   BUF_X32 FE_PHC2382_U_dsdc_N4344 (.Z(FE_PHN2382_U_dsdc_N4344), 
	.A(FE_PHN4344_U_dsdc_N4344));
   BUF_X32 FE_PHC2381_U_dsdc_N4348 (.Z(FE_PHN2381_U_dsdc_N4348), 
	.A(FE_PHN4315_U_dsdc_N4348));
   BUF_X32 FE_PHC2380_U_dsdc_N4490 (.Z(FE_PHN2380_U_dsdc_N4490), 
	.A(FE_PHN4306_U_dsdc_N4490));
   BUF_X32 FE_PHC2377_U_dsdc_N4366 (.Z(FE_PHN2377_U_dsdc_N4366), 
	.A(U_dsdc_N4366));
   BUF_X32 FE_PHC2373_U_dsdc_N4387 (.Z(FE_PHN2373_U_dsdc_N4387), 
	.A(FE_PHN4277_U_dsdc_N4387));
   BUF_X16 FE_PHC2146_U_addrdec_N131 (.Z(FE_PHN2146_U_addrdec_N131), 
	.A(U_addrdec_N131));
   BUF_X32 FE_PHC2051_U_cr_n18 (.Z(FE_PHN2051_U_cr_n18), 
	.A(U_cr_n18));
   BUF_X32 FE_PHC2044_U_dsdc_n273 (.Z(FE_PHN2044_U_dsdc_n273), 
	.A(U_dsdc_n273));
   BUF_X32 FE_PHC2040_U_dsdc_n271 (.Z(FE_PHN2040_U_dsdc_n271), 
	.A(FE_PHN3370_U_dsdc_n271));
   BUF_X32 FE_PHC2038_U_dsdc_n277 (.Z(FE_PHN2038_U_dsdc_n277), 
	.A(FE_PHN3346_U_dsdc_n277));
   BUF_X32 FE_PHC2037_U_dsdc_rcar_cnt1_nxt_0_ (.Z(FE_PHN2037_U_dsdc_rcar_cnt1_nxt_0_), 
	.A(FE_PHN4610_U_dsdc_rcar_cnt1_nxt_0_));
   BUF_X32 FE_PHC2036_U_dsdc_cas_latency_cnt_0_ (.Z(FE_PHN2036_U_dsdc_cas_latency_cnt_0_), 
	.A(U_dsdc_cas_latency_cnt_0_));
   BUF_X32 FE_PHC2034_U_dsdc_bm_ras_cnt_max_0_ (.Z(FE_PHN2034_U_dsdc_bm_ras_cnt_max_0_), 
	.A(U_dsdc_bm_ras_cnt_max_0_));
   BUF_X32 FE_PHC2033_U_dsdc_n262 (.Z(FE_PHN2033_U_dsdc_n262), 
	.A(FE_PHN3325_U_dsdc_n262));
   BUF_X32 FE_PHC2032_U_dsdc_n270 (.Z(FE_PHN2032_U_dsdc_n270), 
	.A(FE_PHN3322_U_dsdc_n270));
   BUF_X32 FE_PHC2031_U_dsdc_n264 (.Z(FE_PHN2031_U_dsdc_n264), 
	.A(FE_PHN3318_U_dsdc_n264));
   BUF_X32 FE_PHC2030_U_dsdc_n255 (.Z(FE_PHN2030_U_dsdc_n255), 
	.A(FE_PHN3319_U_dsdc_n255));
   BUF_X32 FE_PHC2029_U_dsdc_n263 (.Z(FE_PHN2029_U_dsdc_n263), 
	.A(FE_PHN3321_U_dsdc_n263));
   BUF_X32 FE_PHC2027_U_dsdc_n268 (.Z(FE_PHN2027_U_dsdc_n268), 
	.A(FE_PHN3311_U_dsdc_n268));
   BUF_X32 FE_PHC2025_U_addrdec_N107 (.Z(FE_PHN2025_U_addrdec_N107), 
	.A(U_addrdec_N107));
   BUF_X32 FE_PHC1921_U_dsdc_n1084 (.Z(FE_PHN1921_U_dsdc_n1084), 
	.A(U_dsdc_n1084));
   BUF_X32 FE_PHC1918_U_cr_n285 (.Z(FE_PHN1918_U_cr_n285), 
	.A(FE_PHN4612_U_cr_n285));
   BUF_X32 FE_PHC1917_U_cr_N304 (.Z(FE_PHN1917_U_cr_N304), 
	.A(U_cr_N304));
   BUF_X32 FE_PHC1916_U_cr_N556 (.Z(FE_PHN1916_U_cr_N556), 
	.A(FE_PHN5112_U_cr_N556));
   BUF_X32 FE_PHC1913_U_cr_N389 (.Z(FE_PHN1913_U_cr_N389), 
	.A(U_cr_N389));
   BUF_X32 FE_PHC1911_U_cr_N399 (.Z(FE_PHN1911_U_cr_N399), 
	.A(U_cr_N399));
   BUF_X16 FE_PHC1897_U_dsdc_n1002 (.Z(FE_PHN1897_U_dsdc_n1002), 
	.A(U_dsdc_n1002));
   BUF_X32 FE_PHC1896_U_dsdc_r_burst_size_1_ (.Z(FE_PHN1896_U_dsdc_r_burst_size_1_), 
	.A(U_dsdc_r_burst_size_1_));
   BUF_X32 FE_PHC1895_U_dsdc_n996 (.Z(FE_PHN1895_U_dsdc_n996), 
	.A(U_dsdc_n996));
   BUF_X32 FE_PHC1893_U_dsdc_n1392 (.Z(FE_PHN1893_U_dsdc_n1392), 
	.A(U_dsdc_n1392));
   CLKBUF_X1 FE_PHC1892_U_dsdc_r_burst_size_3_ (.Z(FE_PHN1892_U_dsdc_r_burst_size_3_), 
	.A(U_dsdc_r_burst_size_3_));
   BUF_X32 FE_PHC1891_U_dsdc_bm_ras_cnt_3__2_ (.Z(FE_PHN1891_U_dsdc_bm_ras_cnt_3__2_), 
	.A(U_dsdc_bm_ras_cnt_3__2_));
   CLKBUF_X1 FE_PHC1890_U_dsdc_r_burst_size_5_ (.Z(FE_PHN1890_U_dsdc_r_burst_size_5_), 
	.A(U_dsdc_r_burst_size_5_));
   BUF_X32 FE_PHC1889_U_dsdc_bm_ras_cnt_1__2_ (.Z(FE_PHN1889_U_dsdc_bm_ras_cnt_1__2_), 
	.A(U_dsdc_bm_ras_cnt_1__2_));
   CLKBUF_X1 FE_PHC1888_U_dsdc_r_burst_size_4_ (.Z(FE_PHN1888_U_dsdc_r_burst_size_4_), 
	.A(U_dsdc_r_burst_size_4_));
   CLKBUF_X1 FE_PHC1887_U_dsdc_n166 (.Z(FE_PHN1887_U_dsdc_n166), 
	.A(U_dsdc_n166));
   BUF_X32 FE_PHC1868_U_addrdec_n309 (.Z(FE_PHN1868_U_addrdec_n309), 
	.A(U_addrdec_n309));
   BUF_X32 FE_PHC1855_cr_block_size1_7_ (.Z(FE_PHN1855_cr_block_size1_7_), 
	.A(cr_block_size1[7]));
   BUF_X32 FE_PHC1854_U_addrdec_n346 (.Z(FE_PHN1854_U_addrdec_n346), 
	.A(U_addrdec_n346));
   BUF_X32 FE_PHC1848_U_cr_N464 (.Z(FE_PHN1848_U_cr_N464), 
	.A(U_cr_N464));
   BUF_X32 FE_PHC1845_U_cr_N465 (.Z(FE_PHN1845_U_cr_N465), 
	.A(U_cr_N465));
   BUF_X32 FE_PHC1747_U_cr_N555 (.Z(FE_PHN1747_U_cr_N555), 
	.A(FE_PHN3712_U_cr_N555));
   BUF_X32 FE_PHC1746_U_cr_N554 (.Z(FE_PHN1746_U_cr_N554), 
	.A(FE_PHN3651_U_cr_N554));
   BUF_X32 FE_PHC1745_U_cr_N557 (.Z(FE_PHN1745_U_cr_N557), 
	.A(U_cr_N557));
   BUF_X32 FE_PHC1740_U_cr_N564 (.Z(FE_PHN1740_U_cr_N564), 
	.A(FE_PHN4922_U_cr_N564));
   BUF_X32 FE_PHC1739_U_cr_N392 (.Z(FE_PHN1739_U_cr_N392), 
	.A(U_cr_N392));
   BUF_X32 FE_PHC1738_U_cr_N402 (.Z(FE_PHN1738_U_cr_N402), 
	.A(FE_PHN3766_U_cr_N402));
   BUF_X32 FE_PHC1737_U_cr_N390 (.Z(FE_PHN1737_U_cr_N390), 
	.A(U_cr_N390));
   BUF_X32 FE_PHC1736_U_cr_N394 (.Z(FE_PHN1736_U_cr_N394), 
	.A(FE_PHN3759_U_cr_N394));
   BUF_X32 FE_PHC1735_U_cr_N395 (.Z(FE_PHN1735_U_cr_N395), 
	.A(FE_PHN4849_U_cr_N395));
   BUF_X32 FE_PHC1734_U_cr_N396 (.Z(FE_PHN1734_U_cr_N396), 
	.A(FE_PHN3724_U_cr_N396));
   BUF_X32 FE_PHC1733_U_cr_N563 (.Z(FE_PHN1733_U_cr_N563), 
	.A(FE_PHN4574_U_cr_N563));
   BUF_X32 FE_PHC1732_U_cr_N479 (.Z(FE_PHN1732_U_cr_N479), 
	.A(FE_PHN4763_U_cr_N479));
   BUF_X32 FE_PHC1731_U_cr_N560 (.Z(FE_PHN1731_U_cr_N560), 
	.A(FE_PHN3758_U_cr_N560));
   BUF_X32 FE_PHC1730_U_cr_N472 (.Z(FE_PHN1730_U_cr_N472), 
	.A(FE_PHN3844_U_cr_N472));
   BUF_X32 FE_PHC1729_U_cr_N397 (.Z(FE_PHN1729_U_cr_N397), 
	.A(FE_PHN4760_U_cr_N397));
   BUF_X32 FE_PHC1728_U_cr_N475 (.Z(FE_PHN1728_U_cr_N475), 
	.A(FE_PHN3640_U_cr_N475));
   BUF_X32 FE_PHC1727_U_cr_N473 (.Z(FE_PHN1727_U_cr_N473), 
	.A(FE_PHN4893_U_cr_N473));
   BUF_X32 FE_PHC1726_U_cr_N558 (.Z(FE_PHN1726_U_cr_N558), 
	.A(FE_PHN4776_U_cr_N558));
   BUF_X32 FE_PHC1725_U_cr_N400 (.Z(FE_PHN1725_U_cr_N400), 
	.A(U_cr_N400));
   BUF_X32 FE_PHC1724_U_cr_N398 (.Z(FE_PHN1724_U_cr_N398), 
	.A(FE_PHN5110_U_cr_N398));
   BUF_X32 FE_PHC1723_U_cr_N644 (.Z(FE_PHN1723_U_cr_N644), 
	.A(FE_PHN4429_U_cr_N644));
   BUF_X32 FE_PHC1722_U_cr_N647 (.Z(FE_PHN1722_U_cr_N647), 
	.A(FE_PHN3660_U_cr_N647));
   BUF_X32 FE_PHC1721_U_cr_N641 (.Z(FE_PHN1721_U_cr_N641), 
	.A(FE_PHN3643_U_cr_N641));
   BUF_X32 FE_PHC1720_U_cr_N643 (.Z(FE_PHN1720_U_cr_N643), 
	.A(FE_PHN3684_U_cr_N643));
   BUF_X32 FE_PHC1719_U_cr_N476 (.Z(FE_PHN1719_U_cr_N476), 
	.A(FE_PHN4775_U_cr_N476));
   BUF_X32 FE_PHC1718_U_cr_N640 (.Z(FE_PHN1718_U_cr_N640), 
	.A(FE_PHN4360_U_cr_N640));
   BUF_X32 FE_PHC1716_U_cr_n82 (.Z(FE_PHN1716_U_cr_n82), 
	.A(FE_PHN3757_U_cr_n82));
   BUF_X32 FE_PHC1715_U_cr_N642 (.Z(FE_PHN1715_U_cr_N642), 
	.A(FE_PHN3833_U_cr_N642));
   BUF_X32 FE_PHC1714_U_cr_N635 (.Z(FE_PHN1714_U_cr_N635), 
	.A(FE_PHN4792_U_cr_N635));
   BUF_X32 FE_PHC1713_U_cr_N636 (.Z(FE_PHN1713_U_cr_N636), 
	.A(FE_PHN4842_U_cr_N636));
   BUF_X32 FE_PHC1712_U_cr_N738 (.Z(FE_PHN1712_U_cr_N738), 
	.A(FE_PHN3645_U_cr_N738));
   BUF_X32 FE_PHC1711_U_cr_N471 (.Z(FE_PHN1711_U_cr_N471), 
	.A(FE_PHN3760_U_cr_N471));
   BUF_X32 FE_PHC1710_U_cr_n83 (.Z(FE_PHN1710_U_cr_n83), 
	.A(FE_PHN3826_U_cr_n83));
   BUF_X32 FE_PHC1709_U_cr_N739 (.Z(FE_PHN1709_U_cr_N739), 
	.A(FE_PHN3638_U_cr_N739));
   BUF_X32 FE_PHC1708_U_cr_N468 (.Z(FE_PHN1708_U_cr_N468), 
	.A(FE_PHN4805_U_cr_N468));
   BUF_X32 FE_PHC1707_U_cr_N740 (.Z(FE_PHN1707_U_cr_N740), 
	.A(FE_PHN3698_U_cr_N740));
   BUF_X32 FE_PHC1706_U_cr_N301 (.Z(FE_PHN1706_U_cr_N301), 
	.A(FE_PHN4609_U_cr_N301));
   BUF_X32 FE_PHC1705_U_cr_N470 (.Z(FE_PHN1705_U_cr_N470), 
	.A(FE_PHN3665_U_cr_N470));
   BUF_X32 FE_PHC1704_U_cr_N469 (.Z(FE_PHN1704_U_cr_N469), 
	.A(FE_PHN4818_U_cr_N469));
   BUF_X32 FE_PHC1703_U_cr_N691 (.Z(FE_PHN1703_U_cr_N691), 
	.A(FE_PHN4851_U_cr_N691));
   BUF_X32 FE_PHC1702_U_cr_N693 (.Z(FE_PHN1702_U_cr_N693), 
	.A(FE_PHN3680_U_cr_N693));
   BUF_X32 FE_PHC1701_U_cr_N737 (.Z(FE_PHN1701_U_cr_N737), 
	.A(FE_PHN3737_U_cr_N737));
   BUF_X32 FE_PHC1700_U_cr_N300 (.Z(FE_PHN1700_U_cr_N300), 
	.A(U_cr_N300));
   BUF_X32 FE_PHC1699_U_cr_N299 (.Z(FE_PHN1699_U_cr_N299), 
	.A(FE_PHN3713_U_cr_N299));
   BUF_X32 FE_PHC1698_U_cr_N696 (.Z(FE_PHN1698_U_cr_N696), 
	.A(FE_PHN3831_U_cr_N696));
   BUF_X32 FE_PHC1697_U_cr_N697 (.Z(FE_PHN1697_U_cr_N697), 
	.A(FE_PHN3777_U_cr_N697));
   BUF_X32 FE_PHC1696_U_cr_N698 (.Z(FE_PHN1696_U_cr_N698), 
	.A(FE_PHN3657_U_cr_N698));
   BUF_X32 FE_PHC1695_U_cr_N700 (.Z(FE_PHN1695_U_cr_N700), 
	.A(FE_PHN3666_U_cr_N700));
   BUF_X32 FE_PHC1694_U_cr_n89 (.Z(FE_PHN1694_U_cr_n89), 
	.A(FE_PHN3697_U_cr_n89));
   BUF_X32 FE_PHC1693_U_cr_n91 (.Z(FE_PHN1693_U_cr_n91), 
	.A(FE_PHN3687_U_cr_n91));
   BUF_X32 FE_PHC1692_U_cr_N745 (.Z(FE_PHN1692_U_cr_N745), 
	.A(FE_PHN4759_U_cr_N745));
   BUF_X32 FE_PHC1690_U_cr_n92 (.Z(FE_PHN1690_U_cr_n92), 
	.A(FE_PHN3628_U_cr_n92));
   BUF_X32 FE_PHC1683_U_dsdc_N4229 (.Z(FE_PHN1683_U_dsdc_N4229), 
	.A(FE_PHN4785_U_dsdc_N4229));
   BUF_X32 FE_PHC1663_U_refctl_count_0_ (.Z(FE_PHN1663_U_refctl_count_0_), 
	.A(U_refctl_count_0_));
   CLKBUF_X1 FE_PHC1662_U_addrdec_n58 (.Z(FE_PHN1662_U_addrdec_n58), 
	.A(U_addrdec_n58));
   BUF_X32 FE_PHC1661_U_cr_N574 (.Z(FE_PHN1661_U_cr_N574), 
	.A(U_cr_N574));
   BUF_X32 FE_PHC1659_U_dsdc_n386 (.Z(FE_PHN1659_U_dsdc_n386), 
	.A(FE_PHN4613_U_dsdc_n386));
   BUF_X32 FE_PHC1658_U_dsdc_n403 (.Z(FE_PHN1658_U_dsdc_n403), 
	.A(U_dsdc_n403));
   BUF_X32 FE_PHC1656_U_cr_N577 (.Z(FE_PHN1656_U_cr_N577), 
	.A(U_cr_N577));
   BUF_X32 FE_PHC1647_U_cr_n86 (.Z(FE_PHN1647_U_cr_n86), 
	.A(FE_PHN3349_U_cr_n86));
   CLKBUF_X1 FE_PHC1645_U_cr_n65 (.Z(FE_PHN1645_U_cr_n65), 
	.A(FE_PHN4966_U_cr_n65));
   BUF_X32 FE_PHC1643_U_cr_N688 (.Z(FE_PHN1643_U_cr_N688), 
	.A(U_cr_N688));
   BUF_X32 FE_PHC1642_U_cr_n119 (.Z(FE_PHN1642_U_cr_n119), 
	.A(U_cr_n119));
   BUF_X32 FE_PHC1641_U_addrdec_n345 (.Z(FE_PHN1641_U_addrdec_n345), 
	.A(U_addrdec_n345));
   BUF_X16 FE_PHC1640_U_cr_N576 (.Z(FE_PHN1640_U_cr_N576), 
	.A(U_cr_N576));
   BUF_X32 FE_PHC1639_U_cr_N733 (.Z(FE_PHN1639_U_cr_N733), 
	.A(FE_PHN3379_U_cr_N733));
   BUF_X32 FE_PHC1638_U_cr_N689 (.Z(FE_PHN1638_U_cr_N689), 
	.A(U_cr_N689));
   BUF_X32 FE_PHC1637_U_cr_N734 (.Z(FE_PHN1637_U_cr_N734), 
	.A(FE_PHN3389_U_cr_N734));
   BUF_X32 FE_PHC1634_U_cr_n167 (.Z(FE_PHN1634_U_cr_n167), 
	.A(U_cr_n167));
   BUF_X32 FE_PHC1628_U_cr_n286 (.Z(FE_PHN1628_U_cr_n286), 
	.A(FE_PHN4589_U_cr_n286));
   BUF_X32 FE_PHC1623_U_dsdc_n366 (.Z(FE_PHN1623_U_dsdc_n366), 
	.A(FE_PHN4878_U_dsdc_n366));
   BUF_X32 FE_PHC1617_U_cr_N406 (.Z(FE_PHN1617_U_cr_N406), 
	.A(U_cr_N406));
   BUF_X32 FE_PHC1608_cr_reg_data_out_18_ (.Z(FE_PHN1608_cr_reg_data_out_18_), 
	.A(cr_reg_data_out[18]));
   CLKBUF_X1 FE_PHC1597_U_dmc_n1 (.Z(FE_PHN1597_U_dmc_n1), 
	.A(U_dmc_n1));
   BUF_X16 FE_PHC1596_U_dsdc_n1091 (.Z(FE_PHN1596_U_dsdc_n1091), 
	.A(U_dsdc_n1091));
   CLKBUF_X1 FE_PHC1594_U_addrdec_N133 (.Z(FE_PHN1594_U_addrdec_N133), 
	.A(U_addrdec_N133));
   BUF_X32 FE_PHC1593_U_dsdc_bm_bank_status_1_ (.Z(FE_PHN1593_U_dsdc_bm_bank_status_1_), 
	.A(U_dsdc_bm_bank_status_1_));
   BUF_X32 FE_PHC1590_U_dsdc_N4322 (.Z(FE_PHN1590_U_dsdc_N4322), 
	.A(U_dsdc_N4322));
   BUF_X32 FE_PHC1589_U_cr_N552 (.Z(FE_PHN1589_U_cr_N552), 
	.A(U_cr_N552));
   BUF_X32 FE_PHC1587_U_cr_N391 (.Z(FE_PHN1587_U_cr_N391), 
	.A(U_cr_N391));
   BUF_X32 FE_PHC1585_U_dsdc_n1094 (.Z(FE_PHN1585_U_dsdc_n1094), 
	.A(U_dsdc_n1094));
   BUF_X32 FE_PHC1583_U_refctl_n80 (.Z(FE_PHN1583_U_refctl_n80), 
	.A(U_refctl_n80));
   BUF_X32 FE_PHC1582_U_dsdc_N4340 (.Z(FE_PHN1582_U_dsdc_N4340), 
	.A(FE_PHN4537_U_dsdc_N4340));
   BUF_X32 FE_PHC1581_U_dsdc_N4482 (.Z(FE_PHN1581_U_dsdc_N4482), 
	.A(FE_PHN4473_U_dsdc_N4482));
   BUF_X32 FE_PHC1580_U_dsdc_N4436 (.Z(FE_PHN1580_U_dsdc_N4436), 
	.A(FE_PHN4521_U_dsdc_N4436));
   BUF_X32 FE_PHC1578_U_dsdc_N4434 (.Z(FE_PHN1578_U_dsdc_N4434), 
	.A(FE_PHN4546_U_dsdc_N4434));
   BUF_X32 FE_PHC1576_U_dsdc_N4481 (.Z(FE_PHN1576_U_dsdc_N4481), 
	.A(FE_PHN4498_U_dsdc_N4481));
   BUF_X32 FE_PHC1575_U_dsdc_N4435 (.Z(FE_PHN1575_U_dsdc_N4435), 
	.A(FE_PHN4443_U_dsdc_N4435));
   BUF_X32 FE_PHC1574_U_refctl_n78 (.Z(FE_PHN1574_U_refctl_n78), 
	.A(U_refctl_n78));
   BUF_X32 FE_PHC1573_U_dsdc_N4487 (.Z(FE_PHN1573_U_dsdc_N4487), 
	.A(FE_PHN4423_U_dsdc_N4487));
   BUF_X32 FE_PHC1572_U_dsdc_N4485 (.Z(FE_PHN1572_U_dsdc_N4485), 
	.A(FE_PHN4365_U_dsdc_N4485));
   BUF_X32 FE_PHC1570_U_dsdc_N4346 (.Z(FE_PHN1570_U_dsdc_N4346), 
	.A(FE_PHN4323_U_dsdc_N4346));
   BUF_X32 FE_PHC1569_U_cr_N735 (.Z(FE_PHN1569_U_cr_N735), 
	.A(FE_PHN3378_U_cr_N735));
   BUF_X32 FE_PHC1568_U_cr_N466 (.Z(FE_PHN1568_U_cr_N466), 
	.A(U_cr_N466));
   BUF_X32 FE_PHC1567_U_cr_N690 (.Z(FE_PHN1567_U_cr_N690), 
	.A(FE_PHN3456_U_cr_N690));
   BUF_X32 FE_PHC1557_U_refctl_count_next_1_ (.Z(FE_PHN1557_U_refctl_count_next_1_), 
	.A(FE_PHN4934_U_refctl_count_next_1_));
   BUF_X32 FE_PHC1555_U_cr_N571 (.Z(FE_PHN1555_U_cr_N571), 
	.A(U_cr_N571));
   BUF_X32 FE_PHC1549_U_refctl_n89 (.Z(FE_PHN1549_U_refctl_n89), 
	.A(U_refctl_n89));
   BUF_X32 FE_PHC1548_U_refctl_n85 (.Z(FE_PHN1548_U_refctl_n85), 
	.A(U_refctl_n85));
   BUF_X32 FE_PHC1537_U_cr_N553 (.Z(FE_PHN1537_U_cr_N553), 
	.A(FE_PHN4568_U_cr_N553));
   BUF_X32 FE_PHC1536_U_cr_N478 (.Z(FE_PHN1536_U_cr_N478), 
	.A(FE_PHN3751_U_cr_N478));
   BUF_X32 FE_PHC1535_U_cr_N477 (.Z(FE_PHN1535_U_cr_N477), 
	.A(FE_PHN3669_U_cr_N477));
   BUF_X32 FE_PHC1534_U_cr_N637 (.Z(FE_PHN1534_U_cr_N637), 
	.A(FE_PHN3768_U_cr_N637));
   BUF_X32 FE_PHC1533_U_cr_N639 (.Z(FE_PHN1533_U_cr_N639), 
	.A(FE_PHN3659_U_cr_N639));
   BUF_X32 FE_PHC1532_U_cr_N638 (.Z(FE_PHN1532_U_cr_N638), 
	.A(FE_PHN4483_U_cr_N638));
   BUF_X32 FE_PHC1531_U_cr_N694 (.Z(FE_PHN1531_U_cr_N694), 
	.A(FE_PHN3714_U_cr_N694));
   BUF_X32 FE_PHC1530_U_cr_N695 (.Z(FE_PHN1530_U_cr_N695), 
	.A(FE_PHN3702_U_cr_N695));
   BUF_X32 FE_PHC1529_U_dsdc_n215 (.Z(FE_PHN1529_U_dsdc_n215), 
	.A(U_dsdc_n215));
   BUF_X32 FE_PHC1528_U_cr_n88 (.Z(FE_PHN1528_U_cr_n88), 
	.A(FE_PHN3672_U_cr_n88));
   BUF_X32 FE_PHC1526_U_cr_N407 (.Z(FE_PHN1526_U_cr_N407), 
	.A(U_cr_N407));
   BUF_X16 FE_PHC1524_U_cr_N408 (.Z(FE_PHN1524_U_cr_N408), 
	.A(U_cr_N408));
   BUF_X32 FE_PHC1523_U_cr_N409 (.Z(FE_PHN1523_U_cr_N409), 
	.A(FE_PHN4594_U_cr_N409));
   BUF_X32 FE_PHC1522_U_cr_n94 (.Z(FE_PHN1522_U_cr_n94), 
	.A(FE_PHN3619_U_cr_n94));
   BUF_X32 FE_PHC1521_U_dsdc_n423 (.Z(FE_PHN1521_U_dsdc_n423), 
	.A(FE_PHN3160_U_dsdc_n423));
   BUF_X32 FE_PHC1520_U_cr_n75 (.Z(FE_PHN1520_U_cr_n75), 
	.A(FE_PHN3476_U_cr_n75));
   BUF_X32 FE_PHC1519_U_cr_n74 (.Z(FE_PHN1519_U_cr_n74), 
	.A(FE_PHN3475_U_cr_n74));
   BUF_X32 FE_PHC1518_U_cr_n76 (.Z(FE_PHN1518_U_cr_n76), 
	.A(FE_PHN3215_U_cr_n76));
   BUF_X32 FE_PHC1517_U_cr_n78 (.Z(FE_PHN1517_U_cr_n78), 
	.A(U_cr_n78));
   BUF_X32 FE_PHC1516_U_cr_n79 (.Z(FE_PHN1516_U_cr_n79), 
	.A(U_cr_n79));
   BUF_X32 FE_PHC1514_U_cr_N311 (.Z(FE_PHN1514_U_cr_N311), 
	.A(FE_PHN3250_U_cr_N311));
   BUF_X16 FE_PHC1504_U_cr_N551 (.Z(FE_PHN1504_U_cr_N551), 
	.A(U_cr_N551));
   BUF_X32 FE_PHC1497_U_dsdc_n1238 (.Z(FE_PHN1497_U_dsdc_n1238), 
	.A(U_dsdc_n1238));
   BUF_X32 FE_PHC1496_U_dsdc_N4369 (.Z(FE_PHN1496_U_dsdc_N4369), 
	.A(U_dsdc_N4369));
   BUF_X32 FE_PHC1495_U_dsdc_N4416 (.Z(FE_PHN1495_U_dsdc_N4416), 
	.A(U_dsdc_N4416));
   BUF_X32 FE_PHC1494_U_refctl_next_state_0_ (.Z(FE_PHN1494_U_refctl_next_state_0_), 
	.A(FE_PHN3449_U_refctl_next_state_0_));
   BUF_X32 FE_PHC1493_U_dsdc_n282 (.Z(FE_PHN1493_U_dsdc_n282), 
	.A(FE_PHN3443_U_dsdc_n282));
   BUF_X32 FE_PHC1492_U_dsdc_n1180 (.Z(FE_PHN1492_U_dsdc_n1180), 
	.A(U_dsdc_n1180));
   BUF_X32 FE_PHC1491_U_dsdc_N4140 (.Z(FE_PHN1491_U_dsdc_N4140), 
	.A(FE_PHN4587_U_dsdc_N4140));
   BUF_X32 FE_PHC1489_U_dsdc_N4429 (.Z(FE_PHN1489_U_dsdc_N4429), 
	.A(FE_PHN3337_U_dsdc_N4429));
   BUF_X32 FE_PHC1487_U_dsdc_n1194 (.Z(FE_PHN1487_U_dsdc_n1194), 
	.A(U_dsdc_n1194));
   BUF_X32 FE_PHC1486_U_dsdc_N4476 (.Z(FE_PHN1486_U_dsdc_N4476), 
	.A(FE_PHN3328_U_dsdc_N4476));
   BUF_X32 FE_PHC1485_U_dsdc_N4442 (.Z(FE_PHN1485_U_dsdc_N4442), 
	.A(FE_PHN4502_U_dsdc_N4442));
   BUF_X32 FE_PHC1484_U_dsdc_n319 (.Z(FE_PHN1484_U_dsdc_n319), 
	.A(FE_PHN3464_U_dsdc_n319));
   BUF_X32 FE_PHC1483_U_dsdc_n280 (.Z(FE_PHN1483_U_dsdc_n280), 
	.A(FE_PHN3083_U_dsdc_n280));
   CLKBUF_X1 FE_PHC1482_U_cr_n151 (.Z(FE_PHN1482_U_cr_n151), 
	.A(U_cr_n151));
   BUF_X32 FE_PHC1481_U_dsdc_N4489 (.Z(FE_PHN1481_U_dsdc_N4489), 
	.A(FE_PHN4381_U_dsdc_N4489));
   BUF_X32 FE_PHC1480_U_dsdc_n259 (.Z(FE_PHN1480_U_dsdc_n259), 
	.A(FE_PHN3317_U_dsdc_n259));
   BUF_X32 FE_PHC1479_U_dsdc_n260 (.Z(FE_PHN1479_U_dsdc_n260), 
	.A(FE_PHN3316_U_dsdc_n260));
   BUF_X32 FE_PHC1478_U_dsdc_n261 (.Z(FE_PHN1478_U_dsdc_n261), 
	.A(FE_PHN3314_U_dsdc_n261));
   CLKBUF_X1 FE_PHC1477_U_cr_stmg0r_0_ (.Z(FE_PHN1477_U_cr_stmg0r_0_), 
	.A(U_cr_stmg0r_0_));
   BUF_X32 FE_PHC1476_U_refctl_count_next_15_ (.Z(FE_PHN1476_U_refctl_count_next_15_), 
	.A(FE_PHN3326_U_refctl_count_next_15_));
   BUF_X32 FE_PHC1475_cr_s_data_width_early_0_ (.Z(FE_PHN1475_cr_s_data_width_early_0_), 
	.A(FE_PHN3111_cr_s_data_width_early_0_));
   BUF_X32 FE_PHC1473_U_cr_n27 (.Z(FE_PHN1473_U_cr_n27), 
	.A(U_cr_n27));
   BUF_X32 FE_PHC1470_U_dsdc_write_start_nxt (.Z(FE_PHN1470_U_dsdc_write_start_nxt), 
	.A(U_dsdc_write_start_nxt));
   BUF_X32 FE_PHC1456_U_cr_N310 (.Z(FE_PHN1456_U_cr_N310), 
	.A(FE_PHN3683_U_cr_N310));
   BUF_X32 FE_PHC1455_U_cr_N303 (.Z(FE_PHN1455_U_cr_N303), 
	.A(FE_PHN4398_U_cr_N303));
   BUF_X32 FE_PHC1449_U_cr_N561 (.Z(FE_PHN1449_U_cr_N561), 
	.A(U_cr_N561));
   BUF_X32 FE_PHC1447_U_dsdc_N429 (.Z(FE_PHN1447_U_dsdc_N429), 
	.A(U_dsdc_N429));
   BUF_X32 FE_PHC1445_U_dsdc_n157 (.Z(FE_PHN1445_U_dsdc_n157), 
	.A(U_dsdc_n157));
   BUF_X32 FE_PHC1444_U_cr_N646 (.Z(FE_PHN1444_U_cr_N646), 
	.A(FE_PHN4470_U_cr_N646));
   BUF_X32 FE_PHC1430_U_dsdc_N4228 (.Z(FE_PHN1430_U_dsdc_N4228), 
	.A(FE_PHN5042_U_dsdc_N4228));
   BUF_X32 FE_PHC1427_cr_reg_data_out_17_ (.Z(FE_PHN1427_cr_reg_data_out_17_), 
	.A(cr_reg_data_out[17]));
   BUF_X32 FE_PHC1424_U_refctl_count_12_ (.Z(FE_PHN1424_U_refctl_count_12_), 
	.A(U_refctl_count_12_));
   BUF_X32 FE_PHC1421_U_refctl_count_10_ (.Z(FE_PHN1421_U_refctl_count_10_), 
	.A(U_refctl_count_10_));
   BUF_X32 FE_PHC1420_U_refctl_count_8_ (.Z(FE_PHN1420_U_refctl_count_8_), 
	.A(U_refctl_count_8_));
   BUF_X32 FE_PHC1419_U_refctl_count_6_ (.Z(FE_PHN1419_U_refctl_count_6_), 
	.A(U_refctl_count_6_));
   BUF_X32 FE_PHC1418_U_dmc_data_cnt_2_ (.Z(FE_PHN1418_U_dmc_data_cnt_2_), 
	.A(U_dmc_data_cnt_2_));
   BUF_X32 FE_PHC1416_U_dsdc_r_col_addr_1_ (.Z(FE_PHN1416_U_dsdc_r_col_addr_1_), 
	.A(U_dsdc_r_col_addr_1_));
   BUF_X32 FE_PHC1415_U_refctl_n86 (.Z(FE_PHN1415_U_refctl_n86), 
	.A(U_refctl_n86));
   BUF_X32 FE_PHC1414_U_refctl_count_next_14_ (.Z(FE_PHN1414_U_refctl_count_next_14_), 
	.A(U_refctl_count_next_14_));
   BUF_X32 FE_PHC1413_U_dsdc_N4281 (.Z(FE_PHN1413_U_dsdc_N4281), 
	.A(U_dsdc_N4281));
   BUF_X32 FE_PHC1412_U_cr_N634 (.Z(FE_PHN1412_U_cr_N634), 
	.A(U_cr_N634));
   BUF_X32 FE_PHC1411_U_refctl_n91 (.Z(FE_PHN1411_U_refctl_n91), 
	.A(U_refctl_n91));
   BUF_X32 FE_PHC1410_U_dsdc_N4413 (.Z(FE_PHN1410_U_dsdc_N4413), 
	.A(U_dsdc_N4413));
   BUF_X32 FE_PHC1409_U_cr_n85 (.Z(FE_PHN1409_U_cr_n85), 
	.A(FE_PHN3286_U_cr_n85));
   CLKBUF_X1 FE_PHC1407_U_cr_n104 (.Z(FE_PHN1407_U_cr_n104), 
	.A(U_cr_n104));
   BUF_X32 FE_PHC1403_U_refctl_count_next_5_ (.Z(FE_PHN1403_U_refctl_count_next_5_), 
	.A(U_refctl_count_next_5_));
   BUF_X32 FE_PHC1402_U_dsdc_n1462 (.Z(FE_PHN1402_U_dsdc_n1462), 
	.A(U_dsdc_n1462));
   CLKBUF_X1 FE_PHC1401_U_cr_cr_cs_1_ (.Z(FE_PHN1401_U_cr_cr_cs_1_), 
	.A(U_cr_cr_cs_1_));
   BUF_X32 FE_PHC1400_U_cr_n197 (.Z(FE_PHN1400_U_cr_n197), 
	.A(U_cr_n197));
   BUF_X32 FE_PHC1388_U_cr_N393 (.Z(FE_PHN1388_U_cr_N393), 
	.A(U_cr_N393));
   BUF_X32 FE_PHC1387_U_cr_N401 (.Z(FE_PHN1387_U_cr_N401), 
	.A(FE_PHN3575_U_cr_N401));
   BUF_X32 FE_PHC1386_U_cr_N474 (.Z(FE_PHN1386_U_cr_N474), 
	.A(FE_PHN3738_U_cr_N474));
   BUF_X32 FE_PHC1384_U_cr_N467 (.Z(FE_PHN1384_U_cr_N467), 
	.A(FE_PHN3579_U_cr_N467));
   BUF_X32 FE_PHC1383_U_cr_N736 (.Z(FE_PHN1383_U_cr_N736), 
	.A(FE_PHN4787_U_cr_N736));
   BUF_X32 FE_PHC1382_U_cr_N692 (.Z(FE_PHN1382_U_cr_N692), 
	.A(FE_PHN4428_U_cr_N692));
   BUF_X32 FE_PHC1381_U_dsdc_wr_cnt_nxt_1_ (.Z(FE_PHN1381_U_dsdc_wr_cnt_nxt_1_), 
	.A(U_dsdc_wr_cnt_nxt[1]));
   BUF_X32 FE_PHC1380_U_cr_N699 (.Z(FE_PHN1380_U_cr_N699), 
	.A(FE_PHN3722_U_cr_N699));
   BUF_X32 FE_PHC1378_U_cr_n90 (.Z(FE_PHN1378_U_cr_n90), 
	.A(FE_PHN3704_U_cr_n90));
   BUF_X32 FE_PHC1376_U_cr_N648 (.Z(FE_PHN1376_U_cr_N648), 
	.A(U_cr_N648));
   BUF_X32 FE_PHC1375_U_cr_N649 (.Z(FE_PHN1375_U_cr_N649), 
	.A(U_cr_N649));
   BUF_X32 FE_PHC1372_cr_reg_data_out_26_ (.Z(FE_PHN1372_cr_reg_data_out_26_), 
	.A(cr_reg_data_out[26]));
   BUF_X32 FE_PHC1371_cr_reg_data_out_19_ (.Z(FE_PHN1371_cr_reg_data_out_19_), 
	.A(cr_reg_data_out[19]));
   BUF_X32 FE_PHC1369_cr_reg_data_out_23_ (.Z(FE_PHN1369_cr_reg_data_out_23_), 
	.A(cr_reg_data_out[23]));
   CLKBUF_X1 FE_PHC1343_U_dsdc_n1276 (.Z(FE_PHN1343_U_dsdc_n1276), 
	.A(U_dsdc_n1276));
   BUF_X16 FE_PHC1340_U_dmc_data_cnt_nxt_1_ (.Z(FE_PHN1340_U_dmc_data_cnt_nxt_1_), 
	.A(U_dmc_data_cnt_nxt[1]));
   BUF_X16 FE_PHC1338_U_dsdc_cas_cnt_nxt_5_ (.Z(FE_PHN1338_U_dsdc_cas_cnt_nxt_5_), 
	.A(U_dsdc_cas_cnt_nxt[5]));
   BUF_X32 FE_PHC1337_U_dsdc_n363 (.Z(FE_PHN1337_U_dsdc_n363), 
	.A(U_dsdc_n363));
   BUF_X32 FE_PHC1336_U_dsdc_n364 (.Z(FE_PHN1336_U_dsdc_n364), 
	.A(U_dsdc_n364));
   BUF_X32 FE_PHC1335_U_dsdc_n1281 (.Z(FE_PHN1335_U_dsdc_n1281), 
	.A(U_dsdc_n1281));
   BUF_X32 FE_PHC1334_U_dsdc_n365 (.Z(FE_PHN1334_U_dsdc_n365), 
	.A(U_dsdc_n365));
   BUF_X32 FE_PHC1333_U_dsdc_n382 (.Z(FE_PHN1333_U_dsdc_n382), 
	.A(U_dsdc_n382));
   BUF_X32 FE_PHC1329_U_dsdc_N4339 (.Z(FE_PHN1329_U_dsdc_N4339), 
	.A(FE_PHN4605_U_dsdc_N4339));
   BUF_X32 FE_PHC1328_U_dsdc_n417 (.Z(FE_PHN1328_U_dsdc_n417), 
	.A(FE_PHN3195_U_dsdc_n417));
   BUF_X32 FE_PHC1326_U_dsdc_n258 (.Z(FE_PHN1326_U_dsdc_n258), 
	.A(U_dsdc_n258));
   BUF_X32 FE_PHC1323_U_dsdc_n393 (.Z(FE_PHN1323_U_dsdc_n393), 
	.A(FE_PHN4600_U_dsdc_n393));
   BUF_X32 FE_PHC1322_U_dsdc_N4337 (.Z(FE_PHN1322_U_dsdc_N4337), 
	.A(FE_PHN4593_U_dsdc_N4337));
   BUF_X32 FE_PHC1321_U_dsdc_n390 (.Z(FE_PHN1321_U_dsdc_n390), 
	.A(FE_PHN4592_U_dsdc_n390));
   BUF_X32 FE_PHC1315_U_dsdc_N4414 (.Z(FE_PHN1315_U_dsdc_N4414), 
	.A(U_dsdc_N4414));
   BUF_X32 FE_PHC1311_U_dsdc_N4427 (.Z(FE_PHN1311_U_dsdc_N4427), 
	.A(U_dsdc_N4427));
   BUF_X32 FE_PHC1310_U_dsdc_N4474 (.Z(FE_PHN1310_U_dsdc_N4474), 
	.A(U_dsdc_N4474));
   BUF_X32 FE_PHC1306_U_dsdc_N4380 (.Z(FE_PHN1306_U_dsdc_N4380), 
	.A(U_dsdc_N4380));
   BUF_X32 FE_PHC1303_U_dsdc_N4383 (.Z(FE_PHN1303_U_dsdc_N4383), 
	.A(FE_PHN4513_U_dsdc_N4383));
   BUF_X32 FE_PHC1300_U_dsdc_N4439 (.Z(FE_PHN1300_U_dsdc_N4439), 
	.A(FE_PHN4469_U_dsdc_N4439));
   BUF_X32 FE_PHC1299_U_dsdc_N4350 (.Z(FE_PHN1299_U_dsdc_N4350), 
	.A(FE_PHN4461_U_dsdc_N4350));
   BUF_X32 FE_PHC1295_U_dsdc_n418 (.Z(FE_PHN1295_U_dsdc_n418), 
	.A(FE_PHN3082_U_dsdc_n418));
   BUF_X32 FE_PHC1294_U_dsdc_N4333 (.Z(FE_PHN1294_U_dsdc_N4333), 
	.A(U_dsdc_N4333));
   BUF_X32 FE_PHC1292_U_dsdc_N4479 (.Z(FE_PHN1292_U_dsdc_N4479), 
	.A(FE_PHN4445_U_dsdc_N4479));
   BUF_X32 FE_PHC1291_U_dsdc_N4431 (.Z(FE_PHN1291_U_dsdc_N4431), 
	.A(FE_PHN4501_U_dsdc_N4431));
   BUF_X32 FE_PHC1288_U_dsdc_N4319 (.Z(FE_PHN1288_U_dsdc_N4319), 
	.A(U_dsdc_N4319));
   BUF_X32 FE_PHC1287_U_dsdc_N4473 (.Z(FE_PHN1287_U_dsdc_N4473), 
	.A(FE_PHN4503_U_dsdc_N4473));
   BUF_X32 FE_PHC1279_U_dsdc_N4484 (.Z(FE_PHN1279_U_dsdc_N4484), 
	.A(FE_PHN4304_U_dsdc_N4484));
   BUF_X32 FE_PHC1275_U_dsdc_N4426 (.Z(FE_PHN1275_U_dsdc_N4426), 
	.A(U_dsdc_N4426));
   BUF_X32 FE_PHC1271_U_dsdc_N4379 (.Z(FE_PHN1271_U_dsdc_N4379), 
	.A(U_dsdc_N4379));
   BUF_X32 FE_PHC1269_U_dsdc_n257 (.Z(FE_PHN1269_U_dsdc_n257), 
	.A(FE_PHN3312_U_dsdc_n257));
   BUF_X32 FE_PHC1268_U_dsdc_N4332 (.Z(FE_PHN1268_U_dsdc_N4332), 
	.A(FE_PHN3242_U_dsdc_N4332));
   BUF_X32 FE_PHC1262_U_dsdc_N4139 (.Z(FE_PHN1262_U_dsdc_N4139), 
	.A(FE_PHN3951_U_dsdc_N4139));
   BUF_X32 FE_PHC1256_U_cr_N573 (.Z(FE_PHN1256_U_cr_N573), 
	.A(U_cr_N573));
   BUF_X32 FE_PHC1254_U_cr_n55 (.Z(FE_PHN1254_U_cr_n55), 
	.A(U_cr_n55));
   BUF_X32 FE_PHC1253_U_cr_N306 (.Z(FE_PHN1253_U_cr_N306), 
	.A(FE_PHN4029_U_cr_N306));
   BUF_X32 FE_PHC1252_U_cr_N307 (.Z(FE_PHN1252_U_cr_N307), 
	.A(U_cr_N307));
   BUF_X32 FE_PHC1251_U_refctl_ref_req_next (.Z(FE_PHN1251_U_refctl_ref_req_next), 
	.A(U_refctl_ref_req_next));
   CLKBUF_X1 FE_PHC1249_U_dsdc_add_x_2600_1_n8 (.Z(FE_PHN1249_U_dsdc_add_x_2600_1_n8), 
	.A(U_dsdc_add_x_2600_1_n8));
   BUF_X32 FE_PHC1247_U_dsdc_n373 (.Z(FE_PHN1247_U_dsdc_n373), 
	.A(FE_PHN3216_U_dsdc_n373));
   BUF_X32 FE_PHC1243_U_cr_N655 (.Z(FE_PHN1243_U_cr_N655), 
	.A(U_cr_N655));
   BUF_X32 FE_PHC1242_U_dsdc_wtr_cnt_nxt_1_ (.Z(FE_PHN1242_U_dsdc_wtr_cnt_nxt_1_), 
	.A(FE_PHN3450_U_dsdc_wtr_cnt_nxt_1_));
   BUF_X32 FE_PHC1240_U_cr_N312 (.Z(FE_PHN1240_U_cr_N312), 
	.A(FE_PHN3249_U_cr_N312));
   BUF_X32 FE_PHC1236_cr_reg_data_out_25_ (.Z(FE_PHN1236_cr_reg_data_out_25_), 
	.A(cr_reg_data_out[25]));
   BUF_X32 FE_PHC1235_cr_reg_data_out_5_ (.Z(FE_PHN1235_cr_reg_data_out_5_), 
	.A(cr_reg_data_out[5]));
   BUF_X32 FE_PHC1234_cr_reg_data_out_4_ (.Z(FE_PHN1234_cr_reg_data_out_4_), 
	.A(cr_reg_data_out[4]));
   BUF_X32 FE_PHC1230_cr_reg_data_out_11_ (.Z(FE_PHN1230_cr_reg_data_out_11_), 
	.A(cr_reg_data_out[11]));
   CLKBUF_X1 FE_PHC1228_U_dmc_data_cnt_3_ (.Z(FE_PHN1228_U_dmc_data_cnt_3_), 
	.A(U_dmc_data_cnt_3_));
   CLKBUF_X1 FE_PHC1227_U_dsdc_cas_cnt_2_ (.Z(FE_PHN1227_U_dsdc_cas_cnt_2_), 
	.A(U_dsdc_cas_cnt_2_));
   CLKBUF_X1 FE_PHC1224_ctl_sd_in_sf_mode (.Z(FE_PHN1224_ctl_sd_in_sf_mode), 
	.A(ctl_sd_in_sf_mode));
   BUF_X32 FE_PHC1222_U_dsdc_bm_rc_cnt_2__2_ (.Z(FE_PHN1222_U_dsdc_bm_rc_cnt_2__2_), 
	.A(U_dsdc_bm_rc_cnt_2__2_));
   BUF_X32 FE_PHC1221_U_dsdc_bm_rc_cnt_1__2_ (.Z(FE_PHN1221_U_dsdc_bm_rc_cnt_1__2_), 
	.A(U_dsdc_bm_rc_cnt_1__2_));
   BUF_X16 FE_PHC1220_U_dsdc_n407 (.Z(FE_PHN1220_U_dsdc_n407), 
	.A(U_dsdc_n407));
   BUF_X32 FE_PHC1219_U_dsdc_bm_rc_cnt_3__2_ (.Z(FE_PHN1219_U_dsdc_bm_rc_cnt_3__2_), 
	.A(U_dsdc_bm_rc_cnt_3__2_));
   CLKBUF_X1 FE_PHC1218_U_dsdc_cas_cnt_nxt_1_ (.Z(FE_PHN1218_U_dsdc_cas_cnt_nxt_1_), 
	.A(U_dsdc_cas_cnt_nxt[1]));
   BUF_X8 FE_PHC1217_U_dmc_data_cnt_nxt_2_ (.Z(FE_PHN1217_U_dmc_data_cnt_nxt_2_), 
	.A(U_dmc_data_cnt_nxt[2]));
   BUF_X32 FE_PHC1216_U_dsdc_n413 (.Z(FE_PHN1216_U_dsdc_n413), 
	.A(U_dsdc_n413));
   BUF_X32 FE_PHC1215_U_dsdc_n409 (.Z(FE_PHN1215_U_dsdc_n409), 
	.A(FE_PHN4614_U_dsdc_n409));
   BUF_X16 FE_PHC1214_U_dsdc_n411 (.Z(FE_PHN1214_U_dsdc_n411), 
	.A(U_dsdc_n411));
   BUF_X32 FE_PHC1213_U_dsdc_rcar_cnt2_nxt_0_ (.Z(FE_PHN1213_U_dsdc_rcar_cnt2_nxt_0_), 
	.A(U_dsdc_rcar_cnt2_nxt[0]));
   BUF_X32 FE_PHC1212_U_dsdc_cas_latency_cnt_1_ (.Z(FE_PHN1212_U_dsdc_cas_latency_cnt_1_), 
	.A(U_dsdc_cas_latency_cnt_1_));
   BUF_X8 FE_PHC1211_U_dmc_data_cnt_nxt_5_ (.Z(FE_PHN1211_U_dmc_data_cnt_nxt_5_), 
	.A(U_dmc_data_cnt_nxt[5]));
   BUF_X32 FE_PHC1210_U_dsdc_n388 (.Z(FE_PHN1210_U_dsdc_n388), 
	.A(FE_PHN3191_U_dsdc_n388));
   BUF_X32 FE_PHC1209_U_dsdc_N4349 (.Z(FE_PHN1209_U_dsdc_N4349), 
	.A(FE_PHN4591_U_dsdc_N4349));
   BUF_X32 FE_PHC1208_U_dsdc_rcar_cnt1_nxt_1_ (.Z(FE_PHN1208_U_dsdc_rcar_cnt1_nxt_1_), 
	.A(U_dsdc_rcar_cnt1_nxt[1]));
   BUF_X32 FE_PHC1207_U_refctl_count_next_11_ (.Z(FE_PHN1207_U_refctl_count_next_11_), 
	.A(U_refctl_count_next_11_));
   BUF_X32 FE_PHC1206_U_dsdc_N4398 (.Z(FE_PHN1206_U_dsdc_N4398), 
	.A(FE_PHN4434_U_dsdc_N4398));
   BUF_X32 FE_PHC1205_U_dsdc_N4441 (.Z(FE_PHN1205_U_dsdc_N4441), 
	.A(FE_PHN4480_U_dsdc_N4441));
   BUF_X32 FE_PHC1204_U_dsdc_N4445 (.Z(FE_PHN1204_U_dsdc_N4445), 
	.A(FE_PHN4359_U_dsdc_N4445));
   BUF_X32 FE_PHC1203_U_refctl_count_next_9_ (.Z(FE_PHN1203_U_refctl_count_next_9_), 
	.A(U_refctl_count_next_9_));
   BUF_X32 FE_PHC1202_U_dsdc_N4394 (.Z(FE_PHN1202_U_dsdc_N4394), 
	.A(FE_PHN4388_U_dsdc_N4394));
   BUF_X32 FE_PHC1201_U_refctl_count_next_13_ (.Z(FE_PHN1201_U_refctl_count_next_13_), 
	.A(U_refctl_count_next_13_));
   BUF_X32 FE_PHC1200_U_dsdc_n1161 (.Z(FE_PHN1200_U_dsdc_n1161), 
	.A(U_dsdc_n1161));
   BUF_X32 FE_PHC1199_U_dsdc_rp_cnt1_nxt_2_ (.Z(FE_PHN1199_U_dsdc_rp_cnt1_nxt_2_), 
	.A(FE_PHN3045_U_dsdc_rp_cnt1_nxt_2_));
   BUF_X32 FE_PHC1198_U_dsdc_rp_cnt1_nxt_0_ (.Z(FE_PHN1198_U_dsdc_rp_cnt1_nxt_0_), 
	.A(FE_PHN3503_U_dsdc_rp_cnt1_nxt_0_));
   BUF_X32 FE_PHC1185_U_refctl_count_next_7_ (.Z(FE_PHN1185_U_refctl_count_next_7_), 
	.A(U_refctl_count_next_7_));
   BUF_X32 FE_PHC1176_U_cr_n84 (.Z(FE_PHN1176_U_cr_n84), 
	.A(U_cr_n84));
   BUF_X32 FE_PHC1173_U_dsdc_wr_cnt_nxt_0_ (.Z(FE_PHN1173_U_dsdc_wr_cnt_nxt_0_), 
	.A(FE_PHN3327_U_dsdc_wr_cnt_nxt_0_));
   BUF_X32 FE_PHC1171_U_cr_n297 (.Z(FE_PHN1171_U_cr_n297), 
	.A(U_cr_n297));
   BUF_X32 FE_PHC1170_U_cr_N313 (.Z(FE_PHN1170_U_cr_N313), 
	.A(FE_PHN4841_U_cr_N313));
   BUF_X32 FE_PHC1169_cr_reg_data_out_24_ (.Z(FE_PHN1169_cr_reg_data_out_24_), 
	.A(FE_PHN3283_cr_reg_data_out_24_));
   BUF_X32 FE_PHC1168_U_cr_N413 (.Z(FE_PHN1168_U_cr_N413), 
	.A(FE_PHN3043_U_cr_N413));
   BUF_X32 FE_PHC1167_cr_reg_data_out_1_ (.Z(FE_PHN1167_cr_reg_data_out_1_), 
	.A(cr_reg_data_out[1]));
   BUF_X32 FE_PHC1166_cr_reg_data_out_29_ (.Z(FE_PHN1166_cr_reg_data_out_29_), 
	.A(cr_reg_data_out[29]));
   BUF_X32 FE_PHC1165_cr_reg_data_out_14_ (.Z(FE_PHN1165_cr_reg_data_out_14_), 
	.A(cr_reg_data_out[14]));
   BUF_X32 FE_PHC1163_U_cr_n482 (.Z(FE_PHN1163_U_cr_n482), 
	.A(U_cr_n482));
   CLKBUF_X1 FE_PHC1161_U_dsdc_n1339 (.Z(FE_PHN1161_U_dsdc_n1339), 
	.A(U_dsdc_n1339));
   CLKBUF_X1 FE_PHC1160_U_dmc_n48 (.Z(FE_PHN1160_U_dmc_n48), 
	.A(U_dmc_n48));
   BUF_X32 FE_PHC1158_U_dsdc_bm_ras_cnt_max_1_ (.Z(FE_PHN1158_U_dsdc_bm_ras_cnt_max_1_), 
	.A(U_dsdc_bm_ras_cnt_max_1_));
   BUF_X32 FE_PHC1156_U_dsdc_n1182 (.Z(FE_PHN1156_U_dsdc_n1182), 
	.A(U_dsdc_n1182));
   BUF_X32 FE_PHC1155_U_dsdc_n1210 (.Z(FE_PHN1155_U_dsdc_n1210), 
	.A(U_dsdc_n1210));
   BUF_X32 FE_PHC1154_U_dsdc_n1196 (.Z(FE_PHN1154_U_dsdc_n1196), 
	.A(U_dsdc_n1196));
   BUF_X32 FE_PHC1153_U_dsdc_cas_latency_cnt_3_ (.Z(FE_PHN1153_U_dsdc_cas_latency_cnt_3_), 
	.A(U_dsdc_cas_latency_cnt_3_));
   BUF_X32 FE_PHC1152_U_dsdc_r_row_addr_5_ (.Z(FE_PHN1152_U_dsdc_r_row_addr_5_), 
	.A(U_dsdc_r_row_addr_5_));
   BUF_X32 FE_PHC1151_U_dsdc_r_row_addr_8_ (.Z(FE_PHN1151_U_dsdc_r_row_addr_8_), 
	.A(U_dsdc_r_row_addr_8_));
   BUF_X32 FE_PHC1150_U_cr_sctlr_14_ (.Z(FE_PHN1150_U_cr_sctlr_14_), 
	.A(U_cr_sctlr_14_));
   BUF_X32 FE_PHC1149_U_dsdc_r_row_addr_12_ (.Z(FE_PHN1149_U_dsdc_r_row_addr_12_), 
	.A(U_dsdc_r_row_addr_12_));
   BUF_X32 FE_PHC1148_U_dsdc_r_row_addr_10_ (.Z(FE_PHN1148_U_dsdc_r_row_addr_10_), 
	.A(U_dsdc_r_row_addr_10_));
   BUF_X32 FE_PHC1147_U_dsdc_r_row_addr_4_ (.Z(FE_PHN1147_U_dsdc_r_row_addr_4_), 
	.A(U_dsdc_r_row_addr_4_));
   BUF_X32 FE_PHC1146_U_dsdc_r_row_addr_6_ (.Z(FE_PHN1146_U_dsdc_r_row_addr_6_), 
	.A(U_dsdc_r_row_addr_6_));
   BUF_X32 FE_PHC1144_U_dsdc_wrapped_pop_flag_nxt (.Z(FE_PHN1144_U_dsdc_wrapped_pop_flag_nxt), 
	.A(FE_PHN4497_U_dsdc_wrapped_pop_flag_nxt));
   BUF_X32 FE_PHC1143_U_dsdc_num_init_ref_cnt_nxt_2_ (.Z(FE_PHN1143_U_dsdc_num_init_ref_cnt_nxt_2_), 
	.A(FE_PHN3110_U_dsdc_num_init_ref_cnt_nxt_2_));
   BUF_X16 FE_PHC1140_U_refctl_count_next_2_ (.Z(FE_PHN1140_U_refctl_count_next_2_), 
	.A(U_refctl_count_next_2_));
   BUF_X32 FE_PHC1127_U_cr_N305 (.Z(FE_PHN1127_U_cr_N305), 
	.A(FE_PHN4409_U_cr_N305));
   BUF_X32 FE_PHC1124_U_cr_N645 (.Z(FE_PHN1124_U_cr_N645), 
	.A(FE_PHN3736_U_cr_N645));
   BUF_X32 FE_PHC1123_U_dsdc_n372 (.Z(FE_PHN1123_U_dsdc_n372), 
	.A(FE_PHN3227_U_dsdc_n372));
   BUF_X32 FE_PHC1122_U_dsdc_n371 (.Z(FE_PHN1122_U_dsdc_n371), 
	.A(FE_PHN5012_U_dsdc_n371));
   BUF_X32 FE_PHC1121_U_dsdc_n367 (.Z(FE_PHN1121_U_dsdc_n367), 
	.A(FE_PHN3169_U_dsdc_n367));
   BUF_X32 FE_PHC1120_U_dsdc_n369 (.Z(FE_PHN1120_U_dsdc_n369), 
	.A(FE_PHN3162_U_dsdc_n369));
   BUF_X32 FE_PHC1119_U_cr_N653 (.Z(FE_PHN1119_U_cr_N653), 
	.A(U_cr_N653));
   BUF_X32 FE_PHC1118_U_cr_N654 (.Z(FE_PHN1118_U_cr_N654), 
	.A(U_cr_N654));
   BUF_X32 FE_PHC1117_cr_reg_data_out_20_ (.Z(FE_PHN1117_cr_reg_data_out_20_), 
	.A(cr_reg_data_out[20]));
   BUF_X32 FE_PHC1116_U_cr_N415 (.Z(FE_PHN1116_U_cr_N415), 
	.A(U_cr_N415));
   BUF_X32 FE_PHC1103_U_cr_n455 (.Z(FE_PHN1103_U_cr_n455), 
	.A(FE_PHN5237_U_cr_n455));
   CLKBUF_X1 FE_PHC1101_U_dsdc_n1275 (.Z(FE_PHN1101_U_dsdc_n1275), 
	.A(FE_PHN3086_U_dsdc_n1275));
   BUF_X32 FE_PHC1099_U_dsdc_n404 (.Z(FE_PHN1099_U_dsdc_n404), 
	.A(U_dsdc_n404));
   BUF_X16 FE_PHC1098_U_dsdc_N4334 (.Z(FE_PHN1098_U_dsdc_N4334), 
	.A(U_dsdc_N4334));
   BUF_X8 FE_PHC1097_U_dsdc_N4428 (.Z(FE_PHN1097_U_dsdc_N4428), 
	.A(U_dsdc_N4428));
   BUF_X8 FE_PHC1096_U_dsdc_N4381 (.Z(FE_PHN1096_U_dsdc_N4381), 
	.A(U_dsdc_N4381));
   BUF_X32 FE_PHC1095_U_dsdc_n392 (.Z(FE_PHN1095_U_dsdc_n392), 
	.A(U_dsdc_n392));
   BUF_X32 FE_PHC1094_U_dsdc_n394 (.Z(FE_PHN1094_U_dsdc_n394), 
	.A(FE_PHN3461_U_dsdc_n394));
   BUF_X32 FE_PHC1093_U_dsdc_n340 (.Z(FE_PHN1093_U_dsdc_n340), 
	.A(U_dsdc_n340));
   BUF_X16 FE_PHC1092_U_dsdc_N4128 (.Z(FE_PHN1092_U_dsdc_N4128), 
	.A(U_dsdc_N4128));
   BUF_X32 FE_PHC1091_U_refctl_count_next_3_ (.Z(FE_PHN1091_U_refctl_count_next_3_), 
	.A(FE_PHN3343_U_refctl_count_next_3_));
   BUF_X32 FE_PHC1090_U_dsdc_N4460 (.Z(FE_PHN1090_U_dsdc_N4460), 
	.A(U_dsdc_N4460));
   BUF_X32 FE_PHC1089_U_refctl_count_next_4_ (.Z(FE_PHN1089_U_refctl_count_next_4_), 
	.A(FE_PHN4410_U_refctl_count_next_4_));
   BUF_X32 FE_PHC1088_U_cr_n558 (.Z(FE_PHN1088_U_cr_n558), 
	.A(U_cr_n558));
   BUF_X32 FE_PHC1087_U_dsdc_rp_cnt1_nxt_1_ (.Z(FE_PHN1087_U_dsdc_rp_cnt1_nxt_1_), 
	.A(FE_PHN3238_U_dsdc_rp_cnt1_nxt_1_));
   BUF_X32 FE_PHC1083_U_cr_N650 (.Z(FE_PHN1083_U_cr_N650), 
	.A(U_cr_N650));
   BUF_X32 FE_PHC1082_U_cr_n77 (.Z(FE_PHN1082_U_cr_n77), 
	.A(FE_PHN3485_U_cr_n77));
   BUF_X32 FE_PHC1081_U_dsdc_n1671 (.Z(FE_PHN1081_U_dsdc_n1671), 
	.A(U_dsdc_n1671));
   BUF_X32 FE_PHC1080_cr_reg_data_out_0_ (.Z(FE_PHN1080_cr_reg_data_out_0_), 
	.A(cr_reg_data_out[0]));
   BUF_X32 FE_PHC1077_cr_reg_data_out_22_ (.Z(FE_PHN1077_cr_reg_data_out_22_), 
	.A(cr_reg_data_out[22]));
   BUF_X32 FE_PHC1076_U_cr_N418 (.Z(FE_PHN1076_U_cr_N418), 
	.A(U_cr_N418));
   CLKBUF_X1 FE_PHC1064_cr_row_addr_width_3_ (.Z(FE_PHN1064_cr_row_addr_width_3_), 
	.A(cr_row_addr_width[3]));
   BUF_X32 FE_PHC1062_U_dsdc_init_cnt_3_ (.Z(FE_PHN1062_U_dsdc_init_cnt_3_), 
	.A(U_dsdc_init_cnt_3_));
   BUF_X8 FE_PHC1061_U_dsdc_N4475 (.Z(FE_PHN1061_U_dsdc_N4475), 
	.A(U_dsdc_N4475));
   BUF_X16 FE_PHC1060_U_dsdc_N4321 (.Z(FE_PHN1060_U_dsdc_N4321), 
	.A(U_dsdc_N4321));
   BUF_X16 FE_PHC1059_U_dsdc_N4462 (.Z(FE_PHN1059_U_dsdc_N4462), 
	.A(U_dsdc_N4462));
   BUF_X16 FE_PHC1058_U_dsdc_N4141 (.Z(FE_PHN1058_U_dsdc_N4141), 
	.A(U_dsdc_N4141));
   BUF_X16 FE_PHC1057_U_dsdc_N4415 (.Z(FE_PHN1057_U_dsdc_N4415), 
	.A(U_dsdc_N4415));
   CLKBUF_X1 FE_PHC1056_U_dmc_terminate (.Z(FE_PHN1056_U_dmc_terminate), 
	.A(U_dmc_terminate));
   BUF_X16 FE_PHC1055_U_dsdc_N4368 (.Z(FE_PHN1055_U_dsdc_N4368), 
	.A(U_dsdc_N4368));
   BUF_X32 FE_PHC1054_U_dsdc_rp_cnt2_nxt_0_ (.Z(FE_PHN1054_U_dsdc_rp_cnt2_nxt_0_), 
	.A(FE_PHN3085_U_dsdc_rp_cnt2_nxt_0_));
   BUF_X32 FE_PHC1053_U_dsdc_rcar_cnt1_nxt_3_ (.Z(FE_PHN1053_U_dsdc_rcar_cnt1_nxt_3_), 
	.A(FE_PHN3187_U_dsdc_rcar_cnt1_nxt_3_));
   CLKBUF_X1 FE_PHC1052_U_cr_n127 (.Z(FE_PHN1052_U_cr_n127), 
	.A(U_cr_n127));
   BUF_X32 FE_PHC1051_U_dsdc_rcar_cnt1_nxt_2_ (.Z(FE_PHN1051_U_dsdc_rcar_cnt1_nxt_2_), 
	.A(U_dsdc_rcar_cnt1_nxt[2]));
   BUF_X32 FE_PHC1050_U_dsdc_n218 (.Z(FE_PHN1050_U_dsdc_n218), 
	.A(U_dsdc_n218));
   BUF_X32 FE_PHC1048_U_cr_N550 (.Z(FE_PHN1048_U_cr_N550), 
	.A(FE_PHN3614_U_cr_N550));
   BUF_X32 FE_PHC1047_U_dsdc_n405 (.Z(FE_PHN1047_U_dsdc_n405), 
	.A(FE_PHN3613_U_dsdc_n405));
   BUF_X32 FE_PHC1046_U_dsdc_n380 (.Z(FE_PHN1046_U_dsdc_n380), 
	.A(FE_PHN3168_U_dsdc_n380));
   BUF_X32 FE_PHC1045_U_dsdc_n376 (.Z(FE_PHN1045_U_dsdc_n376), 
	.A(FE_PHN5056_U_dsdc_n376));
   BUF_X32 FE_PHC1044_U_cr_N652 (.Z(FE_PHN1044_U_cr_N652), 
	.A(U_cr_N652));
   BUF_X16 FE_PHC1043_U_cr_N412 (.Z(FE_PHN1043_U_cr_N412), 
	.A(U_cr_N412));
   BUF_X32 FE_PHC1042_cr_reg_data_out_28_ (.Z(FE_PHN1042_cr_reg_data_out_28_), 
	.A(cr_reg_data_out[28]));
   BUF_X32 FE_PHC1041_cr_reg_data_out_2_ (.Z(FE_PHN1041_cr_reg_data_out_2_), 
	.A(cr_reg_data_out[2]));
   BUF_X32 FE_PHC1040_U_cr_N419 (.Z(FE_PHN1040_U_cr_N419), 
	.A(U_cr_N419));
   CLKBUF_X1 FE_PHC1035_U_dsdc_n327 (.Z(FE_PHN1035_U_dsdc_n327), 
	.A(U_dsdc_n327));
   CLKBUF_X1 FE_PHC1034_cr_bank_addr_width_1_ (.Z(FE_PHN1034_cr_bank_addr_width_1_), 
	.A(cr_bank_addr_width[1]));
   BUF_X32 FE_PHC1033_U_dsdc_xsr_cnt_1_ (.Z(FE_PHN1033_U_dsdc_xsr_cnt_1_), 
	.A(U_dsdc_xsr_cnt_1_));
   BUF_X32 FE_PHC1032_U_dsdc_init_cnt_9_ (.Z(FE_PHN1032_U_dsdc_init_cnt_9_), 
	.A(U_dsdc_init_cnt_9_));
   BUF_X32 FE_PHC1031_U_dsdc_init_cnt_7_ (.Z(FE_PHN1031_U_dsdc_init_cnt_7_), 
	.A(U_dsdc_init_cnt_7_));
   BUF_X32 FE_PHC1030_U_dsdc_xsr_cnt_3_ (.Z(FE_PHN1030_U_dsdc_xsr_cnt_3_), 
	.A(U_dsdc_xsr_cnt_3_));
   BUF_X16 FE_PHC1029_U_dsdc_n414 (.Z(FE_PHN1029_U_dsdc_n414), 
	.A(U_dsdc_n414));
   BUF_X16 FE_PHC1028_U_dsdc_N4127 (.Z(FE_PHN1028_U_dsdc_N4127), 
	.A(U_dsdc_N4127));
   BUF_X32 FE_PHC1026_U_dsdc_N4367 (.Z(FE_PHN1026_U_dsdc_N4367), 
	.A(U_dsdc_N4367));
   BUF_X32 FE_PHC1023_U_dsdc_n387 (.Z(FE_PHN1023_U_dsdc_n387), 
	.A(U_dsdc_n387));
   BUF_X32 FE_PHC1020_U_dsdc_n1085 (.Z(FE_PHN1020_U_dsdc_n1085), 
	.A(U_dsdc_n1085));
   BUF_X32 FE_PHC1017_U_cr_N651 (.Z(FE_PHN1017_U_cr_N651), 
	.A(U_cr_N651));
   BUF_X32 FE_PHC1016_U_dsdc_n281 (.Z(FE_PHN1016_U_dsdc_n281), 
	.A(FE_PHN3156_U_dsdc_n281));
   BUF_X32 FE_PHC1015_U_cr_n295 (.Z(FE_PHN1015_U_cr_n295), 
	.A(U_cr_n295));
   BUF_X32 FE_PHC1014_U_cr_N567 (.Z(FE_PHN1014_U_cr_N567), 
	.A(U_cr_N567));
   BUF_X32 FE_PHC1013_U_cr_n73 (.Z(FE_PHN1013_U_cr_n73), 
	.A(FE_PHN3185_U_cr_n73));
   BUF_X32 FE_PHC1012_U_dsdc_n_2088_ (.Z(FE_PHN1012_U_dsdc_n_2088_), 
	.A(U_dsdc_n[2088]));
   BUF_X32 FE_PHC1001_U_dsdc_n391 (.Z(FE_PHN1001_U_dsdc_n391), 
	.A(FE_PHN3445_U_dsdc_n391));
   BUF_X16 FE_PHC1000_U_dmc_n14 (.Z(FE_PHN1000_U_dmc_n14), 
	.A(U_dmc_n14));
   BUF_X32 FE_PHC998_U_dsdc_n221 (.Z(FE_PHN998_U_dsdc_n221), 
	.A(FE_PHN4599_U_dsdc_n221));
   BUF_X32 FE_PHC997_U_dsdc_N4320 (.Z(FE_PHN997_U_dsdc_N4320), 
	.A(U_dsdc_N4320));
   BUF_X32 FE_PHC996_U_dsdc_num_init_ref_cnt_nxt_0_ (.Z(FE_PHN996_U_dsdc_num_init_ref_cnt_nxt_0_), 
	.A(FE_PHN3186_U_dsdc_num_init_ref_cnt_nxt_0_));
   BUF_X32 FE_PHC995_U_dsdc_N4283 (.Z(FE_PHN995_U_dsdc_N4283), 
	.A(U_dsdc_N4283));
   BUF_X32 FE_PHC994_U_dsdc_n212 (.Z(FE_PHN994_U_dsdc_n212), 
	.A(FE_PHN3241_U_dsdc_n212));
   BUF_X32 FE_PHC992_U_dsdc_n209 (.Z(FE_PHN992_U_dsdc_n209), 
	.A(FE_PHN4391_U_dsdc_n209));
   BUF_X32 FE_PHC990_U_dsdc_n_2089_ (.Z(FE_PHN990_U_dsdc_n_2089_), 
	.A(U_dsdc_n[2089]));
   BUF_X32 FE_PHC989_U_dsdc_n214 (.Z(FE_PHN989_U_dsdc_n214), 
	.A(FE_PHN4777_U_dsdc_n214));
   BUF_X32 FE_PHC988_U_cr_N298 (.Z(FE_PHN988_U_cr_N298), 
	.A(FE_PHN3692_U_cr_N298));
   BUF_X32 FE_PHC987_U_dsdc_n370 (.Z(FE_PHN987_U_dsdc_n370), 
	.A(FE_PHN3232_U_dsdc_n370));
   BUF_X32 FE_PHC986_U_dsdc_n368 (.Z(FE_PHN986_U_dsdc_n368), 
	.A(FE_PHN3228_U_dsdc_n368));
   BUF_X32 FE_PHC985_U_dsdc_n377 (.Z(FE_PHN985_U_dsdc_n377), 
	.A(FE_PHN3233_U_dsdc_n377));
   BUF_X32 FE_PHC984_U_dsdc_n381 (.Z(FE_PHN984_U_dsdc_n381), 
	.A(FE_PHN3221_U_dsdc_n381));
   BUF_X32 FE_PHC983_U_dsdc_n378 (.Z(FE_PHN983_U_dsdc_n378), 
	.A(FE_PHN5142_U_dsdc_n378));
   BUF_X32 FE_PHC982_U_cr_n93 (.Z(FE_PHN982_U_cr_n93), 
	.A(FE_PHN3212_U_cr_n93));
   BUF_X32 FE_PHC981_U_dsdc_n329 (.Z(FE_PHN981_U_dsdc_n329), 
	.A(U_dsdc_n329));
   BUF_X32 FE_PHC980_cr_reg_data_out_16_ (.Z(FE_PHN980_cr_reg_data_out_16_), 
	.A(cr_reg_data_out[16]));
   BUF_X32 FE_PHC979_cr_reg_data_out_30_ (.Z(FE_PHN979_cr_reg_data_out_30_), 
	.A(cr_reg_data_out[30]));
   BUF_X32 FE_PHC978_U_cr_N416 (.Z(FE_PHN978_U_cr_N416), 
	.A(U_cr_N416));
   BUF_X32 FE_PHC977_U_cr_N417 (.Z(FE_PHN977_U_cr_N417), 
	.A(U_cr_N417));
   BUF_X32 FE_PHC971_U_dsdc_init_cnt_5_ (.Z(FE_PHN971_U_dsdc_init_cnt_5_), 
	.A(U_dsdc_init_cnt_5_));
   BUF_X32 FE_PHC970_U_dsdc_init_cnt_11_ (.Z(FE_PHN970_U_dsdc_init_cnt_11_), 
	.A(U_dsdc_init_cnt_11_));
   BUF_X32 FE_PHC969_U_dsdc_n1727 (.Z(FE_PHN969_U_dsdc_n1727), 
	.A(U_dsdc_n1727));
   BUF_X16 FE_PHC968_U_dsdc_n415 (.Z(FE_PHN968_U_dsdc_n415), 
	.A(U_dsdc_n415));
   BUF_X32 FE_PHC967_U_dmc_n4 (.Z(FE_PHN967_U_dmc_n4), 
	.A(U_dmc_n4));
   BUF_X16 FE_PHC966_U_dsdc_n416 (.Z(FE_PHN966_U_dsdc_n416), 
	.A(U_dsdc_n416));
   BUF_X32 FE_PHC964_U_dsdc_n431 (.Z(FE_PHN964_U_dsdc_n431), 
	.A(FE_PHN3080_U_dsdc_n431));
   BUF_X16 FE_PHC961_U_dsdc_n231 (.Z(FE_PHN961_U_dsdc_n231), 
	.A(U_dsdc_n231));
   BUF_X32 FE_PHC960_U_dsdc_rcar_cnt2_nxt_3_ (.Z(FE_PHN960_U_dsdc_rcar_cnt2_nxt_3_), 
	.A(FE_PHN3079_U_dsdc_rcar_cnt2_nxt_3_));
   BUF_X32 FE_PHC959_U_dsdc_n226 (.Z(FE_PHN959_U_dsdc_n226), 
	.A(FE_PHN5144_U_dsdc_n226));
   BUF_X32 FE_PHC958_U_dsdc_n353 (.Z(FE_PHN958_U_dsdc_n353), 
	.A(U_dsdc_n353));
   BUF_X32 FE_PHC957_U_cr_N559 (.Z(FE_PHN957_U_cr_N559), 
	.A(FE_PHN5011_U_cr_N559));
   CLKBUF_X1 FE_PHC955_s_read_pipe_1_ (.Z(FE_PHN955_s_read_pipe_1_), 
	.A(s_read_pipe[1]));
   BUF_X32 FE_PHC953_U_dsdc_n375 (.Z(FE_PHN953_U_dsdc_n375), 
	.A(FE_PHN3222_U_dsdc_n375));
   BUF_X32 FE_PHC952_U_cr_N410 (.Z(FE_PHN952_U_cr_N410), 
	.A(FE_PHN3224_U_cr_N410));
   BUF_X32 FE_PHC951_U_dsdc_n216 (.Z(FE_PHN951_U_dsdc_n216), 
	.A(FE_PHN2975_U_dsdc_n216));
   BUF_X32 FE_PHC949_cr_reg_data_out_21_ (.Z(FE_PHN949_cr_reg_data_out_21_), 
	.A(cr_reg_data_out[21]));
   BUF_X32 FE_PHC948_U_cr_n442 (.Z(FE_PHN948_U_cr_n442), 
	.A(U_cr_n442));
   BUF_X32 FE_PHC945_U_dsdc_n1175 (.Z(FE_PHN945_U_dsdc_n1175), 
	.A(U_dsdc_n1175));
   CLKBUF_X1 FE_PHC944_U_dmc_n54 (.Z(FE_PHN944_U_dmc_n54), 
	.A(U_dmc_n54));
   BUF_X32 FE_PHC943_U_dmc_n7 (.Z(FE_PHN943_U_dmc_n7), 
	.A(U_dmc_n7));
   BUF_X32 FE_PHC942_U_dsdc_n408 (.Z(FE_PHN942_U_dsdc_n408), 
	.A(U_dsdc_n408));
   BUF_X32 FE_PHC940_U_dsdc_n294 (.Z(FE_PHN940_U_dsdc_n294), 
	.A(FE_PHN4582_U_dsdc_n294));
   BUF_X32 FE_PHC938_U_dsdc_n406 (.Z(FE_PHN938_U_dsdc_n406), 
	.A(FE_PHN3355_U_dsdc_n406));
   BUF_X32 FE_PHC937_U_dsdc_n297 (.Z(FE_PHN937_U_dsdc_n297), 
	.A(FE_PHN3115_U_dsdc_n297));
   BUF_X32 FE_PHC934_U_dsdc_n_2090_ (.Z(FE_PHN934_U_dsdc_n_2090_), 
	.A(U_dsdc_n[2090]));
   BUF_X32 FE_PHC933_U_dsdc_wtr_cnt_nxt_0_ (.Z(FE_PHN933_U_dsdc_wtr_cnt_nxt_0_), 
	.A(FE_PHN4395_U_dsdc_wtr_cnt_nxt_0_));
   BUF_X16 FE_PHC932_U_cr_N315 (.Z(FE_PHN932_U_cr_N315), 
	.A(U_cr_N315));
   BUF_X32 FE_PHC931_U_dsdc_n2094 (.Z(FE_PHN931_U_dsdc_n2094), 
	.A(U_dsdc_n2094));
   BUF_X8 FE_PHC927_U_addrdec_N108 (.Z(FE_PHN927_U_addrdec_N108), 
	.A(U_addrdec_N108));
   BUF_X16 FE_PHC926_U_cr_n98 (.Z(FE_PHN926_U_cr_n98), 
	.A(U_cr_n98));
   BUF_X32 FE_PHC925_U_dsdc_n410 (.Z(FE_PHN925_U_dsdc_n410), 
	.A(FE_PHN3452_U_dsdc_n410));
   BUF_X32 FE_PHC924_U_dsdc_rp_cnt2_nxt_2_ (.Z(FE_PHN924_U_dsdc_rp_cnt2_nxt_2_), 
	.A(FE_PHN3427_U_dsdc_rp_cnt2_nxt_2_));
   BUF_X32 FE_PHC922_U_dsdc_n412 (.Z(FE_PHN922_U_dsdc_n412), 
	.A(FE_PHN3399_U_dsdc_n412));
   BUF_X32 FE_PHC921_U_dsdc_N4461 (.Z(FE_PHN921_U_dsdc_N4461), 
	.A(U_dsdc_N4461));
   BUF_X32 FE_PHC918_cr_bank_addr_width_0_ (.Z(FE_PHN918_cr_bank_addr_width_0_), 
	.A(cr_bank_addr_width[0]));
   BUF_X32 FE_PHC917_U_dsdc_n223 (.Z(FE_PHN917_U_dsdc_n223), 
	.A(U_dsdc_n223));
   BUF_X32 FE_PHC916_U_cr_cr_cs_2_ (.Z(FE_PHN916_U_cr_cr_cs_2_), 
	.A(U_cr_cr_cs_2_));
   CLKBUF_X1 FE_PHC907_U_dsdc_cas_latency_1_ (.Z(FE_PHN907_U_dsdc_cas_latency_1_), 
	.A(U_dsdc_cas_latency_1_));
   BUF_X32 FE_PHC906_U_dsdc_n379 (.Z(FE_PHN906_U_dsdc_n379), 
	.A(FE_PHN3231_U_dsdc_n379));
   BUF_X32 FE_PHC905_U_dsdc_n374 (.Z(FE_PHN905_U_dsdc_n374), 
	.A(FE_PHN3166_U_dsdc_n374));
   BUF_X32 FE_PHC902_U_dmc_data_cnt_4_ (.Z(FE_PHN902_U_dmc_data_cnt_4_), 
	.A(U_dmc_data_cnt_4_));
   BUF_X32 FE_PHC901_U_dsdc_n295 (.Z(FE_PHN901_U_dsdc_n295), 
	.A(FE_PHN4603_U_dsdc_n295));
   BUF_X32 FE_PHC900_U_dsdc_rcar_cnt2_nxt_1_ (.Z(FE_PHN900_U_dsdc_rcar_cnt2_nxt_1_), 
	.A(U_dsdc_rcar_cnt2_nxt[1]));
   BUF_X32 FE_PHC899_U_dsdc_n227 (.Z(FE_PHN899_U_dsdc_n227), 
	.A(FE_PHN3244_U_dsdc_n227));
   BUF_X32 FE_PHC898_U_dsdc_n213 (.Z(FE_PHN898_U_dsdc_n213), 
	.A(FE_PHN4308_U_dsdc_n213));
   CLKBUF_X1 FE_PHC897_U_dsdc_n352 (.Z(FE_PHN897_U_dsdc_n352), 
	.A(U_dsdc_n352));
   BUF_X32 FE_PHC896_U_dsdc_n389 (.Z(FE_PHN896_U_dsdc_n389), 
	.A(FE_PHN4718_U_dsdc_n389));
   BUF_X32 FE_PHC895_U_dsdc_n283 (.Z(FE_PHN895_U_dsdc_n283), 
	.A(FE_PHN3297_U_dsdc_n283));
   BUF_X32 FE_PHC894_U_dsdc_n1464 (.Z(FE_PHN894_U_dsdc_n1464), 
	.A(U_dsdc_n1464));
   BUF_X32 FE_PHC893_U_dsdc_n1092 (.Z(FE_PHN893_U_dsdc_n1092), 
	.A(U_dsdc_n1092));
   BUF_X32 FE_PHC891_U_dsdc_wr_cnt_nxt_2_ (.Z(FE_PHN891_U_dsdc_wr_cnt_nxt_2_), 
	.A(FE_PHN3047_U_dsdc_wr_cnt_nxt_2_));
   BUF_X32 FE_PHC889_U_cr_N411 (.Z(FE_PHN889_U_cr_N411), 
	.A(U_cr_N411));
   BUF_X32 FE_PHC887_n4 (.Z(FE_PHN887_n4), 
	.A(FE_PHN3031_n4));
   BUF_X32 FE_PHC886_n6 (.Z(FE_PHN886_n6), 
	.A(FE_PHN3030_n6));
   BUF_X32 FE_PHC884_n1 (.Z(FE_PHN884_n1), 
	.A(n1));
   BUF_X32 FE_PHC883_n2 (.Z(FE_PHN883_n2), 
	.A(n2));
   BUF_X32 FE_PHC882_U_dsdc_n2097 (.Z(FE_PHN882_U_dsdc_n2097), 
	.A(U_dsdc_n2097));
   BUF_X32 FE_PHC881_n3 (.Z(FE_PHN881_n3), 
	.A(n3));
   BUF_X32 FE_PHC880_cr_reg_data_out_12_ (.Z(FE_PHN880_cr_reg_data_out_12_), 
	.A(cr_reg_data_out[12]));
   BUF_X16 FE_PHC866_U_dmc_n13 (.Z(FE_PHN866_U_dmc_n13), 
	.A(U_dmc_n13));
   BUF_X32 FE_PHC865_U_dsdc_n296 (.Z(FE_PHN865_U_dsdc_n296), 
	.A(FE_PHN3432_U_dsdc_n296));
   BUF_X32 FE_PHC864_U_dsdc_n222 (.Z(FE_PHN864_U_dsdc_n222), 
	.A(FE_PHN3320_U_dsdc_n222));
   BUF_X32 FE_PHC863_U_dsdc_n211 (.Z(FE_PHN863_U_dsdc_n211), 
	.A(FE_PHN3315_U_dsdc_n211));
   BUF_X32 FE_PHC862_U_dsdc_n230 (.Z(FE_PHN862_U_dsdc_n230), 
	.A(FE_PHN4962_U_dsdc_n230));
   BUF_X32 FE_PHC855_cr_reg_data_out_8_ (.Z(FE_PHN855_cr_reg_data_out_8_), 
	.A(cr_reg_data_out[8]));
   BUF_X32 FE_PHC854_U_dsdc_n2093 (.Z(FE_PHN854_U_dsdc_n2093), 
	.A(U_dsdc_n2093));
   BUF_X32 FE_PHC853_cr_reg_data_out_13_ (.Z(FE_PHN853_cr_reg_data_out_13_), 
	.A(cr_reg_data_out[13]));
   BUF_X32 FE_PHC850_cr_reg_data_out_7_ (.Z(FE_PHN850_cr_reg_data_out_7_), 
	.A(cr_reg_data_out[7]));
   CLKBUF_X1 FE_PHC843_U_dsdc_num_init_ref_cnt_1_ (.Z(FE_PHN843_U_dsdc_num_init_ref_cnt_1_), 
	.A(U_dsdc_num_init_ref_cnt_1_));
   BUF_X32 FE_PHC842_U_dsdc_n220 (.Z(FE_PHN842_U_dsdc_n220), 
	.A(U_dsdc_n220));
   BUF_X32 FE_PHC841_U_dsdc_bm_ras_cnt_max_3_ (.Z(FE_PHN841_U_dsdc_bm_ras_cnt_max_3_), 
	.A(U_dsdc_bm_ras_cnt_max_3_));
   BUF_X32 FE_PHC840_U_cr_n99 (.Z(FE_PHN840_U_cr_n99), 
	.A(FE_PHN3196_U_cr_n99));
   BUF_X32 FE_PHC838_U_dsdc_rp_cnt2_nxt_1_ (.Z(FE_PHN838_U_dsdc_rp_cnt2_nxt_1_), 
	.A(U_dsdc_rp_cnt2_nxt[1]));
   CLKBUF_X1 FE_PHC837_U_cr_cr_cs_0_ (.Z(FE_PHN837_U_cr_cr_cs_0_), 
	.A(U_cr_cr_cs_0_));
   BUF_X32 FE_PHC836_U_dsdc_n287 (.Z(FE_PHN836_U_dsdc_n287), 
	.A(U_dsdc_n287));
   BUF_X32 FE_PHC835_U_dsdc_term_cnt_nxt_4_ (.Z(FE_PHN835_U_dsdc_term_cnt_nxt_4_), 
	.A(FE_PHN3028_U_dsdc_term_cnt_nxt_4_));
   BUF_X32 FE_PHC834_U_dsdc_term_cnt_nxt_3_ (.Z(FE_PHN834_U_dsdc_term_cnt_nxt_3_), 
	.A(U_dsdc_term_cnt_nxt[3]));
   BUF_X32 FE_PHC833_U_dsdc_term_cnt_nxt_2_ (.Z(FE_PHN833_U_dsdc_term_cnt_nxt_2_), 
	.A(FE_PHN3011_U_dsdc_term_cnt_nxt_2_));
   BUF_X32 FE_PHC832_cr_reg_data_out_9_ (.Z(FE_PHN832_cr_reg_data_out_9_), 
	.A(cr_reg_data_out[9]));
   BUF_X32 FE_PHC831_cr_reg_data_out_6_ (.Z(FE_PHN831_cr_reg_data_out_6_), 
	.A(cr_reg_data_out[6]));
   BUF_X32 FE_PHC816_U_dsdc_n359 (.Z(FE_PHN816_U_dsdc_n359), 
	.A(U_dsdc_n359));
   BUF_X32 FE_PHC814_U_dsdc_n228 (.Z(FE_PHN814_U_dsdc_n228), 
	.A(FE_PHN5047_U_dsdc_n228));
   BUF_X32 FE_PHC807_U_cr_N420 (.Z(FE_PHN807_U_cr_N420), 
	.A(U_cr_N420));
   BUF_X32 FE_PHC800_U_cr_n96 (.Z(FE_PHN800_U_cr_n96), 
	.A(U_cr_n96));
   BUF_X32 FE_PHC799_U_dsdc_n225 (.Z(FE_PHN799_U_dsdc_n225), 
	.A(U_dsdc_n225));
   BUF_X32 FE_PHC797_U_dsdc_num_init_ref_cnt_nxt_1_ (.Z(FE_PHN797_U_dsdc_num_init_ref_cnt_nxt_1_), 
	.A(FE_PHN3324_U_dsdc_num_init_ref_cnt_nxt_1_));
   BUF_X32 FE_PHC796_U_dsdc_N4174 (.Z(FE_PHN796_U_dsdc_N4174), 
	.A(FE_PHN3104_U_dsdc_N4174));
   BUF_X16 FE_PHC792_U_dsdc_n219 (.Z(FE_PHN792_U_dsdc_n219), 
	.A(U_dsdc_n219));
   CLKBUF_X1 FE_PHC791_U_dsdc_n1491 (.Z(FE_PHN791_U_dsdc_n1491), 
	.A(U_dsdc_n1491));
   BUF_X32 FE_PHC790_U_dsdc_n289 (.Z(FE_PHN790_U_dsdc_n289), 
	.A(U_dsdc_n289));
   CLKBUF_X1 FE_PHC788_U_dsdc_n554 (.Z(FE_PHN788_U_dsdc_n554), 
	.A(U_dsdc_n554));
   BUF_X32 FE_PHC787_n90 (.Z(FE_PHN787_n90), 
	.A(n90));
   BUF_X32 FE_PHC786_U_dsdc_n291 (.Z(FE_PHN786_U_dsdc_n291), 
	.A(U_dsdc_n291));
   BUF_X16 FE_PHC781_U_dsdc_n224 (.Z(FE_PHN781_U_dsdc_n224), 
	.A(U_dsdc_n224));
   BUF_X32 FE_PHC777_U_dmc_N23 (.Z(FE_PHN777_U_dmc_N23), 
	.A(U_dmc_N23));
   BUF_X32 FE_PHC773_U_dsdc_n1823 (.Z(FE_PHN773_U_dsdc_n1823), 
	.A(U_dsdc_n1823));
   BUF_X32 FE_PHC772_U_dsdc_n2095 (.Z(FE_PHN772_U_dsdc_n2095), 
	.A(U_dsdc_n2095));
   CLKBUF_X1 FE_PHC771_U_dsdc_n1540 (.Z(FE_PHN771_U_dsdc_n1540), 
	.A(U_dsdc_n1540));
   BUF_X32 FE_PHC767_U_dsdc_term_cnt_nxt_1_ (.Z(FE_PHN767_U_dsdc_term_cnt_nxt_1_), 
	.A(U_dsdc_term_cnt_nxt[1]));
   BUF_X32 FE_PHC764_U_dsdc_n210 (.Z(FE_PHN764_U_dsdc_n210), 
	.A(U_dsdc_n210));
   BUF_X32 FE_PHC759_U_cr_N565 (.Z(FE_PHN759_U_cr_N565), 
	.A(U_cr_N565));
   BUF_X32 FE_PHC758_U_dsdc_n2096 (.Z(FE_PHN758_U_dsdc_n2096), 
	.A(FE_PHN3208_U_dsdc_n2096));
   BUF_X32 FE_PHC757_U_dsdc_auto_ref_en_nxt (.Z(FE_PHN757_U_dsdc_auto_ref_en_nxt), 
	.A(U_dsdc_auto_ref_en_nxt));
   BUF_X32 FE_PHC751_U_dsdc_rcar_cnt2_nxt_2_ (.Z(FE_PHN751_U_dsdc_rcar_cnt2_nxt_2_), 
	.A(U_dsdc_rcar_cnt2_nxt[2]));
   BUF_X32 FE_PHC745_U_dsdc_n229 (.Z(FE_PHN745_U_dsdc_n229), 
	.A(U_dsdc_n229));
   BUF_X32 FE_PHC742_U_dsdc_wtr_cnt_nxt_2_ (.Z(FE_PHN742_U_dsdc_wtr_cnt_nxt_2_), 
	.A(U_dsdc_wtr_cnt_nxt[2]));
   BUF_X32 FE_PHC740_U_dsdc_term_cnt_nxt_0_ (.Z(FE_PHN740_U_dsdc_term_cnt_nxt_0_), 
	.A(FE_PHN2941_U_dsdc_term_cnt_nxt_0_));
   BUF_X32 FE_PHC726_n7 (.Z(FE_PHN726_n7), 
	.A(n7));
   BUF_X32 FE_PHC725_cr_reg_data_out_10_ (.Z(FE_PHN725_cr_reg_data_out_10_), 
	.A(cr_reg_data_out[10]));
   BUF_X32 FE_PHC713_U_dmc_N24 (.Z(FE_PHN713_U_dmc_N24), 
	.A(U_dmc_N24));
   BUF_X32 FE_PHC710_cr_reg_data_out_3_ (.Z(FE_PHN710_cr_reg_data_out_3_), 
	.A(cr_reg_data_out[3]));
   BUF_X32 FE_PHC706_U_dsdc_n290 (.Z(FE_PHN706_U_dsdc_n290), 
	.A(U_dsdc_n290));
   BUF_X32 FE_PHC698_U_cr_N414 (.Z(FE_PHN698_U_cr_N414), 
	.A(U_cr_N414));
   BUF_X32 FE_PHC697_U_dsdc_n288 (.Z(FE_PHN697_U_dsdc_n288), 
	.A(U_dsdc_n288));
   BUF_X32 FE_PHC696_U_dsdc_n286 (.Z(FE_PHN696_U_dsdc_n286), 
	.A(U_dsdc_n286));
   BUF_X32 FE_PHC694_cr_reg_data_out_15_ (.Z(FE_PHN694_cr_reg_data_out_15_), 
	.A(cr_reg_data_out[15]));
   BUF_X32 FE_PHC691_n5 (.Z(FE_PHN691_n5), 
	.A(FE_PHN3029_n5));
   BUF_X16 FE_PHC683_U_dsdc_n1394 (.Z(FE_PHN683_U_dsdc_n1394), 
	.A(U_dsdc_n1394));
   BUF_X32 FE_PHC678_U_dsdc_n896 (.Z(FE_PHN678_U_dsdc_n896), 
	.A(U_dsdc_n896));
   BUF_X32 FE_PHC672_U_dsdc_n1436 (.Z(FE_PHN672_U_dsdc_n1436), 
	.A(U_dsdc_n1436));
   CLKBUF_X1 FE_PHC671_U_dsdc_n1637 (.Z(FE_PHN671_U_dsdc_n1637), 
	.A(FE_PHN5176_U_dsdc_n1637));
   BUF_X4 FE_OFC371_cr_t_ras_min_3_ (.Z(FE_OFN371_cr_t_ras_min_3_), 
	.A(cr_t_ras_min[3]));
   BUF_X4 FE_OFC365_n95 (.Z(FE_OFN365_n95), 
	.A(n95));
   BUF_X4 FE_OFC360_U_addrdec_n26 (.Z(FE_OFN360_U_addrdec_n26), 
	.A(U_addrdec_n26));
   BUF_X4 FE_OFC357_U_addrdec_n40 (.Z(FE_OFN357_U_addrdec_n40), 
	.A(U_addrdec_n40));
   BUF_X4 FE_OFC353_U_addrdec_n272 (.Z(FE_OFN353_U_addrdec_n272), 
	.A(U_addrdec_n272));
   BUF_X4 FE_OFC348_U_cr_n169 (.Z(FE_OFN348_U_cr_n169), 
	.A(U_cr_n169));
   BUF_X4 FE_OFC347_U_cr_n290 (.Z(FE_OFN347_U_cr_n290), 
	.A(U_cr_n290));
   BUF_X4 FE_OFC345_U_cr_n291 (.Z(FE_OFN345_U_cr_n291), 
	.A(U_cr_n291));
   BUF_X4 FE_OFC336_U_cr_n527 (.Z(FE_OFN336_U_cr_n527), 
	.A(U_cr_n527));
   BUF_X4 FE_OFC333_U_cr_n528 (.Z(FE_OFN333_U_cr_n528), 
	.A(U_cr_n528));
   BUF_X4 FE_OFC332_U_cr_n529 (.Z(FE_OFN332_U_cr_n529), 
	.A(U_cr_n529));
   BUF_X4 FE_OFC326_U_cr_n531 (.Z(FE_OFN326_U_cr_n531), 
	.A(U_cr_n531));
   BUF_X4 FE_OFC319_U_cr_n548 (.Z(FE_OFN319_U_cr_n548), 
	.A(U_cr_n548));
   BUF_X4 FE_OFC316_U_dsdc_n310 (.Z(FE_OFN316_U_dsdc_n310), 
	.A(U_dsdc_n310));
   BUF_X4 FE_OFC314_U_dsdc_n313 (.Z(FE_OFN314_U_dsdc_n313), 
	.A(U_dsdc_n313));
   BUF_X4 FE_OFC311_U_dsdc_n620 (.Z(FE_OFN311_U_dsdc_n620), 
	.A(U_dsdc_n620));
   BUF_X4 FE_OFC304_U_dsdc_n2014 (.Z(FE_OFN304_U_dsdc_n2014), 
	.A(U_dsdc_n2014));
   BUF_X4 FE_OFC303_U_dsdc_n2038 (.Z(FE_OFN303_U_dsdc_n2038), 
	.A(U_dsdc_n2038));
   BUF_X4 FE_OFC227_hiu_data_25_ (.Z(FE_OFN227_hiu_data_25_), 
	.A(hiu_wr_data[25]));
   BUF_X4 FE_OFC226_hiu_data_26_ (.Z(FE_OFN226_hiu_data_26_), 
	.A(hiu_wr_data[26]));
   BUF_X4 FE_OFC224_hiu_data_29_ (.Z(FE_OFN224_hiu_data_29_), 
	.A(hiu_wr_data[29]));
   BUF_X4 FE_OFC223_hiu_data_30_ (.Z(FE_OFN223_hiu_data_30_), 
	.A(hiu_wr_data[30]));
   BUF_X4 FE_OFC221_hiu_burst_size_0_ (.Z(FE_OFN221_hiu_burst_size_0_), 
	.A(hiu_burst_size[0]));
   BUF_X4 FE_OFC218_hiu_burst_size_2_ (.Z(FE_OFN218_hiu_burst_size_2_), 
	.A(hiu_burst_size[2]));
   BUF_X4 FE_OFC215_hiu_burst_size_4_ (.Z(FE_OFN215_hiu_burst_size_4_), 
	.A(hiu_burst_size[4]));
   BUF_X4 FE_OFC211_debug_ad_col_addr_13_ (.Z(FE_OFN211_debug_ad_col_addr_13_), 
	.A(debug_ad_col_addr_13__BAR_BAR));
   BUF_X4 FE_OFC189_HRESETn (.Z(FE_OFN189_HRESETn), 
	.A(FE_OFN36_HRESETn));
   BUF_X4 FE_OFC188_HRESETn (.Z(FE_OFN188_HRESETn), 
	.A(FE_OFN36_HRESETn));
   BUF_X4 FE_OFC187_HRESETn (.Z(FE_OFN187_HRESETn), 
	.A(FE_OFN36_HRESETn));
   BUF_X4 FE_OFC186_HRESETn (.Z(FE_OFN186_HRESETn), 
	.A(FE_OFN36_HRESETn));
   BUF_X4 FE_OFC183_HRESETn (.Z(FE_OFN183_HRESETn), 
	.A(FE_OFN39_HRESETn));
   BUF_X4 FE_OFC173_HRESETn (.Z(FE_OFN173_HRESETn), 
	.A(FE_OFN45_HRESETn));
   BUF_X4 FE_OFC172_HRESETn (.Z(FE_OFN172_HRESETn), 
	.A(FE_OFN46_HRESETn));
   BUF_X4 FE_OFC148_HRESETn (.Z(FE_OFN148_HRESETn), 
	.A(FE_OFN59_HRESETn));
   BUF_X4 FE_OFC142_HRESETn (.Z(FE_OFN142_HRESETn), 
	.A(FE_OFN63_HRESETn));
   BUF_X4 FE_OFC141_HRESETn (.Z(FE_OFN141_HRESETn), 
	.A(FE_OFN64_HRESETn));
   BUF_X8 FE_OFC64_HRESETn (.Z(FE_OFN64_HRESETn), 
	.A(FE_OFN39_HRESETn));
   BUF_X8 FE_OFC63_HRESETn (.Z(FE_OFN63_HRESETn), 
	.A(FE_OFN39_HRESETn));
   CLKBUF_X3 FE_OFC59_HRESETn (.Z(FE_OFN59_HRESETn), 
	.A(FE_OFN39_HRESETn));
   CLKBUF_X3 FE_OFC50_HRESETn (.Z(FE_OFN50_HRESETn), 
	.A(FE_OFN36_HRESETn));
   INV_X8 FE_OFC45_HRESETn (.ZN(FE_OFN45_HRESETn), 
	.A(hresetn));
   INV_X8 FE_OFC44_HRESETn (.ZN(FE_OFN44_HRESETn), 
	.A(hresetn));
   INV_X8 FE_OFC39_HRESETn (.ZN(FE_OFN39_HRESETn), 
	.A(hresetn));
   INV_X8 FE_OFC36_HRESETn (.ZN(FE_OFN36_HRESETn), 
	.A(hresetn));
   CLKBUF_X3 FE_OFC25_ctl_push_n (.Z(FE_OFN25_ctl_push_n), 
	.A(ctl_push_n));
   CLKBUF_X3 FE_OFC23_U_cr_n64 (.Z(FE_OFN23_U_cr_n64), 
	.A(U_cr_n64));
   CLKBUF_X3 FE_OFC1_U_cr_n541 (.Z(FE_OFN1_U_cr_n541), 
	.A(U_cr_n541));
   CLKBUF_X3 FE_OFC0_U_cr_n314 (.Z(FE_OFN0_U_cr_n314), 
	.A(U_cr_n314));
   DFFS_X2 cr_push_reg_n_reg (.SN(FE_OFN31_HRESETn), 
	.Q(cr_push_reg_n), 
	.D(FE_PHN3075_cr_push_n), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_31_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[31]), 
	.D(cr_reg_data_out[31]), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_30_ (.RN(FE_OFN28_HRESETn), 
	.Q(miu_rd_data_reg[30]), 
	.D(FE_PHN979_cr_reg_data_out_30_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_29_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[29]), 
	.D(FE_PHN1166_cr_reg_data_out_29_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_28_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[28]), 
	.D(FE_PHN1042_cr_reg_data_out_28_), 
	.CK(HCLK__L5_N6));
   DFFR_X1 miu_rd_data_reg_reg_27_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[27]), 
	.D(cr_reg_data_out[27]), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_26_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[26]), 
	.D(FE_PHN1372_cr_reg_data_out_26_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_25_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[25]), 
	.D(FE_PHN1236_cr_reg_data_out_25_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_24_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[24]), 
	.D(FE_PHN1169_cr_reg_data_out_24_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_23_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[23]), 
	.D(FE_PHN1369_cr_reg_data_out_23_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_22_ (.RN(FE_OFN28_HRESETn), 
	.Q(miu_rd_data_reg[22]), 
	.D(FE_PHN1077_cr_reg_data_out_22_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_21_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[21]), 
	.D(FE_PHN949_cr_reg_data_out_21_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_20_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[20]), 
	.D(FE_PHN1117_cr_reg_data_out_20_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_19_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[19]), 
	.D(FE_PHN1371_cr_reg_data_out_19_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_18_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[18]), 
	.D(FE_PHN1608_cr_reg_data_out_18_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_17_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[17]), 
	.D(FE_PHN1427_cr_reg_data_out_17_), 
	.CK(HCLK__L5_N6));
   DFFR_X1 miu_rd_data_reg_reg_16_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[16]), 
	.D(FE_PHN980_cr_reg_data_out_16_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_15_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[15]), 
	.D(FE_PHN2929_cr_reg_data_out_15_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_14_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[14]), 
	.D(FE_PHN1165_cr_reg_data_out_14_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_13_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[13]), 
	.D(FE_PHN853_cr_reg_data_out_13_), 
	.CK(HCLK__L5_N6));
   DFFR_X1 miu_rd_data_reg_reg_12_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[12]), 
	.D(FE_PHN880_cr_reg_data_out_12_), 
	.CK(HCLK__L5_N6));
   DFFR_X1 miu_rd_data_reg_reg_11_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[11]), 
	.D(FE_PHN1230_cr_reg_data_out_11_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_10_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[10]), 
	.D(FE_PHN725_cr_reg_data_out_10_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_9_ (.RN(FE_OFN28_HRESETn), 
	.Q(miu_rd_data_reg[9]), 
	.D(FE_PHN832_cr_reg_data_out_9_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_8_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[8]), 
	.D(FE_PHN855_cr_reg_data_out_8_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_7_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[7]), 
	.D(FE_PHN850_cr_reg_data_out_7_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_6_ (.RN(FE_OFN28_HRESETn), 
	.Q(miu_rd_data_reg[6]), 
	.D(FE_PHN831_cr_reg_data_out_6_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_5_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[5]), 
	.D(FE_PHN1235_cr_reg_data_out_5_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_4_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[4]), 
	.D(FE_PHN1234_cr_reg_data_out_4_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_3_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[3]), 
	.D(FE_PHN710_cr_reg_data_out_3_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_2_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[2]), 
	.D(FE_PHN1041_cr_reg_data_out_2_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_1_ (.RN(FE_OFN160_HRESETn), 
	.Q(miu_rd_data_reg[1]), 
	.D(FE_PHN1167_cr_reg_data_out_1_), 
	.CK(HCLK__L5_N17));
   DFFR_X1 miu_rd_data_reg_reg_0_ (.RN(FE_OFN51_HRESETn), 
	.Q(miu_rd_data_reg[0]), 
	.D(FE_PHN1080_cr_reg_data_out_0_), 
	.CK(HCLK__L5_N17));
   AOI22_X1 U3 (.ZN(n1), 
	.B2(miu_rd_data_reg[2]), 
	.B1(FE_OFN25_ctl_push_n), 
	.A2(n82), 
	.A1(s_rd_data[2]));
   INV_X1 U4 (.ZN(miu_rd_data_out[2]), 
	.A(FE_PHN884_n1));
   AOI22_X1 U5 (.ZN(n2), 
	.B2(miu_rd_data_reg[8]), 
	.B1(FE_OFN25_ctl_push_n), 
	.A2(n82), 
	.A1(s_rd_data[8]));
   INV_X1 U6 (.ZN(miu_rd_data_out[8]), 
	.A(FE_PHN883_n2));
   AOI22_X1 U7 (.ZN(n3), 
	.B2(miu_rd_data_reg[4]), 
	.B1(FE_OFN25_ctl_push_n), 
	.A2(n82), 
	.A1(s_rd_data[4]));
   INV_X1 U8 (.ZN(miu_rd_data_out[4]), 
	.A(FE_PHN881_n3));
   AOI22_X1 U9 (.ZN(n4), 
	.B2(miu_rd_data_reg[11]), 
	.B1(FE_OFN25_ctl_push_n), 
	.A2(n82), 
	.A1(s_rd_data[11]));
   INV_X1 U10 (.ZN(miu_rd_data_out[11]), 
	.A(FE_PHN887_n4));
   AOI22_X1 U11 (.ZN(n5), 
	.B2(miu_rd_data_reg[14]), 
	.B1(FE_OFN25_ctl_push_n), 
	.A2(n82), 
	.A1(s_rd_data[14]));
   INV_X1 U12 (.ZN(miu_rd_data_out[14]), 
	.A(FE_PHN691_n5));
   AOI22_X1 U13 (.ZN(n6), 
	.B2(miu_rd_data_reg[13]), 
	.B1(FE_OFN25_ctl_push_n), 
	.A2(n82), 
	.A1(s_rd_data[13]));
   INV_X1 U14 (.ZN(miu_rd_data_out[13]), 
	.A(FE_PHN886_n6));
   AOI22_X1 U15 (.ZN(n7), 
	.B2(miu_rd_data_reg[15]), 
	.B1(FE_OFN25_ctl_push_n), 
	.A2(n82), 
	.A1(s_rd_data[15]));
   INV_X1 U16 (.ZN(miu_rd_data_out[15]), 
	.A(FE_PHN726_n7));
   AND3_X4 U18 (.ZN(miu_push_n), 
	.A3(FE_OFN25_ctl_push_n), 
	.A2(cr_push_reg_n), 
	.A1(dmc_push_n));
   NAND2_X1 U20 (.ZN(n19), 
	.A2(hiu_mem_req), 
	.A1(n21));
   INV_X1 U21 (.ZN(n21), 
	.A(sdram_req_i));
   OAI22_X2 U25 (.ZN(N28), 
	.B2(n19), 
	.B1(ad_static_mem_req), 
	.A2(U_cr_n39), 
	.A1(n21));
   INV_X4 U26 (.ZN(n14), 
	.A(n44));
   MUX2_X2 U29 (.Z(miu_rd_data_out[22]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[22]), 
	.A(s_rd_data[22]));
   MUX2_X2 U30 (.Z(miu_rd_data_out[30]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[30]), 
	.A(s_rd_data[30]));
   MUX2_X2 U31 (.Z(miu_rd_data_out[20]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[20]), 
	.A(s_rd_data[20]));
   MUX2_X2 U32 (.Z(miu_rd_data_out[31]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[31]), 
	.A(s_rd_data[31]));
   MUX2_X2 U33 (.Z(miu_rd_data_out[24]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[24]), 
	.A(s_rd_data[24]));
   MUX2_X2 U34 (.Z(miu_rd_data_out[28]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[28]), 
	.A(s_rd_data[28]));
   MUX2_X2 U35 (.Z(miu_rd_data_out[27]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[27]), 
	.A(s_rd_data[27]));
   MUX2_X2 U36 (.Z(miu_rd_data_out[18]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[18]), 
	.A(s_rd_data[18]));
   MUX2_X2 U37 (.Z(miu_rd_data_out[16]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[16]), 
	.A(s_rd_data[16]));
   MUX2_X2 U38 (.Z(miu_rd_data_out[23]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[23]), 
	.A(s_rd_data[23]));
   MUX2_X2 U39 (.Z(miu_rd_data_out[21]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[21]), 
	.A(s_rd_data[21]));
   MUX2_X2 U40 (.Z(miu_rd_data_out[19]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[19]), 
	.A(s_rd_data[19]));
   MUX2_X2 U41 (.Z(miu_rd_data_out[17]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[17]), 
	.A(s_rd_data[17]));
   MUX2_X2 U42 (.Z(miu_rd_data_out[25]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[25]), 
	.A(s_rd_data[25]));
   MUX2_X2 U43 (.Z(miu_rd_data_out[26]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[26]), 
	.A(s_rd_data[26]));
   MUX2_X2 U44 (.Z(miu_rd_data_out[29]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[29]), 
	.A(s_rd_data[29]));
   AND3_X4 U45 (.ZN(miu_pop_n), 
	.A3(dmc_pop_n), 
	.A2(ctl_pop_n), 
	.A1(cr_pop_n));
   MUX2_X2 U48 (.Z(miu_rd_data_out[0]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[0]), 
	.A(s_rd_data[0]));
   MUX2_X2 U49 (.Z(miu_rd_data_out[10]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[10]), 
	.A(s_rd_data[10]));
   MUX2_X2 U50 (.Z(miu_rd_data_out[12]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[12]), 
	.A(s_rd_data[12]));
   MUX2_X2 U51 (.Z(miu_rd_data_out[1]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[1]), 
	.A(s_rd_data[1]));
   MUX2_X2 U52 (.Z(miu_rd_data_out[3]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[3]), 
	.A(s_rd_data[3]));
   MUX2_X2 U53 (.Z(miu_rd_data_out[5]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[5]), 
	.A(s_rd_data[5]));
   MUX2_X2 U54 (.Z(miu_rd_data_out[6]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[6]), 
	.A(s_rd_data[6]));
   MUX2_X2 U55 (.Z(miu_rd_data_out[7]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[7]), 
	.A(s_rd_data[7]));
   MUX2_X2 U56 (.Z(miu_rd_data_out[9]), 
	.S(FE_OFN25_ctl_push_n), 
	.B(miu_rd_data_reg[9]), 
	.A(s_rd_data[9]));
   OAI211_X1 U_dsdc_U2200 (.ZN(U_dsdc_n1673), 
	.C2(U_dsdc_n482), 
	.C1(U_dsdc_init_cnt_14_), 
	.B(U_dsdc_n1676), 
	.A(U_dsdc_init_cnt_15_));
   OAI211_X1 U_dsdc_U2198 (.ZN(U_dsdc_n1559), 
	.C2(FE_PHN1887_U_dsdc_n166), 
	.C1(U_dsdc_r_wrapped_burst), 
	.B(U_dsdc_n299), 
	.A(U_dsdc_r_burst_size_0_));
   NOR4_X1 U_dsdc_U2197 (.ZN(U_dsdc_n1479), 
	.A4(U_dsdc_n1506), 
	.A3(U_dsdc_n341), 
	.A2(U_dsdc_n432), 
	.A1(U_dsdc_operation_cs_3_));
   AOI21_X1 U_dsdc_U2196 (.ZN(U_dsdc_n1486), 
	.B2(U_dsdc_n1522), 
	.B1(U_dsdc_n1450), 
	.A(U_dsdc_n432));
   XNOR2_X2 U_dsdc_U2195 (.ZN(U_dsdc_n1306), 
	.B(cr_t_wr[0]), 
	.A(cr_t_wr[1]));
   XOR2_X2 U_dsdc_U2194 (.Z(U_dsdc_n1277), 
	.B(U_dsdc_n1278), 
	.A(FE_PHN1343_U_dsdc_n1276));
   XOR2_X2 U_dsdc_U2193 (.Z(U_dsdc_n1271), 
	.B(U_dsdc_n1267), 
	.A(U_dsdc_n1272));
   XNOR2_X2 U_dsdc_U2192 (.ZN(U_dsdc_n1247), 
	.B(cr_t_wtr[0]), 
	.A(cr_t_wtr[1]));
   MUX2_X2 U_dsdc_U2191 (.Z(U_dsdc_N4463), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_n1245), 
	.A(cr_t_ras_min[3]));
   MUX2_X2 U_dsdc_U2190 (.Z(U_dsdc_N4476), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_n1235), 
	.A(cr_t_rc[3]));
   MUX2_X2 U_dsdc_U2189 (.Z(U_dsdc_N4477), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__0_), 
	.A(U_dsdc_n1225));
   MUX2_X2 U_dsdc_U2188 (.Z(U_dsdc_N4478), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__1_), 
	.A(U_dsdc_n1224));
   MUX2_X2 U_dsdc_U2187 (.Z(U_dsdc_N4479), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__2_), 
	.A(U_dsdc_n1223));
   MUX2_X2 U_dsdc_U2186 (.Z(U_dsdc_N4480), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__3_), 
	.A(U_dsdc_n1222));
   MUX2_X2 U_dsdc_U2185 (.Z(U_dsdc_N4481), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__4_), 
	.A(U_dsdc_n1221));
   MUX2_X2 U_dsdc_U2184 (.Z(U_dsdc_N4482), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__5_), 
	.A(U_dsdc_n1220));
   MUX2_X2 U_dsdc_U2183 (.Z(U_dsdc_N4483), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__6_), 
	.A(U_dsdc_n1219));
   MUX2_X2 U_dsdc_U2182 (.Z(U_dsdc_N4490), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__13_), 
	.A(U_dsdc_n1218));
   MUX2_X2 U_dsdc_U2181 (.Z(U_dsdc_N4491), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__14_), 
	.A(U_dsdc_n1217));
   MUX2_X2 U_dsdc_U2180 (.Z(U_dsdc_N4492), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__15_), 
	.A(U_dsdc_n1216));
   MUX2_X2 U_dsdc_U2179 (.Z(U_dsdc_N4416), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_n1215), 
	.A(cr_t_ras_min[3]));
   MUX2_X2 U_dsdc_U2178 (.Z(U_dsdc_N4429), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_n1208), 
	.A(cr_t_rc[3]));
   MUX2_X2 U_dsdc_U2177 (.Z(U_dsdc_N4430), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__0_), 
	.A(U_dsdc_n1225));
   MUX2_X2 U_dsdc_U2176 (.Z(U_dsdc_N4431), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__1_), 
	.A(U_dsdc_n1224));
   MUX2_X2 U_dsdc_U2175 (.Z(U_dsdc_N4432), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__2_), 
	.A(U_dsdc_n1223));
   MUX2_X2 U_dsdc_U2174 (.Z(U_dsdc_N4433), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__3_), 
	.A(U_dsdc_n1222));
   MUX2_X2 U_dsdc_U2173 (.Z(U_dsdc_N4434), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__4_), 
	.A(U_dsdc_n1221));
   MUX2_X2 U_dsdc_U2172 (.Z(U_dsdc_N4435), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__5_), 
	.A(U_dsdc_n1220));
   MUX2_X2 U_dsdc_U2171 (.Z(U_dsdc_N4436), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__6_), 
	.A(U_dsdc_n1219));
   MUX2_X2 U_dsdc_U2170 (.Z(U_dsdc_N4443), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__13_), 
	.A(U_dsdc_n1218));
   MUX2_X2 U_dsdc_U2169 (.Z(U_dsdc_N4444), 
	.S(FE_OFN316_U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__14_), 
	.A(U_dsdc_n1217));
   MUX2_X2 U_dsdc_U2168 (.Z(U_dsdc_N4445), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__15_), 
	.A(U_dsdc_n1216));
   MUX2_X2 U_dsdc_U2167 (.Z(U_dsdc_N4369), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_n1201), 
	.A(cr_t_ras_min[3]));
   MUX2_X2 U_dsdc_U2166 (.Z(U_dsdc_N4382), 
	.S(U_dsdc_n620), 
	.B(FE_PHN1487_U_dsdc_n1194), 
	.A(cr_t_rc[3]));
   MUX2_X2 U_dsdc_U2165 (.Z(U_dsdc_N4383), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__0_), 
	.A(U_dsdc_n1225));
   MUX2_X2 U_dsdc_U2164 (.Z(U_dsdc_N4384), 
	.S(FE_OFN311_U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__1_), 
	.A(U_dsdc_n1224));
   MUX2_X2 U_dsdc_U2163 (.Z(U_dsdc_N4385), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__2_), 
	.A(U_dsdc_n1223));
   MUX2_X2 U_dsdc_U2162 (.Z(U_dsdc_N4386), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__3_), 
	.A(U_dsdc_n1222));
   MUX2_X2 U_dsdc_U2161 (.Z(U_dsdc_N4387), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__4_), 
	.A(U_dsdc_n1221));
   MUX2_X2 U_dsdc_U2160 (.Z(U_dsdc_N4388), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__5_), 
	.A(U_dsdc_n1220));
   MUX2_X2 U_dsdc_U2159 (.Z(U_dsdc_N4389), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__6_), 
	.A(U_dsdc_n1219));
   MUX2_X2 U_dsdc_U2158 (.Z(U_dsdc_N4396), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__13_), 
	.A(U_dsdc_n1218));
   MUX2_X2 U_dsdc_U2157 (.Z(U_dsdc_N4397), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__14_), 
	.A(U_dsdc_n1217));
   MUX2_X2 U_dsdc_U2156 (.Z(U_dsdc_N4398), 
	.S(FE_OFN311_U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__15_), 
	.A(U_dsdc_n1216));
   MUX2_X2 U_dsdc_U2155 (.Z(U_dsdc_N4322), 
	.S(n83), 
	.B(U_dsdc_n1187), 
	.A(FE_OFN371_cr_t_ras_min_3_));
   MUX2_X2 U_dsdc_U2154 (.Z(U_dsdc_N4335), 
	.S(n83), 
	.B(FE_PHN1492_U_dsdc_n1180), 
	.A(cr_t_rc[3]));
   MUX2_X2 U_dsdc_U2152 (.Z(U_dsdc_N4336), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__0_), 
	.A(U_dsdc_n1225));
   MUX2_X2 U_dsdc_U2151 (.Z(U_dsdc_N4337), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__1_), 
	.A(U_dsdc_n1224));
   MUX2_X2 U_dsdc_U2150 (.Z(U_dsdc_N4338), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__2_), 
	.A(U_dsdc_n1223));
   MUX2_X2 U_dsdc_U2149 (.Z(U_dsdc_N4339), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__3_), 
	.A(U_dsdc_n1222));
   MUX2_X2 U_dsdc_U2148 (.Z(U_dsdc_N4340), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__4_), 
	.A(U_dsdc_n1221));
   MUX2_X2 U_dsdc_U2147 (.Z(U_dsdc_N4341), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__5_), 
	.A(U_dsdc_n1220));
   MUX2_X2 U_dsdc_U2146 (.Z(U_dsdc_N4342), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__6_), 
	.A(U_dsdc_n1219));
   MUX2_X2 U_dsdc_U2145 (.Z(U_dsdc_N4349), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__13_), 
	.A(U_dsdc_n1218));
   MUX2_X2 U_dsdc_U2144 (.Z(U_dsdc_N4350), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__14_), 
	.A(U_dsdc_n1217));
   MUX2_X2 U_dsdc_U2143 (.Z(U_dsdc_N4351), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__15_), 
	.A(U_dsdc_n1216));
   MUX2_X2 U_dsdc_U2142 (.Z(U_dsdc_N4139), 
	.S(U_dsdc_n1166), 
	.B(cr_t_rcd[0]), 
	.A(U_dsdc_n1164));
   MUX2_X2 U_dsdc_U2141 (.Z(U_dsdc_N4140), 
	.S(U_dsdc_n1166), 
	.B(cr_t_rcd[1]), 
	.A(U_dsdc_n1162));
   MUX2_X2 U_dsdc_U2140 (.Z(U_dsdc_n1157), 
	.S(U_dsdc_n1166), 
	.B(U_cr_n120), 
	.A(U_dsdc_n1156));
   MUX2_X2 U_dsdc_U2139 (.Z(U_dsdc_n1155), 
	.S(U_dsdc_n1166), 
	.B(FE_PHN3192_U_cr_n128), 
	.A(U_dsdc_n1154));
   MUX2_X2 U_dsdc_U2137 (.Z(U_dsdc_N4484), 
	.S(FE_OFN314_U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__7_), 
	.A(U_dsdc_n1151));
   MUX2_X2 U_dsdc_U2136 (.Z(U_dsdc_N4437), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__7_), 
	.A(U_dsdc_n1151));
   MUX2_X2 U_dsdc_U2135 (.Z(U_dsdc_N4390), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__7_), 
	.A(U_dsdc_n1151));
   MUX2_X2 U_dsdc_U2134 (.Z(U_dsdc_N4343), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__7_), 
	.A(U_dsdc_n1151));
   MUX2_X2 U_dsdc_U2133 (.Z(U_dsdc_N4485), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__8_), 
	.A(U_dsdc_n1149));
   MUX2_X2 U_dsdc_U2132 (.Z(U_dsdc_N4438), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__8_), 
	.A(U_dsdc_n1149));
   MUX2_X2 U_dsdc_U2131 (.Z(U_dsdc_N4391), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__8_), 
	.A(U_dsdc_n1149));
   MUX2_X2 U_dsdc_U2130 (.Z(U_dsdc_N4344), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__8_), 
	.A(U_dsdc_n1149));
   MUX2_X2 U_dsdc_U2129 (.Z(U_dsdc_N4486), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__9_), 
	.A(U_dsdc_n1148));
   MUX2_X2 U_dsdc_U2128 (.Z(U_dsdc_N4439), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__9_), 
	.A(U_dsdc_n1148));
   MUX2_X2 U_dsdc_U2127 (.Z(U_dsdc_N4392), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__9_), 
	.A(U_dsdc_n1148));
   MUX2_X2 U_dsdc_U2126 (.Z(U_dsdc_N4345), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__9_), 
	.A(U_dsdc_n1148));
   MUX2_X2 U_dsdc_U2125 (.Z(U_dsdc_N4487), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__10_), 
	.A(U_dsdc_n1146));
   MUX2_X2 U_dsdc_U2124 (.Z(U_dsdc_N4440), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__10_), 
	.A(U_dsdc_n1146));
   MUX2_X2 U_dsdc_U2123 (.Z(U_dsdc_N4393), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__10_), 
	.A(U_dsdc_n1146));
   MUX2_X2 U_dsdc_U2122 (.Z(U_dsdc_N4346), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__10_), 
	.A(U_dsdc_n1146));
   MUX2_X2 U_dsdc_U2121 (.Z(U_dsdc_N4488), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__11_), 
	.A(U_dsdc_n1145));
   MUX2_X2 U_dsdc_U2120 (.Z(U_dsdc_N4441), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__11_), 
	.A(U_dsdc_n1145));
   MUX2_X2 U_dsdc_U2119 (.Z(U_dsdc_N4394), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__11_), 
	.A(U_dsdc_n1145));
   MUX2_X2 U_dsdc_U2118 (.Z(U_dsdc_N4347), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__11_), 
	.A(U_dsdc_n1145));
   MUX2_X2 U_dsdc_U2117 (.Z(U_dsdc_N4489), 
	.S(U_dsdc_n313), 
	.B(U_dsdc_bm_row_addr_3__12_), 
	.A(U_dsdc_n1143));
   MUX2_X2 U_dsdc_U2116 (.Z(U_dsdc_N4442), 
	.S(U_dsdc_n310), 
	.B(U_dsdc_bm_row_addr_2__12_), 
	.A(U_dsdc_n1143));
   MUX2_X2 U_dsdc_U2115 (.Z(U_dsdc_N4395), 
	.S(U_dsdc_n620), 
	.B(U_dsdc_bm_row_addr_1__12_), 
	.A(U_dsdc_n1143));
   MUX2_X2 U_dsdc_U2114 (.Z(U_dsdc_N4348), 
	.S(n83), 
	.B(U_dsdc_bm_row_addr_0__12_), 
	.A(U_dsdc_n1143));
   XNOR2_X2 U_dsdc_U2113 (.ZN(U_dsdc_cas_latency_2_), 
	.B(FE_PHN1596_U_dsdc_n1091), 
	.A(U_dsdc_n1093));
   MUX2_X2 U_dsdc_U2111 (.Z(U_dsdc_n1023), 
	.S(U_dsdc_bm_num_open_bank_3_), 
	.B(U_dsdc_n1326), 
	.A(U_dsdc_n1166));
   MUX2_X2 U_dsdc_U2110 (.Z(U_dsdc_n1015), 
	.S(U_dsdc_bm_num_open_bank_2_), 
	.B(U_dsdc_n1290), 
	.A(U_dsdc_n1159));
   MUX2_X2 U_dsdc_U2109 (.Z(U_dsdc_n1010), 
	.S(U_dsdc_bm_num_open_bank_1_), 
	.B(U_dsdc_n1326), 
	.A(U_dsdc_n1166));
   MUX2_X2 U_dsdc_U2108 (.Z(U_dsdc_n1007), 
	.S(FE_PHN1093_U_dsdc_n340), 
	.B(U_dsdc_n1159), 
	.A(U_dsdc_n1290));
   XNOR2_X2 U_dsdc_U2107 (.ZN(U_dsdc_n827), 
	.B(U_dsdc_n361), 
	.A(ad_sdram_chip_select_0_));
   NAND2_X2 U_dsdc_U2101 (.ZN(U_dsdc_n1258), 
	.A2(U_dsdc_n1163), 
	.A1(U_dsdc_n1418));
   INV_X4 U_dsdc_U2100 (.ZN(U_dsdc_n1817), 
	.A(U_dsdc_n2041));
   NAND2_X2 U_dsdc_U2098 (.ZN(U_dsdc_n2013), 
	.A2(U_dsdc_n1411), 
	.A1(U_dsdc_n891));
   INV_X4 U_dsdc_U2097 (.ZN(U_dsdc_n759), 
	.A(U_dsdc_n1413));
   INV_X4 U_dsdc_U2096 (.ZN(U_dsdc_n1038), 
	.A(U_dsdc_n2014));
   INV_X4 U_dsdc_U2095 (.ZN(U_dsdc_n964), 
	.A(U_dsdc_n966));
   NOR2_X2 U_dsdc_U2093 (.ZN(U_dsdc_n1800), 
	.A2(U_dsdc_n1574), 
	.A1(U_dsdc_n1577));
   NOR2_X2 U_dsdc_U2092 (.ZN(U_dsdc_n604), 
	.A2(U_dsdc_n1127), 
	.A1(debug_ad_bank_addr[1]));
   OAI21_X1 U_dsdc_U2091 (.ZN(U_dsdc_n1005), 
	.B2(U_dsdc_n1166), 
	.B1(U_dsdc_n1326), 
	.A(FE_PHN1093_U_dsdc_n340));
   AOI221_X2 U_dsdc_U2090 (.ZN(U_dsdc_n1576), 
	.C2(U_dsdc_n2059), 
	.C1(U_cr_n39), 
	.B2(U_dsdc_n2059), 
	.B1(U_dsdc_n2066), 
	.A(U_dsdc_n1478));
   AOI222_X1 U_dsdc_U2088 (.ZN(U_dsdc_n749), 
	.C2(hiu_burst_size[3]), 
	.C1(U_dsdc_n983), 
	.B2(FE_PHN1892_U_dsdc_r_burst_size_3_), 
	.B1(U_dsdc_n751), 
	.A2(U_dsdc_data_cnt_3_), 
	.A1(U_dsdc_RSOP_1683_C2_CONTROL1));
   AOI222_X1 U_dsdc_U2087 (.ZN(U_dsdc_n747), 
	.C2(hiu_burst_size[5]), 
	.C1(U_dsdc_n983), 
	.B2(FE_PHN1890_U_dsdc_r_burst_size_5_), 
	.B1(U_dsdc_n751), 
	.A2(U_dsdc_data_cnt_5_), 
	.A1(U_dsdc_RSOP_1683_C2_CONTROL1));
   AOI21_X1 U_dsdc_U2085 (.ZN(U_dsdc_n1316), 
	.B2(U_dsdc_n1558), 
	.B1(U_dsdc_n1312), 
	.A(U_dsdc_n181));
   INV_X4 U_dsdc_U2084 (.ZN(U_dsdc_n1388), 
	.A(U_dsdc_n1112));
   XNOR2_X2 U_dsdc_U2083 (.ZN(U_dsdc_n566), 
	.B(debug_ad_row_addr[2]), 
	.A(U_dsdc_n565));
   XNOR2_X2 U_dsdc_U2082 (.ZN(U_dsdc_n567), 
	.B(U_dsdc_n561), 
	.A(debug_ad_row_addr[0]));
   XNOR2_X2 U_dsdc_U2081 (.ZN(U_dsdc_n568), 
	.B(debug_ad_row_addr[4]), 
	.A(U_dsdc_n557));
   XNOR2_X2 U_dsdc_U2080 (.ZN(U_dsdc_n549), 
	.B(debug_ad_row_addr[14]), 
	.A(U_dsdc_n548));
   XNOR2_X2 U_dsdc_U2079 (.ZN(U_dsdc_n550), 
	.B(debug_ad_row_addr[10]), 
	.A(U_dsdc_n546));
   XNOR2_X2 U_dsdc_U2078 (.ZN(U_dsdc_n539), 
	.B(U_addrdec_n241), 
	.A(U_dsdc_n519));
   XNOR2_X2 U_dsdc_U2077 (.ZN(U_dsdc_n511), 
	.B(debug_ad_row_addr[8]), 
	.A(U_dsdc_n510));
   XNOR2_X2 U_dsdc_U2076 (.ZN(U_dsdc_n512), 
	.B(debug_ad_row_addr[6]), 
	.A(U_dsdc_n504));
   OR2_X4 U_dsdc_U2075 (.ZN(U_dsdc_n399), 
	.A2(U_dsdc_n1661), 
	.A1(U_dsdc_n1660));
   AND2_X4 U_dsdc_U2074 (.ZN(U_dsdc_n360), 
	.A2(FE_PHN1887_U_dsdc_n166), 
	.A1(U_dsdc_n1425));
   OR2_X4 U_dsdc_U2073 (.ZN(U_dsdc_n346), 
	.A2(U_dsdc_n1655), 
	.A1(U_dsdc_n1658));
   OR2_X4 U_dsdc_U2072 (.ZN(U_dsdc_n345), 
	.A2(U_dsdc_n1655), 
	.A1(U_dsdc_n1660));
   AND2_X4 U_dsdc_U2071 (.ZN(U_dsdc_n330), 
	.A2(U_dsdc_bm_row_addr_2__2_), 
	.A1(U_dsdc_n159));
   AND2_X4 U_dsdc_U2070 (.ZN(U_dsdc_n314), 
	.A2(U_dsdc_bm_row_addr_0__8_), 
	.A1(U_dsdc_n998));
   AND2_X4 U_dsdc_U2069 (.ZN(U_dsdc_n312), 
	.A2(U_dsdc_bm_row_addr_0__10_), 
	.A1(U_dsdc_n998));
   AND2_X4 U_dsdc_U2067 (.ZN(U_dsdc_n305), 
	.A2(U_dsdc_n703), 
	.A1(U_dsdc_n1415));
   NAND2_X2 U_dsdc_U2066 (.ZN(U_dsdc_n599), 
	.A2(U_dsdc_n1127), 
	.A1(debug_ad_bank_addr[1]));
   AND2_X4 U_dsdc_U2064 (.ZN(U_dsdc_n184), 
	.A2(U_dsdc_n1258), 
	.A1(U_dsdc_n725));
   INV_X4 U_dsdc_U2062 (.ZN(U_dsdc_n983), 
	.A(U_dsdc_n1546));
   AND3_X4 U_dsdc_U2061 (.ZN(U_dsdc_n810), 
	.A3(U_dsdc_n789), 
	.A2(U_dsdc_n790), 
	.A1(U_dsdc_n791));
   AND3_X4 U_dsdc_U2060 (.ZN(U_dsdc_n802), 
	.A3(U_dsdc_n786), 
	.A2(U_dsdc_n787), 
	.A1(U_dsdc_n788));
   AND3_X4 U_dsdc_U2059 (.ZN(U_dsdc_n808), 
	.A3(U_dsdc_n792), 
	.A2(U_dsdc_n793), 
	.A1(U_dsdc_n794));
   AND3_X4 U_dsdc_U2058 (.ZN(U_dsdc_n805), 
	.A3(U_dsdc_n782), 
	.A2(U_dsdc_n783), 
	.A1(U_dsdc_n784));
   NOR2_X2 U_dsdc_U2057 (.ZN(U_dsdc_n1980), 
	.A2(U_dsdc_n354), 
	.A1(U_dsdc_n1447));
   NOR2_X2 U_dsdc_U2056 (.ZN(U_dsdc_n1364), 
	.A2(FE_PHN1887_U_dsdc_n166), 
	.A1(U_dsdc_n184));
   AND2_X4 U_dsdc_U2055 (.ZN(U_dsdc_n1840), 
	.A2(U_dsdc_r_close_bank_addr_1_), 
	.A1(U_dsdc_n292));
   INV_X4 U_dsdc_U2054 (.ZN(U_dsdc_n1309), 
	.A(U_dsdc_n1411));
   NOR2_X2 U_dsdc_U2053 (.ZN(U_dsdc_n1425), 
	.A2(U_dsdc_n667), 
	.A1(U_dsdc_n712));
   INV_X1 U_dsdc_U2052 (.ZN(U_dsdc_n1561), 
	.A(U_dsdc_n663));
   NOR2_X1 U_dsdc_U2051 (.ZN(U_dsdc_n691), 
	.A2(U_dsdc_n167), 
	.A1(U_dsdc_n1427));
   NOR2_X1 U_dsdc_U2050 (.ZN(U_dsdc_n866), 
	.A2(U_dsdc_n355), 
	.A1(U_dsdc_n692));
   AND4_X4 U_dsdc_U2049 (.ZN(U_dsdc_n886), 
	.A4(U_dsdc_n1438), 
	.A3(U_dsdc_n988), 
	.A2(sdram_req_i), 
	.A1(U_dsdc_n885));
   NOR2_X2 U_dsdc_U2048 (.ZN(U_dsdc_n1299), 
	.A2(U_dsdc_n165), 
	.A1(U_dsdc_n880));
   NOR2_X2 U_dsdc_U2047 (.ZN(U_dsdc_n1499), 
	.A2(U_dsdc_n1521), 
	.A1(U_dsdc_n1455));
   NOR3_X2 U_dsdc_U2046 (.ZN(U_dsdc_n1584), 
	.A3(U_dsdc_rcar_cnt1_0_), 
	.A2(U_dsdc_rcar_cnt1_1_), 
	.A1(U_dsdc_rcar_cnt1_2_));
   NOR3_X2 U_dsdc_U2045 (.ZN(U_dsdc_n1728), 
	.A3(FE_PHN969_U_dsdc_n1727), 
	.A2(U_dsdc_xsr_cnt_7_), 
	.A1(U_dsdc_xsr_cnt_8_));
   NAND2_X1 U_dsdc_U2043 (.ZN(U_dsdc_n867), 
	.A2(U_dsdc_access_cs_0_), 
	.A1(U_dsdc_n1296));
   INV_X4 U_dsdc_U2042 (.ZN(U_dsdc_n2063), 
	.A(U_dsdc_n1577));
   AND3_X4 U_dsdc_U2041 (.ZN(ctl_init_done), 
	.A3(U_dsdc_n1489), 
	.A2(U_dsdc_n1430), 
	.A1(U_dsdc_n1728));
   NAND3_X1 U_dsdc_U2039 (.ZN(U_dsdc_n653), 
	.A3(U_dsdc_n170), 
	.A2(U_dsdc_access_cs_4_), 
	.A1(U_dsdc_n1427));
   AOI22_X1 U_dsdc_U2038 (.ZN(U_dsdc_n729), 
	.B2(U_dsdc_n165), 
	.B1(U_dsdc_n1412), 
	.A2(U_dsdc_n1425), 
	.A1(U_dsdc_n1424));
   XOR2_X2 U_dsdc_U2037 (.Z(U_dsdc_num_row[3]), 
	.B(U_dsdc_n612), 
	.A(U_dsdc_N4241));
   OAI21_X1 U_dsdc_U2036 (.ZN(U_dsdc_n1370), 
	.B2(U_dsdc_access_cs_0_), 
	.B1(U_dsdc_n1356), 
	.A(U_dsdc_n1355));
   XNOR2_X2 U_dsdc_U2035 (.ZN(U_dsdc_n1657), 
	.B(U_dsdc_n1662), 
	.A(FE_PHN3054_cr_row_addr_width_2_));
   XOR2_X2 U_dsdc_U2034 (.Z(U_dsdc_num_row[15]), 
	.B(U_dsdc_n611), 
	.A(U_dsdc_N4253));
   XOR2_X2 U_dsdc_U2032 (.Z(U_dsdc_num_row[2]), 
	.B(U_dsdc_n598), 
	.A(U_dsdc_N4240));
   XNOR2_X2 U_dsdc_U2031 (.ZN(U_dsdc_num_row[7]), 
	.B(U_dsdc_n346), 
	.A(U_dsdc_n616));
   XNOR2_X2 U_dsdc_U2030 (.ZN(U_dsdc_num_row[13]), 
	.B(U_dsdc_n399), 
	.A(U_dsdc_n609));
   XNOR2_X2 U_dsdc_U2029 (.ZN(U_dsdc_num_row[5]), 
	.B(U_dsdc_n345), 
	.A(U_dsdc_n614));
   XNOR2_X2 U_dsdc_U2028 (.ZN(U_dsdc_num_row[10]), 
	.B(U_dsdc_n606), 
	.A(U_dsdc_N4248));
   XNOR2_X2 U_dsdc_U2027 (.ZN(U_dsdc_num_row[6]), 
	.B(U_dsdc_n615), 
	.A(U_dsdc_N4244));
   XNOR2_X2 U_dsdc_U2026 (.ZN(U_dsdc_num_row[8]), 
	.B(U_dsdc_n617), 
	.A(U_dsdc_N4246));
   XNOR2_X2 U_dsdc_U2025 (.ZN(U_dsdc_num_row[4]), 
	.B(U_dsdc_n613), 
	.A(U_dsdc_N4242));
   XNOR2_X2 U_dsdc_U2024 (.ZN(U_dsdc_num_row[14]), 
	.B(U_dsdc_n610), 
	.A(U_dsdc_N4252));
   XNOR2_X2 U_dsdc_U2023 (.ZN(U_dsdc_num_row[12]), 
	.B(U_dsdc_n608), 
	.A(U_dsdc_N4250));
   AOI222_X1 U_dsdc_U2022 (.ZN(U_dsdc_n1267), 
	.C2(hiu_burst_size[5]), 
	.C1(U_dsdc_n1270), 
	.B2(U_dsdc_n1269), 
	.B1(FE_PHN1890_U_dsdc_r_burst_size_5_), 
	.A2(U_dsdc_cas_cnt_5_), 
	.A1(U_dsdc_n1268));
   OR3_X4 U_dsdc_U2021 (.ZN(U_dsdc_n1881), 
	.A3(U_dsdc_n1875), 
	.A2(U_dsdc_n1876), 
	.A1(U_dsdc_n2073));
   MUX2_X2 U_dsdc_U2020 (.Z(U_dsdc_n215), 
	.S(U_dsdc_delta_delay_1_), 
	.B(U_dsdc_n1879), 
	.A(U_dsdc_n1880));
   NAND3_X1 U_dsdc_U2019 (.ZN(U_dsdc_n1347), 
	.A3(U_dsdc_n1395), 
	.A2(ad_sdram_chip_select_0_), 
	.A1(U_dsdc_n1345));
   NAND3_X2 U_dsdc_U2018 (.ZN(U_dsdc_n1815), 
	.A3(U_dsdc_n2013), 
	.A2(U_dsdc_n1546), 
	.A1(U_dsdc_n1409));
   NOR2_X2 U_dsdc_U2016 (.ZN(U_dsdc_n1750), 
	.A2(U_dsdc_n1754), 
	.A1(U_dsdc_n1728));
   OR3_X4 U_dsdc_U2015 (.ZN(U_dsdc_n2079), 
	.A3(U_dsdc_n2074), 
	.A2(U_dsdc_n1415), 
	.A1(U_dsdc_n1425));
   NOR2_X2 U_dsdc_U2014 (.ZN(U_dsdc_n687), 
	.A2(U_dsdc_r_burst_size_1_), 
	.A1(U_dsdc_r_burst_size_2_));
   NOR2_X2 U_dsdc_U2011 (.ZN(U_dsdc_n1415), 
	.A2(U_dsdc_n690), 
	.A1(U_dsdc_n660));
   NOR2_X2 U_dsdc_U2010 (.ZN(U_dsdc_n1082), 
	.A2(FE_PHN1212_U_dsdc_cas_latency_cnt_1_), 
	.A1(FE_PHN2036_U_dsdc_cas_latency_cnt_0_));
   NOR2_X2 U_dsdc_U2008 (.ZN(U_dsdc_n1163), 
	.A2(U_dsdc_rcd_cnt_2_), 
	.A1(U_dsdc_n1165));
   NAND2_X2 U_dsdc_U2007 (.ZN(U_dsdc_n904), 
	.A2(U_dsdc_r_wrapped_burst), 
	.A1(U_dsdc_n1312));
   NOR2_X2 U_dsdc_U2006 (.ZN(U_dsdc_n1296), 
	.A2(U_dsdc_wr_cnt_2_), 
	.A1(U_dsdc_n1297));
   NOR2_X2 U_dsdc_U2005 (.ZN(U_dsdc_n1436), 
	.A2(cr_do_power_down), 
	.A1(power_down));
   NOR2_X2 U_dsdc_U2004 (.ZN(U_dsdc_n1153), 
	.A2(FE_PHN1158_U_dsdc_bm_ras_cnt_max_1_), 
	.A1(FE_PHN2034_U_dsdc_bm_ras_cnt_max_0_));
   NOR2_X2 U_dsdc_U2003 (.ZN(U_dsdc_n1437), 
	.A2(FE_PHN841_U_dsdc_bm_ras_cnt_max_3_), 
	.A1(FE_PHN1200_U_dsdc_n1161));
   OAI21_X2 U_dsdc_U2002 (.ZN(U_dsdc_n1336), 
	.B2(U_dsdc_n1292), 
	.B1(U_dsdc_n1294), 
	.A(U_dsdc_n1978));
   NOR2_X2 U_dsdc_U2001 (.ZN(U_dsdc_n1394), 
	.A2(U_dsdc_n1336), 
	.A1(U_dsdc_n1325));
   NAND2_X2 U_dsdc_U2000 (.ZN(U_dsdc_n725), 
	.A2(U_dsdc_access_cs_4_), 
	.A1(U_dsdc_n964));
   NOR2_X2 U_dsdc_U1999 (.ZN(U_dsdc_n1410), 
	.A2(U_dsdc_n1309), 
	.A1(U_dsdc_n904));
   NOR2_X2 U_dsdc_U1998 (.ZN(U_dsdc_n881), 
	.A2(U_dsdc_n1312), 
	.A1(U_dsdc_n1309));
   NAND2_X2 U_dsdc_U1997 (.ZN(U_dsdc_n1040), 
	.A2(U_dsdc_n433), 
	.A1(U_dsdc_i_col_addr_1_));
   NOR2_X2 U_dsdc_U1996 (.ZN(U_dsdc_n1434), 
	.A2(U_dsdc_n341), 
	.A1(U_dsdc_n641));
   NOR2_X2 U_dsdc_U1995 (.ZN(U_dsdc_n1269), 
	.A2(U_dsdc_n1300), 
	.A1(U_dsdc_n1258));
   NOR3_X2 U_dsdc_U1994 (.ZN(U_dsdc_n1340), 
	.A3(U_dsdc_n1268), 
	.A2(U_dsdc_n1269), 
	.A1(U_dsdc_n1270));
   NAND3_X2 U_dsdc_U1993 (.ZN(U_dsdc_n1975), 
	.A3(n84), 
	.A2(U_dsdc_n1428), 
	.A1(sdram_req_i));
   INV_X4 U_dsdc_U1992 (.ZN(U_dsdc_n670), 
	.A(U_dsdc_n1975));
   NAND2_X2 U_dsdc_U1991 (.ZN(U_dsdc_n903), 
	.A2(U_dsdc_n328), 
	.A1(U_dsdc_n1312));
   NOR2_X2 U_dsdc_U1990 (.ZN(U_dsdc_n663), 
	.A2(U_dsdc_n1446), 
	.A1(FE_PHN1227_U_dsdc_cas_cnt_2_));
   NAND2_X2 U_dsdc_U1989 (.ZN(U_dsdc_n991), 
	.A2(U_dsdc_n305), 
	.A1(U_dsdc_n1061));
   NAND2_X2 U_dsdc_U1988 (.ZN(U_dsdc_n1094), 
	.A2(U_dsdc_n331), 
	.A1(U_dsdc_n1082));
   NOR2_X2 U_dsdc_U1987 (.ZN(U_dsdc_n1414), 
	.A2(FE_PHN1153_U_dsdc_cas_latency_cnt_3_), 
	.A1(FE_PHN1585_U_dsdc_n1094));
   NAND2_X2 U_dsdc_U1986 (.ZN(U_dsdc_n746), 
	.A2(U_dsdc_n735), 
	.A1(U_dsdc_n1344));
   INV_X4 U_dsdc_U1985 (.ZN(U_dsdc_n2071), 
	.A(U_dsdc_n1415));
   NOR2_X2 U_dsdc_U1984 (.ZN(U_dsdc_n936), 
	.A2(U_dsdc_n703), 
	.A1(U_dsdc_n2071));
   NAND2_X2 U_dsdc_U1983 (.ZN(U_dsdc_n741), 
	.A2(U_dsdc_access_cs_2_), 
	.A1(U_dsdc_n654));
   NOR2_X2 U_dsdc_U1982 (.ZN(U_dsdc_n1419), 
	.A2(U_dsdc_data_flag), 
	.A1(U_dsdc_early_term_flag));
   NAND2_X2 U_dsdc_U1981 (.ZN(U_dsdc_n756), 
	.A2(U_dsdc_n737), 
	.A1(U_dsdc_n738));
   NAND2_X2 U_dsdc_U1980 (.ZN(U_dsdc_n745), 
	.A2(U_dsdc_n1079), 
	.A1(U_dsdc_n756));
   INV_X4 U_dsdc_U1979 (.ZN(U_dsdc_n934), 
	.A(U_dsdc_n1412));
   NAND3_X2 U_dsdc_U1976 (.ZN(U_dsdc_RSOP_1683_C2_CONTROL1), 
	.A3(U_dsdc_n744), 
	.A2(U_dsdc_n745), 
	.A1(U_dsdc_n746));
   NOR2_X2 U_dsdc_U1975 (.ZN(U_dsdc_n1418), 
	.A2(U_dsdc_n711), 
	.A1(U_dsdc_n660));
   NAND2_X2 U_dsdc_U1974 (.ZN(U_dsdc_n1165), 
	.A2(U_dsdc_n174), 
	.A1(U_dsdc_n326));
   NAND2_X2 U_dsdc_U1973 (.ZN(U_dsdc_n1637), 
	.A2(U_dsdc_n1484), 
	.A1(cr_s_ready_valid));
   INV_X4 U_dsdc_U1972 (.ZN(U_dsdc_n1444), 
	.A(FE_PHN671_U_dsdc_n1637));
   NAND2_X2 U_dsdc_U1971 (.ZN(U_dsdc_n1876), 
	.A2(U_dsdc_n1414), 
	.A1(U_dsdc_n1444));
   NAND2_X2 U_dsdc_U1970 (.ZN(U_dsdc_n760), 
	.A2(U_dsdc_n305), 
	.A1(U_dsdc_n668));
   NOR2_X2 U_dsdc_U1969 (.ZN(U_dsdc_DP_OP_1642_126_2028_I4), 
	.A2(U_dsdc_n760), 
	.A1(U_dsdc_n1876));
   NAND4_X2 U_dsdc_U1968 (.ZN(U_dsdc_n1380), 
	.A4(U_dsdc_n755), 
	.A3(U_dsdc_n1258), 
	.A2(U_dsdc_n601), 
	.A1(U_dsdc_n1546));
   NAND2_X2 U_dsdc_U1967 (.ZN(U_dsdc_n753), 
	.A2(U_dsdc_n1258), 
	.A1(U_dsdc_n1546));
   NAND2_X2 U_dsdc_U1966 (.ZN(U_dsdc_DP_OP_1642_126_2028_I6), 
	.A2(U_dsdc_n601), 
	.A1(U_dsdc_n754));
   AOI22_X2 U_dsdc_U1965 (.ZN(U_dsdc_n750), 
	.B2(U_dsdc_r_burst_size_2_), 
	.B1(U_dsdc_n751), 
	.A2(U_dsdc_data_cnt_2_), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n85));
   INV_X4 U_dsdc_U1964 (.ZN(U_dsdc_DP_OP_1642_126_2028_I5_1_), 
	.A(U_dsdc_n752));
   OAI211_X2 U_dsdc_U1963 (.ZN(U_dsdc_DP_OP_1642_126_2028_n86), 
	.C2(U_dsdc_n342), 
	.C1(U_dsdc_n754), 
	.B(U_dsdc_n755), 
	.A(U_dsdc_n601));
   NOR2_X2 U_dsdc_U1962 (.ZN(U_dsdc_n1825), 
	.A2(U_dsdc_data_cnt_0_), 
	.A1(U_dsdc_n1444));
   NAND2_X2 U_dsdc_U1961 (.ZN(U_dsdc_n1823), 
	.A2(U_dsdc_n436), 
	.A1(U_dsdc_n1825));
   NOR2_X2 U_dsdc_U1960 (.ZN(U_dsdc_n1822), 
	.A2(FE_PHN773_U_dsdc_n1823), 
	.A1(U_dsdc_data_cnt_2_));
   NAND2_X2 U_dsdc_U1959 (.ZN(U_dsdc_n1820), 
	.A2(U_dsdc_n437), 
	.A1(U_dsdc_n1822));
   NOR2_X2 U_dsdc_U1958 (.ZN(U_dsdc_n762), 
	.A2(U_dsdc_data_cnt_4_), 
	.A1(U_dsdc_n1820));
   AOI21_X2 U_dsdc_U1957 (.ZN(U_dsdc_n757), 
	.B2(U_cr_n58), 
	.B1(U_dsdc_n1344), 
	.A(U_dsdc_n756));
   NOR2_X2 U_dsdc_U1956 (.ZN(U_dsdc_n764), 
	.A2(U_dsdc_n1079), 
	.A1(U_dsdc_n757));
   NAND2_X2 U_dsdc_U1955 (.ZN(U_dsdc_n758), 
	.A2(U_dsdc_n1412), 
	.A1(U_dsdc_n668));
   OAI22_X2 U_dsdc_U1954 (.ZN(U_dsdc_n1381), 
	.B2(U_dsdc_n758), 
	.B1(U_dsdc_n759), 
	.A2(U_dsdc_n760), 
	.A1(U_dsdc_n761));
   INV_X4 U_dsdc_U1953 (.ZN(U_dsdc_n814), 
	.A(debug_ad_row_addr[1]));
   NAND2_X2 U_dsdc_U1951 (.ZN(U_dsdc_n799), 
	.A2(U_dsdc_bm_row_addr_2__1_), 
	.A1(U_dsdc_n159));
   INV_X4 U_dsdc_U1950 (.ZN(U_dsdc_n815), 
	.A(U_dsdc_n813));
   NAND2_X2 U_dsdc_U1948 (.ZN(U_dsdc_n791), 
	.A2(U_dsdc_bm_row_addr_3__11_), 
	.A1(U_dsdc_n978));
   NAND2_X2 U_dsdc_U1947 (.ZN(U_dsdc_n790), 
	.A2(U_dsdc_bm_row_addr_2__11_), 
	.A1(U_dsdc_n159));
   INV_X4 U_dsdc_U1946 (.ZN(U_dsdc_n812), 
	.A(U_dsdc_n810));
   INV_X4 U_dsdc_U1943 (.ZN(U_dsdc_n803), 
	.A(debug_ad_row_addr[9]));
   NAND2_X2 U_dsdc_U1942 (.ZN(U_dsdc_n787), 
	.A2(U_dsdc_bm_row_addr_2__9_), 
	.A1(U_dsdc_n159));
   INV_X4 U_dsdc_U1941 (.ZN(U_dsdc_n804), 
	.A(U_dsdc_n802));
   NOR3_X2 U_dsdc_U1940 (.ZN(U_dsdc_n524), 
	.A3(U_dsdc_n804), 
	.A2(U_dsdc_n803), 
	.A1(U_dsdc_bm_row_addr_0__9_));
   NAND2_X2 U_dsdc_U1939 (.ZN(U_dsdc_n794), 
	.A2(U_dsdc_bm_row_addr_3__5_), 
	.A1(U_dsdc_n978));
   NAND2_X2 U_dsdc_U1938 (.ZN(U_dsdc_n793), 
	.A2(U_dsdc_bm_row_addr_2__5_), 
	.A1(U_dsdc_n159));
   NAND2_X2 U_dsdc_U1937 (.ZN(U_dsdc_n522), 
	.A2(U_dsdc_n808), 
	.A1(debug_ad_row_addr[5]));
   NOR2_X2 U_dsdc_U1936 (.ZN(U_dsdc_n523), 
	.A2(U_dsdc_n522), 
	.A1(U_dsdc_bm_row_addr_0__5_));
   NOR2_X2 U_dsdc_U1935 (.ZN(U_dsdc_n535), 
	.A2(U_dsdc_n523), 
	.A1(U_dsdc_n524));
   NAND2_X2 U_dsdc_U1934 (.ZN(U_dsdc_n784), 
	.A2(U_dsdc_bm_row_addr_3__15_), 
	.A1(U_dsdc_n978));
   NAND2_X2 U_dsdc_U1933 (.ZN(U_dsdc_n783), 
	.A2(U_dsdc_bm_row_addr_2__15_), 
	.A1(U_dsdc_n159));
   INV_X4 U_dsdc_U1932 (.ZN(U_dsdc_n807), 
	.A(U_dsdc_n805));
   NAND2_X2 U_dsdc_U1931 (.ZN(U_dsdc_n527), 
	.A2(U_dsdc_n806), 
	.A1(U_dsdc_n807));
   NAND2_X2 U_dsdc_U1930 (.ZN(U_dsdc_n526), 
	.A2(U_dsdc_n814), 
	.A1(U_dsdc_n815));
   NAND2_X2 U_dsdc_U1929 (.ZN(U_dsdc_n525), 
	.A2(U_dsdc_n812), 
	.A1(U_addrdec_n231));
   NAND3_X2 U_dsdc_U1928 (.ZN(U_dsdc_n528), 
	.A3(U_dsdc_n525), 
	.A2(U_dsdc_n526), 
	.A1(U_dsdc_n527));
   INV_X4 U_dsdc_U1927 (.ZN(U_dsdc_n531), 
	.A(U_dsdc_n528));
   NAND2_X2 U_dsdc_U1926 (.ZN(U_dsdc_n530), 
	.A2(U_dsdc_n804), 
	.A1(U_dsdc_n803));
   INV_X4 U_dsdc_U1925 (.ZN(U_dsdc_n1104), 
	.A(debug_ad_row_addr[5]));
   NAND2_X2 U_dsdc_U1924 (.ZN(U_dsdc_n529), 
	.A2(U_dsdc_n809), 
	.A1(U_dsdc_n1104));
   NAND3_X2 U_dsdc_U1923 (.ZN(U_dsdc_n532), 
	.A3(U_dsdc_n529), 
	.A2(U_dsdc_n530), 
	.A1(U_dsdc_n531));
   NOR2_X2 U_dsdc_U1922 (.ZN(U_dsdc_n533), 
	.A2(U_dsdc_n807), 
	.A1(U_dsdc_n806));
   NOR2_X2 U_dsdc_U1921 (.ZN(U_dsdc_n534), 
	.A2(U_dsdc_n177), 
	.A1(U_dsdc_n532));
   NAND3_X2 U_dsdc_U1920 (.ZN(U_dsdc_n537), 
	.A3(U_dsdc_n534), 
	.A2(U_dsdc_n535), 
	.A1(U_dsdc_n536));
   NAND3_X2 U_dsdc_U1919 (.ZN(U_dsdc_n785), 
	.A3(U_dsdc_n776), 
	.A2(U_dsdc_n777), 
	.A1(U_dsdc_n778));
   NAND3_X2 U_dsdc_U1917 (.ZN(U_dsdc_n602), 
	.A3(U_dsdc_n795), 
	.A2(U_dsdc_n796), 
	.A1(U_dsdc_n797));
   INV_X4 U_dsdc_U1916 (.ZN(U_dsdc_n816), 
	.A(debug_ad_row_addr[7]));
   NAND2_X2 U_dsdc_U1915 (.ZN(U_dsdc_n540), 
	.A2(U_dsdc_n816), 
	.A1(U_dsdc_n602));
   NAND2_X2 U_dsdc_U1914 (.ZN(U_dsdc_n517), 
	.A2(U_dsdc_n515), 
	.A1(U_dsdc_n516));
   AOI21_X2 U_dsdc_U1913 (.ZN(U_dsdc_n519), 
	.B2(U_dsdc_bm_row_addr_2__12_), 
	.B1(U_dsdc_n159), 
	.A(U_dsdc_n517));
   NAND3_X2 U_dsdc_U1912 (.ZN(U_dsdc_n541), 
	.A3(U_dsdc_n539), 
	.A2(U_dsdc_n540), 
	.A1(U_dsdc_n538));
   INV_X4 U_dsdc_U1911 (.ZN(U_dsdc_n487), 
	.A(U_dsdc_n541));
   INV_X4 U_dsdc_U1909 (.ZN(U_dsdc_n801), 
	.A(debug_ad_row_addr[3]));
   NAND2_X2 U_dsdc_U1908 (.ZN(U_dsdc_n502), 
	.A2(U_dsdc_bm_row_addr_3__6_), 
	.A1(U_dsdc_n978));
   NAND3_X2 U_dsdc_U1907 (.ZN(U_dsdc_n503), 
	.A3(U_dsdc_n500), 
	.A2(U_dsdc_n501), 
	.A1(U_dsdc_n502));
   AOI21_X2 U_dsdc_U1906 (.ZN(U_dsdc_n504), 
	.B2(U_dsdc_bm_row_addr_2__6_), 
	.B1(U_dsdc_n159), 
	.A(U_dsdc_n503));
   NAND2_X2 U_dsdc_U1905 (.ZN(U_dsdc_n508), 
	.A2(U_dsdc_bm_row_addr_3__8_), 
	.A1(U_dsdc_n978));
   INV_X4 U_dsdc_U1904 (.ZN(U_dsdc_n600), 
	.A(U_dsdc_n604));
   NOR2_X2 U_dsdc_U1901 (.ZN(U_dsdc_n507), 
	.A2(U_dsdc_n314), 
	.A1(n86));
   NAND2_X2 U_dsdc_U1900 (.ZN(U_dsdc_n509), 
	.A2(U_dsdc_n507), 
	.A1(U_dsdc_n508));
   AOI21_X2 U_dsdc_U1899 (.ZN(U_dsdc_n510), 
	.B2(U_dsdc_bm_row_addr_2__8_), 
	.B1(U_dsdc_n159), 
	.A(U_dsdc_n509));
   NOR2_X2 U_dsdc_U1898 (.ZN(U_dsdc_n513), 
	.A2(U_dsdc_n511), 
	.A1(U_dsdc_n512));
   NAND3_X2 U_dsdc_U1897 (.ZN(U_dsdc_n542), 
	.A3(U_dsdc_n513), 
	.A2(U_dsdc_n514), 
	.A1(U_dsdc_n332));
   NAND2_X2 U_dsdc_U1896 (.ZN(U_dsdc_n555), 
	.A2(U_dsdc_bm_row_addr_3__4_), 
	.A1(U_dsdc_n978));
   NOR2_X2 U_dsdc_U1895 (.ZN(U_dsdc_n552), 
	.A2(U_dsdc_n600), 
	.A1(U_dsdc_n339));
   AOI21_X2 U_dsdc_U1894 (.ZN(U_dsdc_n553), 
	.B2(U_dsdc_bm_row_addr_0__4_), 
	.B1(U_dsdc_n998), 
	.A(U_dsdc_n552));
   NAND2_X2 U_dsdc_U1893 (.ZN(U_dsdc_n556), 
	.A2(U_dsdc_n553), 
	.A1(U_dsdc_n555));
   AOI21_X2 U_dsdc_U1892 (.ZN(U_dsdc_n557), 
	.B2(U_dsdc_bm_row_addr_2__4_), 
	.B1(U_dsdc_n159), 
	.A(U_dsdc_n556));
   NAND2_X2 U_dsdc_U1891 (.ZN(U_dsdc_n559), 
	.A2(U_dsdc_bm_row_addr_3__0_), 
	.A1(U_dsdc_n978));
   NAND2_X2 U_dsdc_U1889 (.ZN(U_dsdc_n560), 
	.A2(U_dsdc_n558), 
	.A1(U_dsdc_n559));
   NAND2_X2 U_dsdc_U1887 (.ZN(U_dsdc_n563), 
	.A2(U_dsdc_bm_row_addr_3__2_), 
	.A1(U_dsdc_n978));
   NAND2_X2 U_dsdc_U1886 (.ZN(U_dsdc_n564), 
	.A2(U_dsdc_n562), 
	.A1(U_dsdc_n563));
   NOR2_X2 U_dsdc_U1885 (.ZN(U_dsdc_n565), 
	.A2(U_dsdc_n330), 
	.A1(U_dsdc_n564));
   NOR3_X2 U_dsdc_U1884 (.ZN(U_dsdc_n569), 
	.A3(U_dsdc_n566), 
	.A2(U_dsdc_n567), 
	.A1(U_dsdc_n568));
   NOR3_X2 U_dsdc_U1883 (.ZN(U_dsdc_n551), 
	.A3(U_dsdc_bm_row_addr_0__3_), 
	.A2(U_dsdc_n801), 
	.A1(U_dsdc_n798));
   NAND2_X2 U_dsdc_U1882 (.ZN(U_dsdc_n544), 
	.A2(U_dsdc_bm_row_addr_3__10_), 
	.A1(U_dsdc_n978));
   NOR2_X2 U_dsdc_U1881 (.ZN(U_dsdc_n543), 
	.A2(U_dsdc_n312), 
	.A1(U_dsdc_n176));
   NAND2_X2 U_dsdc_U1880 (.ZN(U_dsdc_n545), 
	.A2(U_dsdc_n543), 
	.A1(U_dsdc_n544));
   AOI21_X2 U_dsdc_U1879 (.ZN(U_dsdc_n546), 
	.B2(U_dsdc_bm_row_addr_2__10_), 
	.B1(U_dsdc_n159), 
	.A(U_dsdc_n545));
   NAND2_X2 U_dsdc_U1878 (.ZN(U_dsdc_n547), 
	.A2(U_dsdc_bm_row_addr_3__14_), 
	.A1(U_dsdc_n978));
   NOR3_X2 U_dsdc_U1877 (.ZN(U_dsdc_n570), 
	.A3(U_dsdc_n549), 
	.A2(U_dsdc_n550), 
	.A1(U_dsdc_n551));
   NAND2_X2 U_dsdc_U1876 (.ZN(U_dsdc_n486), 
	.A2(U_dsdc_n570), 
	.A1(U_dsdc_n569));
   NOR2_X2 U_dsdc_U1875 (.ZN(U_dsdc_n485), 
	.A2(U_dsdc_n486), 
	.A1(U_dsdc_n542));
   NAND2_X2 U_dsdc_U1874 (.ZN(U_dsdc_n488), 
	.A2(debug_ad_row_addr[5]), 
	.A1(U_dsdc_n808));
   NOR2_X2 U_dsdc_U1872 (.ZN(U_dsdc_n491), 
	.A2(U_dsdc_n801), 
	.A1(U_dsdc_n798));
   NOR3_X2 U_dsdc_U1871 (.ZN(U_dsdc_n498), 
	.A3(U_dsdc_n491), 
	.A2(U_dsdc_n318), 
	.A1(U_dsdc_n492));
   NAND2_X2 U_dsdc_U1870 (.ZN(U_dsdc_n493), 
	.A2(U_dsdc_n1104), 
	.A1(U_dsdc_bm_row_addr_0__5_));
   NOR3_X2 U_dsdc_U1869 (.ZN(U_dsdc_n497), 
	.A3(U_dsdc_n494), 
	.A2(U_dsdc_n495), 
	.A1(U_dsdc_n496));
   AOI21_X2 U_dsdc_U1868 (.ZN(U_dsdc_n571), 
	.B2(U_dsdc_n498), 
	.B1(U_dsdc_n499), 
	.A(U_dsdc_n497));
   INV_X4 U_dsdc_U1867 (.ZN(U_dsdc_n484), 
	.A(U_dsdc_n571));
   NAND3_X2 U_dsdc_U1866 (.ZN(U_dsdc_n483), 
	.A3(U_dsdc_n484), 
	.A2(U_dsdc_n485), 
	.A1(U_dsdc_n487));
   NOR2_X2 U_dsdc_U1865 (.ZN(U_dsdc_n818), 
	.A2(U_dsdc_n827), 
	.A1(U_dsdc_n884));
   NAND2_X2 U_dsdc_U1864 (.ZN(U_dsdc_n1196), 
	.A2(U_dsdc_n420), 
	.A1(U_dsdc_n186));
   NOR2_X2 U_dsdc_U1863 (.ZN(U_dsdc_n1200), 
	.A2(FE_PHN1889_U_dsdc_bm_ras_cnt_1__2_), 
	.A1(FE_PHN1154_U_dsdc_n1196));
   NAND2_X2 U_dsdc_U1862 (.ZN(U_dsdc_n1195), 
	.A2(FE_PHN1336_U_dsdc_n364), 
	.A1(U_dsdc_n1200));
   NAND2_X2 U_dsdc_U1861 (.ZN(U_dsdc_n1297), 
	.A2(U_dsdc_n397), 
	.A1(U_dsdc_n195));
   INV_X4 U_dsdc_U1860 (.ZN(U_dsdc_n1294), 
	.A(U_dsdc_n1296));
   NAND2_X2 U_dsdc_U1859 (.ZN(U_dsdc_n1238), 
	.A2(U_dsdc_n421), 
	.A1(U_dsdc_n187));
   NOR2_X2 U_dsdc_U1858 (.ZN(U_dsdc_n1244), 
	.A2(FE_PHN1891_U_dsdc_bm_ras_cnt_3__2_), 
	.A1(FE_PHN1497_U_dsdc_n1238));
   NAND2_X2 U_dsdc_U1857 (.ZN(U_dsdc_n1237), 
	.A2(FE_PHN1333_U_dsdc_n382), 
	.A1(U_dsdc_n1244));
   NAND2_X2 U_dsdc_U1856 (.ZN(U_dsdc_n1210), 
	.A2(U_dsdc_n422), 
	.A1(U_dsdc_n188));
   NOR2_X2 U_dsdc_U1855 (.ZN(U_dsdc_n1214), 
	.A2(U_dsdc_bm_ras_cnt_2__2_), 
	.A1(FE_PHN1155_U_dsdc_n1210));
   NAND2_X2 U_dsdc_U1854 (.ZN(U_dsdc_n1209), 
	.A2(FE_PHN1334_U_dsdc_n365), 
	.A1(U_dsdc_n1214));
   NAND2_X2 U_dsdc_U1853 (.ZN(U_dsdc_n1182), 
	.A2(U_dsdc_n424), 
	.A1(U_dsdc_n189));
   NOR2_X2 U_dsdc_U1852 (.ZN(U_dsdc_n1186), 
	.A2(U_dsdc_bm_ras_cnt_0__2_), 
	.A1(FE_PHN1156_U_dsdc_n1182));
   NAND2_X2 U_dsdc_U1851 (.ZN(U_dsdc_n1181), 
	.A2(FE_PHN1337_U_dsdc_n363), 
	.A1(U_dsdc_n1186));
   NOR2_X2 U_dsdc_U1850 (.ZN(U_dsdc_n980), 
	.A2(U_dsdc_n1546), 
	.A1(U_dsdc_n979));
   INV_X4 U_dsdc_U1849 (.ZN(U_dsdc_n999), 
	.A(U_dsdc_oldest_bank_0_));
   NOR2_X2 U_dsdc_U1848 (.ZN(U_dsdc_n840), 
	.A2(U_dsdc_n837), 
	.A1(U_dsdc_n999));
   NOR2_X2 U_dsdc_U1847 (.ZN(U_dsdc_n839), 
	.A2(U_dsdc_n838), 
	.A1(U_dsdc_oldest_bank_0_));
   OAI21_X2 U_dsdc_U1846 (.ZN(U_dsdc_n846), 
	.B2(U_dsdc_n839), 
	.B1(U_dsdc_n840), 
	.A(U_dsdc_n1000));
   NOR2_X2 U_dsdc_U1845 (.ZN(U_dsdc_n844), 
	.A2(U_dsdc_n841), 
	.A1(U_dsdc_n999));
   NOR2_X2 U_dsdc_U1844 (.ZN(U_dsdc_n843), 
	.A2(U_dsdc_n842), 
	.A1(U_dsdc_oldest_bank_0_));
   OAI21_X2 U_dsdc_U1843 (.ZN(U_dsdc_n845), 
	.B2(U_dsdc_n843), 
	.B1(U_dsdc_n844), 
	.A(U_dsdc_oldest_bank_1_));
   NAND3_X2 U_dsdc_U1842 (.ZN(U_dsdc_n986), 
	.A3(U_dsdc_n1296), 
	.A2(U_dsdc_n845), 
	.A1(U_dsdc_n846));
   INV_X4 U_dsdc_U1841 (.ZN(U_dsdc_n940), 
	.A(U_dsdc_n1483));
   NOR2_X2 U_dsdc_U1840 (.ZN(U_dsdc_n819), 
	.A2(U_dsdc_n940), 
	.A1(U_dsdc_n827));
   NAND2_X2 U_dsdc_U1839 (.ZN(U_dsdc_n825), 
	.A2(U_dsdc_n819), 
	.A1(U_dsdc_n884));
   INV_X4 U_dsdc_U1838 (.ZN(U_dsdc_n984), 
	.A(U_dsdc_n825));
   NOR2_X2 U_dsdc_U1837 (.ZN(U_dsdc_n1003), 
	.A2(U_dsdc_n985), 
	.A1(U_dsdc_n986));
   INV_X4 U_dsdc_U1836 (.ZN(U_dsdc_n1004), 
	.A(U_dsdc_n1003));
   NAND3_X2 U_dsdc_U1835 (.ZN(U_dsdc_n1017), 
	.A3(FE_PHN1093_U_dsdc_n340), 
	.A2(U_dsdc_n180), 
	.A1(U_dsdc_n1326));
   NOR3_X2 U_dsdc_U1834 (.ZN(U_dsdc_n1022), 
	.A3(U_dsdc_bm_num_open_bank_2_), 
	.A2(U_dsdc_bm_num_open_bank_3_), 
	.A1(U_dsdc_n1017));
   NAND2_X2 U_dsdc_U1833 (.ZN(U_dsdc_n975), 
	.A2(U_dsdc_n826), 
	.A1(U_dsdc_n984));
   NAND2_X2 U_dsdc_U1832 (.ZN(U_dsdc_n1345), 
	.A2(U_dsdc_n1483), 
	.A1(U_dsdc_n975));
   OAI21_X2 U_dsdc_U1831 (.ZN(U_dsdc_n829), 
	.B2(U_dsdc_bm_rc_cnt_0__3_), 
	.B1(U_dsdc_bm_rc_cnt_0__2_), 
	.A(U_dsdc_n998));
   NAND2_X2 U_dsdc_U1830 (.ZN(U_dsdc_n1228), 
	.A2(U_dsdc_n190), 
	.A1(U_dsdc_n400));
   NAND2_X2 U_dsdc_U1829 (.ZN(U_dsdc_n1203), 
	.A2(U_dsdc_n191), 
	.A1(U_dsdc_n401));
   AOI22_X2 U_dsdc_U1828 (.ZN(U_dsdc_n834), 
	.B2(U_dsdc_n1203), 
	.B1(U_dsdc_n159), 
	.A2(U_dsdc_n1228), 
	.A1(U_dsdc_n978));
   NAND2_X2 U_dsdc_U1827 (.ZN(U_dsdc_n1175), 
	.A2(U_dsdc_n192), 
	.A1(U_dsdc_n402));
   NAND2_X2 U_dsdc_U1826 (.ZN(U_dsdc_n1189), 
	.A2(U_dsdc_n193), 
	.A1(U_dsdc_n419));
   AOI22_X2 U_dsdc_U1825 (.ZN(U_dsdc_n833), 
	.B2(U_dsdc_n1189), 
	.B1(U_dsdc_n604), 
	.A2(FE_PHN945_U_dsdc_n1175), 
	.A1(U_dsdc_n998));
   NAND3_X2 U_dsdc_U1824 (.ZN(U_dsdc_n976), 
	.A3(U_dsdc_n833), 
	.A2(U_dsdc_n834), 
	.A1(U_dsdc_n835));
   INV_X4 U_dsdc_U1823 (.ZN(U_dsdc_n988), 
	.A(U_dsdc_n827));
   NAND2_X2 U_dsdc_U1822 (.ZN(U_dsdc_n1362), 
	.A2(U_dsdc_n430), 
	.A1(U_dsdc_n1616));
   INV_X4 U_dsdc_U1821 (.ZN(U_dsdc_n1422), 
	.A(U_dsdc_n1362));
   NOR2_X2 U_dsdc_U1820 (.ZN(U_dsdc_n1384), 
	.A2(U_dsdc_n712), 
	.A1(U_dsdc_n658));
   NAND3_X2 U_dsdc_U1819 (.ZN(U_dsdc_n1020), 
	.A3(U_dsdc_bm_num_open_bank_0_), 
	.A2(U_dsdc_bm_num_open_bank_1_), 
	.A1(U_dsdc_n1166));
   NOR2_X2 U_dsdc_U1818 (.ZN(U_dsdc_n1026), 
	.A2(U_dsdc_n1021), 
	.A1(U_dsdc_n1022));
   INV_X4 U_dsdc_U1817 (.ZN(U_dsdc_n1290), 
	.A(U_dsdc_n1326));
   NAND2_X2 U_dsdc_U1816 (.ZN(U_dsdc_n2056), 
	.A2(U_dsdc_n1465), 
	.A1(U_dsdc_n1449));
   OAI21_X2 U_dsdc_U1815 (.ZN(U_dsdc_n990), 
	.B2(U_dsdc_n988), 
	.B1(U_dsdc_n1546), 
	.A(U_dsdc_n1354));
   NAND2_X2 U_dsdc_U1814 (.ZN(U_dsdc_n1161), 
	.A2(U_dsdc_n428), 
	.A1(U_dsdc_n1153));
   NAND2_X2 U_dsdc_U1813 (.ZN(U_dsdc_n1496), 
	.A2(U_dsdc_n1296), 
	.A1(U_dsdc_n1437));
   NOR2_X2 U_dsdc_U1812 (.ZN(U_dsdc_n989), 
	.A2(U_dsdc_n940), 
	.A1(U_dsdc_n1496));
   NAND2_X2 U_dsdc_U1811 (.ZN(U_dsdc_n1283), 
	.A2(U_dsdc_n989), 
	.A1(U_dsdc_n990));
   NAND2_X2 U_dsdc_U1810 (.ZN(U_dsdc_n1342), 
	.A2(U_dsdc_n1437), 
	.A1(U_dsdc_n1416));
   AOI21_X2 U_dsdc_U1809 (.ZN(U_dsdc_n995), 
	.B2(U_dsdc_n994), 
	.B1(U_dsdc_n1386), 
	.A(U_dsdc_n993));
   NAND2_X2 U_dsdc_U1808 (.ZN(U_dsdc_n1325), 
	.A2(U_dsdc_n995), 
	.A1(U_dsdc_n1283));
   NAND2_X2 U_dsdc_U1807 (.ZN(U_dsdc_n1064), 
	.A2(U_dsdc_n1412), 
	.A1(U_dsdc_n1300));
   NOR2_X2 U_dsdc_U1806 (.ZN(U_dsdc_n715), 
	.A2(U_dsdc_n165), 
	.A1(U_dsdc_n1064));
   NAND2_X2 U_dsdc_U1805 (.ZN(U_dsdc_n1978), 
	.A2(U_dsdc_n715), 
	.A1(U_dsdc_n1980));
   NAND3_X2 U_dsdc_U1804 (.ZN(U_dsdc_n1006), 
	.A3(FE_PHN683_U_dsdc_n1394), 
	.A2(U_dsdc_n1159), 
	.A1(U_dsdc_n1290));
   NAND2_X2 U_dsdc_U1803 (.ZN(U_dsdc_n1011), 
	.A2(U_dsdc_n1006), 
	.A1(U_dsdc_n1007));
   NOR2_X2 U_dsdc_U1802 (.ZN(U_dsdc_n1016), 
	.A2(U_dsdc_n1010), 
	.A1(U_dsdc_n1011));
   NAND2_X2 U_dsdc_U1801 (.ZN(U_dsdc_n1024), 
	.A2(U_dsdc_n1015), 
	.A1(U_dsdc_n1016));
   NAND2_X2 U_dsdc_U1800 (.ZN(U_dsdc_n297), 
	.A2(U_dsdc_n1025), 
	.A1(U_dsdc_n603));
   INV_X4 U_dsdc_U1799 (.ZN(U_dsdc_n900), 
	.A(U_dsdc_n914));
   INV_X4 U_dsdc_U1798 (.ZN(U_dsdc_n821), 
	.A(hiu_wrapped_burst));
   NOR2_X2 U_dsdc_U1797 (.ZN(U_dsdc_n1254), 
	.A2(U_dsdc_n1448), 
	.A1(hiu_burst_size[4]));
   NAND2_X2 U_dsdc_U1796 (.ZN(U_dsdc_n1557), 
	.A2(hiu_burst_size[0]), 
	.A1(U_dsdc_n1254));
   NOR2_X2 U_dsdc_U1795 (.ZN(U_dsdc_n1053), 
	.A2(U_dsdc_n1557), 
	.A1(U_dsdc_n821));
   NAND2_X2 U_dsdc_U1794 (.ZN(U_dsdc_n1248), 
	.A2(U_dsdc_n398), 
	.A1(U_dsdc_n194));
   NOR2_X2 U_dsdc_U1793 (.ZN(U_dsdc_n1284), 
	.A2(U_dsdc_wtr_cnt_2_), 
	.A1(U_dsdc_n1248));
   NAND2_X2 U_dsdc_U1792 (.ZN(U_dsdc_n1090), 
	.A2(U_dsdc_n1079), 
	.A1(U_dsdc_n1393));
   NOR2_X2 U_dsdc_U1791 (.ZN(U_dsdc_n1464), 
	.A2(FE_PHN787_n90), 
	.A1(s_cas_latency[1]));
   OAI221_X2 U_dsdc_U1790 (.ZN(U_dsdc_n1462), 
	.C2(FE_PHN894_U_dsdc_n1464), 
	.C1(s_cas_latency[2]), 
	.B2(U_dsdc_n1461), 
	.B1(n91), 
	.A(U_dsdc_n1460));
   NOR2_X2 U_dsdc_U1789 (.ZN(U_dsdc_n1084), 
	.A2(U_cr_n40), 
	.A1(U_dsdc_n1088));
   NOR2_X2 U_dsdc_U1788 (.ZN(U_dsdc_n1092), 
	.A2(U_dsdc_n1081), 
	.A1(FE_PHN894_U_dsdc_n1464));
   NAND4_X2 U_dsdc_U1787 (.ZN(U_dsdc_n2082), 
	.A4(U_dsdc_n164), 
	.A3(U_dsdc_n185), 
	.A2(U_dsdc_n356), 
	.A1(U_dsdc_n168));
   NOR2_X2 U_dsdc_U1786 (.ZN(U_dsdc_n1826), 
	.A2(U_dsdc_n2082), 
	.A1(U_dsdc_r_bm_close_all));
   NAND2_X2 U_dsdc_U1785 (.ZN(U_dsdc_n1942), 
	.A2(U_dsdc_n1846), 
	.A1(U_dsdc_n1826));
   NOR3_X2 U_dsdc_U1784 (.ZN(U_dsdc_n1867), 
	.A3(U_dsdc_n1942), 
	.A2(U_dsdc_n395), 
	.A1(U_dsdc_r_bm_close_bank_2_));
   INV_X4 U_dsdc_U1783 (.ZN(U_dsdc_n1941), 
	.A(U_dsdc_n2082));
   NOR2_X2 U_dsdc_U1782 (.ZN(U_dsdc_n1850), 
	.A2(U_dsdc_n1941), 
	.A1(U_dsdc_n395));
   NAND2_X2 U_dsdc_U1781 (.ZN(U_dsdc_n1860), 
	.A2(U_dsdc_n1850), 
	.A1(U_dsdc_n164));
   INV_X4 U_dsdc_U1780 (.ZN(U_dsdc_n1859), 
	.A(U_dsdc_n1867));
   NOR2_X2 U_dsdc_U1779 (.ZN(U_dsdc_n1842), 
	.A2(U_dsdc_r_close_bank_addr_1_), 
	.A1(U_dsdc_r_close_bank_addr_0_));
   NAND2_X2 U_dsdc_U1778 (.ZN(U_dsdc_n1841), 
	.A2(U_dsdc_r_close_bank_addr_1_), 
	.A1(U_dsdc_r_close_bank_addr_0_));
   NOR2_X2 U_dsdc_U1777 (.ZN(U_dsdc_n1839), 
	.A2(U_dsdc_n292), 
	.A1(U_dsdc_r_close_bank_addr_1_));
   AOI22_X2 U_dsdc_U1776 (.ZN(U_dsdc_n1827), 
	.B2(U_dsdc_bm_bank_age_1__3_), 
	.B1(U_dsdc_n1839), 
	.A2(U_dsdc_n1840), 
	.A1(U_dsdc_bm_bank_age_2__3_));
   OAI21_X2 U_dsdc_U1775 (.ZN(U_dsdc_n1828), 
	.B2(U_dsdc_n284), 
	.B1(U_dsdc_n1841), 
	.A(U_dsdc_n1827));
   AOI21_X2 U_dsdc_U1774 (.ZN(U_dsdc_n1953), 
	.B2(U_dsdc_bm_bank_age_0__3_), 
	.B1(U_dsdc_n1842), 
	.A(U_dsdc_n1828));
   AOI22_X2 U_dsdc_U1773 (.ZN(U_dsdc_n1829), 
	.B2(U_dsdc_bm_bank_age_1__1_), 
	.B1(U_dsdc_n1839), 
	.A2(U_dsdc_n1840), 
	.A1(U_dsdc_bm_bank_age_2__1_));
   AOI21_X2 U_dsdc_U1772 (.ZN(U_dsdc_n1944), 
	.B2(U_dsdc_bm_bank_age_0__1_), 
	.B1(U_dsdc_n1842), 
	.A(U_dsdc_n1830));
   AOI22_X2 U_dsdc_U1771 (.ZN(U_dsdc_n1831), 
	.B2(U_dsdc_bm_bank_age_1__0_), 
	.B1(U_dsdc_n1839), 
	.A2(U_dsdc_n1840), 
	.A1(U_dsdc_bm_bank_age_2__0_));
   AOI21_X2 U_dsdc_U1770 (.ZN(U_dsdc_n1833), 
	.B2(U_dsdc_bm_bank_age_0__0_), 
	.B1(U_dsdc_n1842), 
	.A(U_dsdc_n1832));
   NOR2_X2 U_dsdc_U1769 (.ZN(U_dsdc_n1945), 
	.A2(U_dsdc_n1833), 
	.A1(U_dsdc_n1944));
   NOR2_X2 U_dsdc_U1768 (.ZN(U_dsdc_n1911), 
	.A2(U_dsdc_n308), 
	.A1(U_dsdc_n477));
   NAND2_X2 U_dsdc_U1767 (.ZN(U_dsdc_n1943), 
	.A2(U_dsdc_n1833), 
	.A1(U_dsdc_n1944));
   AOI22_X2 U_dsdc_U1766 (.ZN(U_dsdc_n1834), 
	.B2(U_dsdc_n1943), 
	.B1(U_dsdc_n178), 
	.A2(U_dsdc_n1951), 
	.A1(U_dsdc_n336));
   OAI221_X2 U_dsdc_U1765 (.ZN(U_dsdc_n1836), 
	.C2(U_dsdc_n1944), 
	.C1(U_dsdc_bm_bank_age_2__0_), 
	.B2(U_dsdc_bm_bank_age_2__1_), 
	.B1(U_dsdc_bm_bank_age_2__0_), 
	.A(U_dsdc_n1834));
   AOI22_X2 U_dsdc_U1762 (.ZN(U_dsdc_n1844), 
	.B2(U_dsdc_bm_bank_age_1__4_), 
	.B1(U_dsdc_n1839), 
	.A2(U_dsdc_n1840), 
	.A1(U_dsdc_bm_bank_age_2__4_));
   AOI22_X2 U_dsdc_U1761 (.ZN(U_dsdc_n1843), 
	.B2(U_dsdc_bm_bank_age_3__4_), 
	.B1(U_dsdc_n476), 
	.A2(U_dsdc_n1842), 
	.A1(U_dsdc_bm_bank_age_0__4_));
   NAND2_X2 U_dsdc_U1760 (.ZN(U_dsdc_n1954), 
	.A2(U_dsdc_n1843), 
	.A1(U_dsdc_n1844));
   NAND3_X2 U_dsdc_U1759 (.ZN(U_dsdc_n1856), 
	.A3(U_dsdc_n1849), 
	.A2(FE_PHN958_U_dsdc_n353), 
	.A1(U_dsdc_n178));
   NOR3_X2 U_dsdc_U1758 (.ZN(U_dsdc_n1961), 
	.A3(U_dsdc_n2082), 
	.A2(U_dsdc_n1846), 
	.A1(U_dsdc_r_bm_close_all));
   AOI21_X2 U_dsdc_U1757 (.ZN(U_dsdc_n1855), 
	.B2(U_dsdc_bm_bank_age_2__0_), 
	.B1(U_dsdc_bm_bank_age_2__1_), 
	.A(U_dsdc_n1860));
   AOI211_X2 U_dsdc_U1756 (.ZN(U_dsdc_n1858), 
	.C2(U_dsdc_n1856), 
	.C1(U_dsdc_n1867), 
	.B(U_dsdc_n1855), 
	.A(U_dsdc_n1961));
   OAI221_X2 U_dsdc_U1755 (.ZN(U_dsdc_n1865), 
	.C2(U_dsdc_n1859), 
	.C1(U_dsdc_n336), 
	.B2(U_dsdc_n1860), 
	.B1(U_dsdc_bm_bank_age_2__2_), 
	.A(U_dsdc_n1858));
   AOI221_X2 U_dsdc_U1754 (.ZN(U_dsdc_n1870), 
	.C2(U_dsdc_n459), 
	.C1(U_dsdc_n1866), 
	.B2(U_dsdc_bm_bank_age_2__3_), 
	.B1(U_dsdc_n1867), 
	.A(U_dsdc_n1865));
   NOR2_X2 U_dsdc_U1753 (.ZN(U_dsdc_n1868), 
	.A2(U_dsdc_n1861), 
	.A1(U_dsdc_n336));
   OAI21_X2 U_dsdc_U1752 (.ZN(U_dsdc_n213), 
	.B2(U_dsdc_n350), 
	.B1(U_dsdc_n1870), 
	.A(U_dsdc_n1869));
   AOI211_X2 U_dsdc_U1751 (.ZN(U_dsdc_n1019), 
	.C2(U_dsdc_bm_num_open_bank_3_), 
	.C1(U_dsdc_n1024), 
	.B(U_dsdc_n1022), 
	.A(U_dsdc_n1018));
   INV_X4 U_dsdc_U1750 (.ZN(U_dsdc_n296), 
	.A(U_dsdc_n1019));
   NOR3_X2 U_dsdc_U1749 (.ZN(U_dsdc_n1937), 
	.A3(U_dsdc_n1942), 
	.A2(U_dsdc_n383), 
	.A1(U_dsdc_r_bm_close_bank_1_));
   NOR3_X2 U_dsdc_U1748 (.ZN(U_dsdc_n1936), 
	.A3(U_dsdc_n383), 
	.A2(U_dsdc_n1941), 
	.A1(U_dsdc_r_bm_open_bank[1]));
   INV_X4 U_dsdc_U1747 (.ZN(U_dsdc_n1930), 
	.A(U_dsdc_n1936));
   INV_X4 U_dsdc_U1746 (.ZN(U_dsdc_n1929), 
	.A(U_dsdc_n1937));
   AOI22_X2 U_dsdc_U1745 (.ZN(U_dsdc_n1912), 
	.B2(U_dsdc_n1951), 
	.B1(U_dsdc_n337), 
	.A2(U_dsdc_n1943), 
	.A1(U_dsdc_n335));
   OAI221_X2 U_dsdc_U1744 (.ZN(U_dsdc_n1914), 
	.C2(U_dsdc_n1944), 
	.C1(U_dsdc_bm_bank_age_1__0_), 
	.B2(U_dsdc_bm_bank_age_1__1_), 
	.B1(U_dsdc_bm_bank_age_1__0_), 
	.A(U_dsdc_n1912));
   AOI221_X2 U_dsdc_U1743 (.ZN(U_dsdc_n1916), 
	.C2(U_dsdc_n1915), 
	.C1(U_dsdc_n1914), 
	.B2(U_dsdc_n1915), 
	.B1(U_dsdc_n1945), 
	.A(U_dsdc_n1913));
   AOI21_X2 U_dsdc_U1742 (.ZN(U_dsdc_n1917), 
	.B2(U_dsdc_n1953), 
	.B1(U_dsdc_bm_bank_age_1__3_), 
	.A(U_dsdc_n1916));
   NAND3_X2 U_dsdc_U1741 (.ZN(U_dsdc_n1926), 
	.A3(U_dsdc_n1920), 
	.A2(FE_PHN897_U_dsdc_n352), 
	.A1(U_dsdc_n335));
   AOI21_X2 U_dsdc_U1740 (.ZN(U_dsdc_n1925), 
	.B2(U_dsdc_bm_bank_age_1__0_), 
	.B1(U_dsdc_bm_bank_age_1__1_), 
	.A(U_dsdc_n1930));
   AOI211_X2 U_dsdc_U1739 (.ZN(U_dsdc_n1928), 
	.C2(U_dsdc_n1926), 
	.C1(U_dsdc_n1937), 
	.B(U_dsdc_n1925), 
	.A(U_dsdc_n1961));
   OAI221_X2 U_dsdc_U1738 (.ZN(U_dsdc_n1935), 
	.C2(U_dsdc_n1929), 
	.C1(U_dsdc_n337), 
	.B2(U_dsdc_n1930), 
	.B1(U_dsdc_bm_bank_age_1__2_), 
	.A(U_dsdc_n1928));
   AOI221_X2 U_dsdc_U1737 (.ZN(U_dsdc_n1940), 
	.C2(FE_PHN3077_U_dsdc_n460), 
	.C1(U_dsdc_n1936), 
	.B2(U_dsdc_bm_bank_age_1__3_), 
	.B1(U_dsdc_n1937), 
	.A(U_dsdc_n1935));
   NAND3_X2 U_dsdc_U1736 (.ZN(U_dsdc_n1931), 
	.A3(U_dsdc_n1936), 
	.A2(U_dsdc_bm_bank_age_1__0_), 
	.A1(U_dsdc_bm_bank_age_1__1_));
   NOR2_X2 U_dsdc_U1735 (.ZN(U_dsdc_n1938), 
	.A2(U_dsdc_n1931), 
	.A1(U_dsdc_n337));
   OAI21_X2 U_dsdc_U1734 (.ZN(U_dsdc_n227), 
	.B2(U_dsdc_n349), 
	.B1(U_dsdc_n1940), 
	.A(U_dsdc_n1939));
   NOR2_X2 U_dsdc_U1733 (.ZN(U_dsdc_n879), 
	.A2(U_dsdc_n1309), 
	.A1(U_dsdc_n903));
   NAND2_X2 U_dsdc_U1732 (.ZN(U_dsdc_n724), 
	.A2(U_dsdc_n758), 
	.A1(U_dsdc_n682));
   NAND2_X2 U_dsdc_U1731 (.ZN(U_dsdc_n650), 
	.A2(U_dsdc_n200), 
	.A1(U_dsdc_n457));
   NOR2_X2 U_dsdc_U1730 (.ZN(U_dsdc_n1638), 
	.A2(U_dsdc_term_cnt_1_), 
	.A1(U_dsdc_term_cnt_0_));
   INV_X4 U_dsdc_U1729 (.ZN(U_dsdc_n1640), 
	.A(U_dsdc_n1638));
   NOR3_X2 U_dsdc_U1728 (.ZN(U_dsdc_n1424), 
	.A3(U_dsdc_n1640), 
	.A2(U_dsdc_term_cnt_3_), 
	.A1(U_dsdc_n650));
   NAND2_X2 U_dsdc_U1727 (.ZN(U_dsdc_n1329), 
	.A2(U_dsdc_n309), 
	.A1(U_dsdc_n171));
   NOR2_X2 U_dsdc_U1726 (.ZN(U_dsdc_n1426), 
	.A2(U_dsdc_rp_cnt2_2_), 
	.A1(U_dsdc_n1329));
   NAND2_X2 U_dsdc_U1725 (.ZN(U_dsdc_n1871), 
	.A2(U_dsdc_n1426), 
	.A1(U_dsdc_n1424));
   INV_X4 U_dsdc_U1724 (.ZN(U_dsdc_n1423), 
	.A(U_dsdc_n1871));
   NAND3_X2 U_dsdc_U1723 (.ZN(U_dsdc_n1627), 
	.A3(U_dsdc_n1425), 
	.A2(U_dsdc_r_rw), 
	.A1(U_dsdc_n1423));
   INV_X4 U_dsdc_U1722 (.ZN(U_dsdc_n722), 
	.A(U_dsdc_n1627));
   NOR2_X2 U_dsdc_U1721 (.ZN(U_dsdc_n1293), 
	.A2(U_dsdc_n690), 
	.A1(U_dsdc_n692));
   INV_X4 U_dsdc_U1720 (.ZN(U_dsdc_n1556), 
	.A(U_dsdc_n1410));
   INV_X4 U_dsdc_U1719 (.ZN(U_dsdc_n673), 
	.A(U_dsdc_n936));
   NOR2_X2 U_dsdc_U1718 (.ZN(U_dsdc_n683), 
	.A2(U_dsdc_n904), 
	.A1(U_dsdc_n673));
   AOI21_X2 U_dsdc_U1717 (.ZN(U_dsdc_n1403), 
	.B2(U_dsdc_n724), 
	.B1(U_dsdc_n1060), 
	.A(U_dsdc_n683));
   NAND2_X2 U_dsdc_U1716 (.ZN(U_dsdc_n1629), 
	.A2(U_dsdc_access_cs_0_), 
	.A1(U_dsdc_n736));
   NOR2_X2 U_dsdc_U1715 (.ZN(U_dsdc_n728), 
	.A2(U_dsdc_n1633), 
	.A1(U_dsdc_n684));
   AOI21_X2 U_dsdc_U1714 (.ZN(U_dsdc_n686), 
	.B2(U_dsdc_n1423), 
	.B1(U_dsdc_n685), 
	.A(U_dsdc_n728));
   NOR2_X2 U_dsdc_U1713 (.ZN(U_dsdc_n1625), 
	.A2(U_dsdc_n1419), 
	.A1(U_dsdc_n686));
   NOR3_X2 U_dsdc_U1712 (.ZN(U_dsdc_n689), 
	.A3(U_dsdc_n688), 
	.A2(U_dsdc_n1258), 
	.A1(U_dsdc_n1559));
   AOI211_X2 U_dsdc_U1711 (.ZN(U_dsdc_n1560), 
	.C2(U_dsdc_wrapped_pop_flag), 
	.C1(U_dsdc_n865), 
	.B(U_dsdc_n689), 
	.A(U_dsdc_n1625));
   OAI221_X2 U_dsdc_U1710 (.ZN(U_dsdc_n1562), 
	.C2(U_dsdc_n1651), 
	.C1(U_dsdc_n1561), 
	.B2(U_dsdc_n1403), 
	.B1(U_dsdc_n1561), 
	.A(U_dsdc_n1560));
   NOR3_X2 U_dsdc_U1709 (.ZN(U_dsdc_n726), 
	.A3(U_dsdc_n1562), 
	.A2(U_dsdc_n1563), 
	.A1(U_dsdc_n1293));
   OAI211_X2 U_dsdc_U1708 (.ZN(ctl_burst_done), 
	.C2(U_dsdc_n181), 
	.C1(U_dsdc_n727), 
	.B(U_dsdc_n725), 
	.A(U_dsdc_n726));
   NOR2_X2 U_dsdc_U1707 (.ZN(U_dsdc_n1179), 
	.A2(U_dsdc_bm_rc_cnt_0__2_), 
	.A1(FE_PHN945_U_dsdc_n1175));
   NOR2_X2 U_dsdc_U1706 (.ZN(U_dsdc_n1180), 
	.A2(U_dsdc_n441), 
	.A1(U_dsdc_n1179));
   AOI21_X2 U_dsdc_U1705 (.ZN(U_dsdc_n1169), 
	.B2(debug_ad_row_addr[13]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1132));
   INV_X4 U_dsdc_U1704 (.ZN(U_dsdc_n1218), 
	.A(U_dsdc_n1169));
   AOI21_X2 U_dsdc_U1703 (.ZN(U_dsdc_n1170), 
	.B2(debug_ad_row_addr[3]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1115));
   INV_X4 U_dsdc_U1702 (.ZN(U_dsdc_n1222), 
	.A(U_dsdc_n1170));
   AOI21_X2 U_dsdc_U1701 (.ZN(U_dsdc_n1147), 
	.B2(debug_ad_row_addr[9]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1073));
   INV_X4 U_dsdc_U1700 (.ZN(U_dsdc_n1148), 
	.A(U_dsdc_n1147));
   AOI21_X2 U_dsdc_U1699 (.ZN(U_dsdc_n1171), 
	.B2(debug_ad_row_addr[2]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1116));
   INV_X4 U_dsdc_U1698 (.ZN(U_dsdc_n1223), 
	.A(U_dsdc_n1171));
   NAND2_X2 U_dsdc_U1697 (.ZN(U_dsdc_n1027), 
	.A2(FE_PHN1148_U_dsdc_r_row_addr_10_), 
	.A1(U_dsdc_n1109));
   OAI21_X2 U_dsdc_U1696 (.ZN(U_dsdc_n1146), 
	.B2(U_dsdc_n1028), 
	.B1(U_dsdc_n1112), 
	.A(U_dsdc_n1027));
   NAND2_X2 U_dsdc_U1695 (.ZN(U_dsdc_n1110), 
	.A2(FE_PHN1147_U_dsdc_r_row_addr_4_), 
	.A1(U_dsdc_n1109));
   OAI21_X2 U_dsdc_U1694 (.ZN(U_dsdc_n1221), 
	.B2(U_dsdc_n1111), 
	.B1(U_dsdc_n1112), 
	.A(U_dsdc_n1110));
   AOI21_X2 U_dsdc_U1693 (.ZN(U_dsdc_n1144), 
	.B2(debug_ad_row_addr[11]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1069));
   INV_X4 U_dsdc_U1692 (.ZN(U_dsdc_n1145), 
	.A(U_dsdc_n1144));
   AOI21_X2 U_dsdc_U1691 (.ZN(U_dsdc_n1172), 
	.B2(debug_ad_row_addr[1]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1117));
   INV_X4 U_dsdc_U1690 (.ZN(U_dsdc_n1224), 
	.A(U_dsdc_n1172));
   NAND2_X2 U_dsdc_U1689 (.ZN(U_dsdc_n1075), 
	.A2(FE_PHN1151_U_dsdc_r_row_addr_8_), 
	.A1(U_dsdc_n1109));
   OAI21_X2 U_dsdc_U1688 (.ZN(U_dsdc_n1149), 
	.B2(U_dsdc_n1076), 
	.B1(U_dsdc_n1112), 
	.A(U_dsdc_n1075));
   AOI21_X2 U_dsdc_U1687 (.ZN(U_dsdc_n1150), 
	.B2(debug_ad_row_addr[7]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1095));
   INV_X4 U_dsdc_U1686 (.ZN(U_dsdc_n1151), 
	.A(U_dsdc_n1150));
   NAND2_X2 U_dsdc_U1685 (.ZN(U_dsdc_n1103), 
	.A2(FE_PHN1152_U_dsdc_r_row_addr_5_), 
	.A1(U_dsdc_n1109));
   OAI21_X2 U_dsdc_U1684 (.ZN(U_dsdc_n1220), 
	.B2(U_dsdc_n1104), 
	.B1(U_dsdc_n1112), 
	.A(U_dsdc_n1103));
   NAND2_X2 U_dsdc_U1683 (.ZN(U_dsdc_n1097), 
	.A2(FE_PHN1146_U_dsdc_r_row_addr_6_), 
	.A1(U_dsdc_n1109));
   OAI21_X2 U_dsdc_U1682 (.ZN(U_dsdc_n1219), 
	.B2(U_dsdc_n1098), 
	.B1(U_dsdc_n1112), 
	.A(U_dsdc_n1097));
   NAND2_X2 U_dsdc_U1681 (.ZN(U_dsdc_n1058), 
	.A2(FE_PHN1149_U_dsdc_r_row_addr_12_), 
	.A1(U_dsdc_n1109));
   OAI21_X2 U_dsdc_U1680 (.ZN(U_dsdc_n1143), 
	.B2(U_addrdec_n241), 
	.B1(U_dsdc_n1112), 
	.A(U_dsdc_n1058));
   AOI21_X2 U_dsdc_U1679 (.ZN(U_dsdc_n1168), 
	.B2(debug_ad_row_addr[14]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1134));
   INV_X4 U_dsdc_U1678 (.ZN(U_dsdc_n1217), 
	.A(U_dsdc_n1168));
   AOI21_X2 U_dsdc_U1677 (.ZN(U_dsdc_n1173), 
	.B2(debug_ad_row_addr[0]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1122));
   INV_X4 U_dsdc_U1676 (.ZN(U_dsdc_n1225), 
	.A(U_dsdc_n1173));
   AOI21_X2 U_dsdc_U1675 (.ZN(U_dsdc_n1167), 
	.B2(debug_ad_row_addr[15]), 
	.B1(U_dsdc_n1388), 
	.A(U_dsdc_n1137));
   INV_X4 U_dsdc_U1674 (.ZN(U_dsdc_n1216), 
	.A(U_dsdc_n1167));
   NOR2_X2 U_dsdc_U1673 (.ZN(U_dsdc_n1234), 
	.A2(FE_PHN1219_U_dsdc_bm_rc_cnt_3__2_), 
	.A1(U_dsdc_n1228));
   NOR2_X2 U_dsdc_U1672 (.ZN(U_dsdc_n1235), 
	.A2(U_dsdc_n442), 
	.A1(U_dsdc_n1234));
   OAI21_X2 U_dsdc_U1671 (.ZN(U_dsdc_n1014), 
	.B2(U_dsdc_n1012), 
	.B1(U_dsdc_n1013), 
	.A(U_dsdc_n338));
   OAI21_X2 U_dsdc_U1670 (.ZN(U_dsdc_n295), 
	.B2(U_dsdc_n338), 
	.B1(U_dsdc_n1016), 
	.A(U_dsdc_n1014));
   NOR2_X2 U_dsdc_U1667 (.ZN(U_dsdc_n967), 
	.A2(U_dsdc_n1163), 
	.A1(U_dsdc_n710));
   NOR2_X2 U_dsdc_U1665 (.ZN(U_dsdc_n1358), 
	.A2(U_dsdc_n1293), 
	.A1(U_dsdc_n691));
   NOR2_X2 U_dsdc_U1664 (.ZN(U_dsdc_n693), 
	.A2(U_dsdc_n871), 
	.A1(U_dsdc_n866));
   NAND2_X2 U_dsdc_U1663 (.ZN(U_dsdc_n1802), 
	.A2(U_dsdc_n693), 
	.A1(U_dsdc_n1358));
   NAND2_X2 U_dsdc_U1662 (.ZN(U_dsdc_n1349), 
	.A2(U_dsdc_n1633), 
	.A1(U_dsdc_n741));
   NOR2_X2 U_dsdc_U1661 (.ZN(U_dsdc_n1041), 
	.A2(n21), 
	.A1(U_dsdc_n914));
   AOI21_X2 U_dsdc_U1660 (.ZN(U_dsdc_n945), 
	.B2(U_dsdc_n712), 
	.B1(U_dsdc_n1348), 
	.A(U_dsdc_n711));
   NAND2_X2 U_dsdc_U1658 (.ZN(U_dsdc_n880), 
	.A2(U_dsdc_n714), 
	.A1(U_dsdc_n1437));
   NAND2_X2 U_dsdc_U1657 (.ZN(U_dsdc_n1033), 
	.A2(U_dsdc_n883), 
	.A1(U_dsdc_n1041));
   NOR2_X2 U_dsdc_U1656 (.ZN(U_dsdc_n960), 
	.A2(U_dsdc_n2013), 
	.A1(U_dsdc_n1033));
   NAND2_X2 U_dsdc_U1655 (.ZN(U_dsdc_n890), 
	.A2(U_dsdc_n886), 
	.A1(U_dsdc_n887));
   NAND2_X2 U_dsdc_U1654 (.ZN(U_dsdc_n896), 
	.A2(U_cr_n56), 
	.A1(FE_PHN2909_U_dsdc_n1436));
   NAND2_X2 U_dsdc_U1653 (.ZN(U_dsdc_n889), 
	.A2(n84), 
	.A1(U_cr_n39));
   NOR2_X2 U_dsdc_U1652 (.ZN(U_dsdc_n1032), 
	.A2(U_dsdc_n889), 
	.A1(FE_PHN678_U_dsdc_n896));
   INV_X4 U_dsdc_U1651 (.ZN(U_dsdc_n892), 
	.A(U_dsdc_n1032));
   NOR2_X2 U_dsdc_U1650 (.ZN(U_dsdc_n1042), 
	.A2(U_dsdc_n1031), 
	.A1(U_dsdc_n892));
   AOI21_X2 U_dsdc_U1649 (.ZN(U_dsdc_n1310), 
	.B2(U_dsdc_n1042), 
	.B1(U_dsdc_n890), 
	.A(U_dsdc_n165));
   NAND2_X2 U_dsdc_U1648 (.ZN(U_dsdc_n893), 
	.A2(U_dsdc_n891), 
	.A1(U_dsdc_n892));
   NAND2_X2 U_dsdc_U1647 (.ZN(U_dsdc_n1298), 
	.A2(U_dsdc_n893), 
	.A1(U_dsdc_n1310));
   NAND2_X2 U_dsdc_U1646 (.ZN(U_dsdc_n1252), 
	.A2(U_dsdc_n1411), 
	.A1(U_dsdc_n1298));
   NAND2_X2 U_dsdc_U1645 (.ZN(U_dsdc_n1979), 
	.A2(U_dsdc_n881), 
	.A1(U_dsdc_n1299));
   NAND3_X2 U_dsdc_U1644 (.ZN(U_dsdc_n1374), 
	.A3(U_dsdc_n1979), 
	.A2(U_dsdc_n1252), 
	.A1(U_dsdc_n894));
   NOR2_X2 U_dsdc_U1642 (.ZN(U_dsdc_n596), 
	.A2(U_dsdc_row_cnt_12_), 
	.A1(U_dsdc_row_cnt_14_));
   NAND3_X2 U_dsdc_U1641 (.ZN(U_dsdc_n597), 
	.A3(U_dsdc_n426), 
	.A2(U_dsdc_n197), 
	.A1(U_dsdc_n596));
   NOR2_X2 U_dsdc_U1640 (.ZN(U_dsdc_n1468), 
	.A2(U_dsdc_n1490), 
	.A1(U_dsdc_n1485));
   INV_X4 U_dsdc_U1639 (.ZN(U_dsdc_n1506), 
	.A(U_dsdc_n1435));
   NOR2_X2 U_dsdc_U1638 (.ZN(U_dsdc_n1467), 
	.A2(U_dsdc_n1451), 
	.A1(U_dsdc_n1506));
   AOI22_X2 U_dsdc_U1637 (.ZN(U_dsdc_n1492), 
	.B2(U_cr_n39), 
	.B1(U_dsdc_n1467), 
	.A2(U_dsdc_n1468), 
	.A1(U_dsdc_n1478));
   NOR2_X2 U_dsdc_U1636 (.ZN(U_dsdc_n1489), 
	.A2(U_dsdc_n1490), 
	.A1(U_dsdc_n1451));
   INV_X4 U_dsdc_U1635 (.ZN(U_dsdc_n1521), 
	.A(U_dsdc_n1512));
   NOR2_X2 U_dsdc_U1634 (.ZN(U_dsdc_n1519), 
	.A2(U_dsdc_n1521), 
	.A1(U_dsdc_operation_cs_1_));
   NOR2_X2 U_dsdc_U1633 (.ZN(U_dsdc_n1450), 
	.A2(U_dsdc_operation_cs_2_), 
	.A1(U_dsdc_operation_cs_3_));
   NAND2_X2 U_dsdc_U1632 (.ZN(U_dsdc_n1454), 
	.A2(U_dsdc_n432), 
	.A1(U_dsdc_n1450));
   NOR2_X2 U_dsdc_U1631 (.ZN(U_dsdc_n1498), 
	.A2(U_dsdc_n1454), 
	.A1(U_dsdc_n1490));
   NOR2_X2 U_dsdc_U1629 (.ZN(U_dsdc_n1534), 
	.A2(U_dsdc_n1485), 
	.A1(U_dsdc_n1506));
   NOR2_X2 U_dsdc_U1628 (.ZN(ctl_sd_in_sf_mode), 
	.A2(U_dsdc_n1455), 
	.A1(U_dsdc_n1451));
   NOR2_X2 U_dsdc_U1627 (.ZN(U_dsdc_n2060), 
	.A2(ctl_sd_in_sf_mode), 
	.A1(U_dsdc_n1534));
   NOR2_X2 U_dsdc_U1626 (.ZN(U_dsdc_n2064), 
	.A2(U_dsdc_n1522), 
	.A1(U_dsdc_n1485));
   NOR2_X2 U_dsdc_U1625 (.ZN(U_dsdc_n1526), 
	.A2(U_dsdc_n1506), 
	.A1(U_dsdc_n1454));
   INV_X4 U_dsdc_U1624 (.ZN(U_dsdc_n1587), 
	.A(U_dsdc_n1584));
   NOR2_X2 U_dsdc_U1623 (.ZN(U_dsdc_n1577), 
	.A2(U_dsdc_n1587), 
	.A1(U_dsdc_rcar_cnt1_3_));
   NOR2_X2 U_dsdc_U1622 (.ZN(U_dsdc_n1574), 
	.A2(U_dsdc_n1468), 
	.A1(U_dsdc_n1467));
   NAND2_X2 U_dsdc_U1621 (.ZN(U_dsdc_n2051), 
	.A2(U_dsdc_n642), 
	.A1(U_dsdc_n1434));
   NOR2_X2 U_dsdc_U1620 (.ZN(U_dsdc_n1565), 
	.A2(U_dsdc_n2051), 
	.A1(U_dsdc_n1577));
   NOR2_X2 U_dsdc_U1619 (.ZN(U_dsdc_n1432), 
	.A2(U_dsdc_n1522), 
	.A1(U_dsdc_n1454));
   NAND2_X2 U_dsdc_U1618 (.ZN(U_dsdc_n1510), 
	.A2(U_dsdc_n1434), 
	.A1(U_dsdc_n661));
   NOR2_X2 U_dsdc_U1617 (.ZN(U_dsdc_n1535), 
	.A2(U_dsdc_n1524), 
	.A1(U_dsdc_n1432));
   NAND3_X2 U_dsdc_U1616 (.ZN(U_dsdc_n1509), 
	.A3(U_dsdc_n169), 
	.A2(U_dsdc_n427), 
	.A1(U_dsdc_n198));
   NOR2_X2 U_dsdc_U1615 (.ZN(U_dsdc_n1617), 
	.A2(U_dsdc_n1431), 
	.A1(U_dsdc_n1535));
   NOR4_X2 U_dsdc_U1614 (.ZN(U_dsdc_n1740), 
	.A4(U_dsdc_xsr_cnt_2_), 
	.A3(FE_PHN1030_U_dsdc_xsr_cnt_3_), 
	.A2(FE_PHN1033_U_dsdc_xsr_cnt_1_), 
	.A1(U_dsdc_xsr_cnt_0_));
   INV_X4 U_dsdc_U1613 (.ZN(U_dsdc_n1737), 
	.A(U_dsdc_n1740));
   NOR3_X2 U_dsdc_U1612 (.ZN(U_dsdc_n1736), 
	.A3(U_dsdc_n1737), 
	.A2(U_dsdc_xsr_cnt_5_), 
	.A1(U_dsdc_xsr_cnt_4_));
   NAND2_X2 U_dsdc_U1611 (.ZN(U_dsdc_n1727), 
	.A2(FE_PHN816_U_dsdc_n359), 
	.A1(U_dsdc_n1736));
   NOR2_X2 U_dsdc_U1610 (.ZN(U_dsdc_n1536), 
	.A2(U_dsdc_n1522), 
	.A1(U_dsdc_n1451));
   NOR2_X2 U_dsdc_U1609 (.ZN(U_dsdc_n1500), 
	.A2(U_dsdc_n1452), 
	.A1(U_dsdc_n1728));
   NAND2_X2 U_dsdc_U1606 (.ZN(U_dsdc_n1491), 
	.A2(U_dsdc_n429), 
	.A1(U_dsdc_n199));
   INV_X4 U_dsdc_U1605 (.ZN(U_dsdc_n1430), 
	.A(FE_PHN791_U_dsdc_n1491));
   NAND2_X2 U_dsdc_U1603 (.ZN(U_dsdc_n2058), 
	.A2(U_dsdc_n661), 
	.A1(U_dsdc_n662));
   NAND3_X2 U_dsdc_U1599 (.ZN(U_dsdc_n899), 
	.A3(U_dsdc_n847), 
	.A2(U_dsdc_n848), 
	.A1(U_dsdc_n913));
   NAND2_X2 U_dsdc_U1591 (.ZN(U_dsdc_n1974), 
	.A2(U_dsdc_n710), 
	.A1(U_dsdc_n725));
   NAND2_X2 U_dsdc_U1587 (.ZN(U_dsdc_n1372), 
	.A2(U_dsdc_n1438), 
	.A1(U_dsdc_n1557));
   INV_X4 U_dsdc_U1586 (.ZN(U_dsdc_n1043), 
	.A(U_dsdc_n1372));
   AOI21_X2 U_dsdc_U1585 (.ZN(U_dsdc_n1367), 
	.B2(U_dsdc_n703), 
	.B1(U_dsdc_n1061), 
	.A(U_dsdc_n2071));
   OAI21_X2 U_dsdc_U1581 (.ZN(U_dsdc_n958), 
	.B2(U_dsdc_n967), 
	.B1(U_dsdc_r_rw), 
	.A(U_dsdc_n1974));
   NOR4_X2 U_dsdc_U1579 (.ZN(U_dsdc_n1564), 
	.A4(U_dsdc_num_init_ref_cnt_3_), 
	.A3(U_dsdc_num_init_ref_cnt_2_), 
	.A2(FE_PHN843_U_dsdc_num_init_ref_cnt_1_), 
	.A1(U_dsdc_num_init_ref_cnt_0_));
   INV_X4 U_dsdc_U1578 (.ZN(U_dsdc_n1433), 
	.A(U_dsdc_n2051));
   NOR2_X2 U_dsdc_U1577 (.ZN(U_dsdc_n1466), 
	.A2(U_dsdc_n1470), 
	.A1(cr_do_initialize));
   NAND2_X2 U_dsdc_U1576 (.ZN(U_dsdc_n2052), 
	.A2(U_dsdc_n1466), 
	.A1(FE_PHN2909_U_dsdc_n1436));
   NOR2_X2 U_dsdc_U1575 (.ZN(U_dsdc_n1758), 
	.A2(U_cr_n39), 
	.A1(U_dsdc_n2052));
   NAND2_X2 U_dsdc_U1574 (.ZN(U_dsdc_n1501), 
	.A2(U_dsdc_n1509), 
	.A1(U_dsdc_n1432));
   NOR2_X2 U_dsdc_U1573 (.ZN(U_dsdc_n1581), 
	.A2(U_dsdc_n1455), 
	.A1(U_dsdc_n1485));
   NAND2_X2 U_dsdc_U1570 (.ZN(U_dsdc_n956), 
	.A2(U_dsdc_n934), 
	.A1(U_dsdc_n2071));
   NOR4_X2 U_dsdc_U1569 (.ZN(U_dsdc_n959), 
	.A4(U_dsdc_n1425), 
	.A3(U_dsdc_n1349), 
	.A2(U_dsdc_n956), 
	.A1(U_dsdc_n1802));
   NAND4_X2 U_dsdc_U1568 (.ZN(U_dsdc_n963), 
	.A4(U_dsdc_n957), 
	.A3(U_dsdc_n958), 
	.A2(U_dsdc_n959), 
	.A1(U_dsdc_n972));
   NOR3_X2 U_dsdc_U1567 (.ZN(U_dsdc_n1907), 
	.A3(U_dsdc_n1942), 
	.A2(U_dsdc_n396), 
	.A1(U_dsdc_r_bm_close_bank_3_));
   NOR3_X2 U_dsdc_U1566 (.ZN(U_dsdc_n1906), 
	.A3(U_dsdc_n396), 
	.A2(U_dsdc_n1941), 
	.A1(U_dsdc_r_bm_open_bank[3]));
   INV_X4 U_dsdc_U1565 (.ZN(U_dsdc_n1900), 
	.A(U_dsdc_n1906));
   INV_X4 U_dsdc_U1564 (.ZN(U_dsdc_n1899), 
	.A(U_dsdc_n1907));
   AOI22_X2 U_dsdc_U1563 (.ZN(U_dsdc_n1882), 
	.B2(U_dsdc_n1951), 
	.B1(U_dsdc_n303), 
	.A2(U_dsdc_n1943), 
	.A1(U_dsdc_n302));
   OAI221_X2 U_dsdc_U1562 (.ZN(U_dsdc_n1884), 
	.C2(U_dsdc_n1944), 
	.C1(U_dsdc_bm_bank_age_3__0_), 
	.B2(U_dsdc_bm_bank_age_3__1_), 
	.B1(U_dsdc_bm_bank_age_3__0_), 
	.A(U_dsdc_n1882));
   AOI221_X2 U_dsdc_U1561 (.ZN(U_dsdc_n1886), 
	.C2(U_dsdc_n1885), 
	.C1(U_dsdc_n1884), 
	.B2(U_dsdc_n1885), 
	.B1(U_dsdc_n1945), 
	.A(U_dsdc_n1883));
   AOI21_X2 U_dsdc_U1560 (.ZN(U_dsdc_n1887), 
	.B2(U_dsdc_n1953), 
	.B1(U_dsdc_bm_bank_age_3__3_), 
	.A(U_dsdc_n1886));
   AOI222_X1 U_dsdc_U1559 (.ZN(U_dsdc_n1890), 
	.C2(U_dsdc_n1954), 
	.C1(U_dsdc_n351), 
	.B2(U_dsdc_n1954), 
	.B1(U_dsdc_n1887), 
	.A2(U_dsdc_n351), 
	.A1(U_dsdc_n1887));
   NAND3_X2 U_dsdc_U1558 (.ZN(U_dsdc_n1896), 
	.A3(U_dsdc_n1890), 
	.A2(U_dsdc_n304), 
	.A1(U_dsdc_n302));
   AOI21_X2 U_dsdc_U1557 (.ZN(U_dsdc_n1895), 
	.B2(U_dsdc_bm_bank_age_3__0_), 
	.B1(U_dsdc_bm_bank_age_3__1_), 
	.A(U_dsdc_n1900));
   AOI211_X2 U_dsdc_U1556 (.ZN(U_dsdc_n1898), 
	.C2(U_dsdc_n1896), 
	.C1(U_dsdc_n1907), 
	.B(U_dsdc_n1895), 
	.A(U_dsdc_n1961));
   OAI221_X2 U_dsdc_U1555 (.ZN(U_dsdc_n1905), 
	.C2(U_dsdc_n1899), 
	.C1(U_dsdc_n303), 
	.B2(U_dsdc_n1900), 
	.B1(U_dsdc_bm_bank_age_3__2_), 
	.A(U_dsdc_n1898));
   AOI221_X2 U_dsdc_U1554 (.ZN(U_dsdc_n1910), 
	.C2(U_dsdc_n284), 
	.C1(U_dsdc_n1906), 
	.B2(U_dsdc_bm_bank_age_3__3_), 
	.B1(U_dsdc_n1907), 
	.A(U_dsdc_n1905));
   NOR2_X2 U_dsdc_U1553 (.ZN(U_dsdc_n1908), 
	.A2(U_dsdc_n1901), 
	.A1(U_dsdc_n303));
   AOI22_X2 U_dsdc_U1552 (.ZN(U_dsdc_n222), 
	.B2(U_dsdc_n351), 
	.B1(U_dsdc_n1909), 
	.A2(U_dsdc_n1910), 
	.A1(U_dsdc_bm_bank_age_3__4_));
   NOR2_X2 U_dsdc_U1551 (.ZN(U_dsdc_n1207), 
	.A2(FE_PHN1222_U_dsdc_bm_rc_cnt_2__2_), 
	.A1(U_dsdc_n1203));
   NOR2_X2 U_dsdc_U1550 (.ZN(U_dsdc_n1208), 
	.A2(U_dsdc_n439), 
	.A1(U_dsdc_n1207));
   NOR2_X2 U_dsdc_U1549 (.ZN(U_dsdc_n1193), 
	.A2(FE_PHN1221_U_dsdc_bm_rc_cnt_1__2_), 
	.A1(U_dsdc_n1189));
   NOR2_X2 U_dsdc_U1548 (.ZN(U_dsdc_n1194), 
	.A2(U_dsdc_n438), 
	.A1(U_dsdc_n1193));
   NAND2_X2 U_dsdc_U1547 (.ZN(U_dsdc_n307), 
	.A2(U_dsdc_n604), 
	.A1(U_dsdc_n1166));
   INV_X4 U_dsdc_U1546 (.ZN(U_dsdc_n621), 
	.A(U_dsdc_n307));
   INV_X4 U_dsdc_U1543 (.ZN(U_dsdc_n1009), 
	.A(U_dsdc_n1011));
   OAI211_X2 U_dsdc_U1542 (.ZN(U_dsdc_n294), 
	.C2(U_dsdc_n180), 
	.C1(U_dsdc_n1009), 
	.B(U_dsdc_n1008), 
	.A(U_dsdc_n1017));
   NAND2_X2 U_dsdc_U1541 (.ZN(U_dsdc_n1289), 
	.A2(U_dsdc_n1032), 
	.A1(U_dsdc_n960));
   NAND2_X2 U_dsdc_U1538 (.ZN(U_dsdc_n1051), 
	.A2(U_dsdc_n1044), 
	.A1(U_dsdc_n1320));
   NAND2_X2 U_dsdc_U1537 (.ZN(U_dsdc_n1314), 
	.A2(FE_PHN1887_U_dsdc_n166), 
	.A1(U_dsdc_n619));
   AOI21_X2 U_dsdc_U1527 (.ZN(U_dsdc_n1409), 
	.B2(U_dsdc_n672), 
	.B1(U_dsdc_n1413), 
	.A(U_dsdc_n669));
   INV_X4 U_dsdc_U1525 (.ZN(U_dsdc_n1260), 
	.A(U_dsdc_n1268));
   NOR2_X2 U_dsdc_U1513 (.ZN(U_dsdc_n1482), 
	.A2(U_dsdc_t_xp_cnt_0_), 
	.A1(U_dsdc_t_xp_cnt_1_));
   INV_X4 U_dsdc_U1512 (.ZN(U_dsdc_n2057), 
	.A(U_dsdc_n1534));
   AOI21_X2 U_dsdc_U1511 (.ZN(U_dsdc_n1540), 
	.B2(U_dsdc_n1465), 
	.B1(U_dsdc_n1466), 
	.A(U_dsdc_n1581));
   INV_X4 U_dsdc_U1510 (.ZN(U_dsdc_n2066), 
	.A(U_dsdc_n1467));
   INV_X4 U_dsdc_U1509 (.ZN(U_dsdc_n2059), 
	.A(U_dsdc_n1468));
   OAI22_X2 U_dsdc_U1508 (.ZN(U_dsdc_n1472), 
	.B2(U_dsdc_n1469), 
	.B1(U_dsdc_n1470), 
	.A2(U_dsdc_n1471), 
	.A1(U_dsdc_n1482));
   NOR4_X2 U_dsdc_U1507 (.ZN(U_dsdc_n1503), 
	.A4(U_dsdc_n1472), 
	.A3(U_dsdc_n362), 
	.A2(U_dsdc_n1576), 
	.A1(U_dsdc_n1800));
   NOR4_X2 U_dsdc_U1506 (.ZN(U_dsdc_n1708), 
	.A4(FE_PHN1062_U_dsdc_init_cnt_3_), 
	.A3(U_dsdc_init_cnt_2_), 
	.A2(U_dsdc_init_cnt_1_), 
	.A1(U_dsdc_init_cnt_0_));
   NOR3_X2 U_dsdc_U1505 (.ZN(U_dsdc_n1701), 
	.A3(U_dsdc_n1704), 
	.A2(U_dsdc_init_cnt_4_), 
	.A1(FE_PHN971_U_dsdc_init_cnt_5_));
   NOR3_X2 U_dsdc_U1504 (.ZN(U_dsdc_n1694), 
	.A3(U_dsdc_n1697), 
	.A2(U_dsdc_init_cnt_6_), 
	.A1(FE_PHN1031_U_dsdc_init_cnt_7_));
   NOR3_X2 U_dsdc_U1503 (.ZN(U_dsdc_n1687), 
	.A3(U_dsdc_n1690), 
	.A2(U_dsdc_init_cnt_8_), 
	.A1(FE_PHN1032_U_dsdc_init_cnt_9_));
   NOR3_X2 U_dsdc_U1502 (.ZN(U_dsdc_n1679), 
	.A3(U_dsdc_n1683), 
	.A2(FE_PHN3268_U_dsdc_init_cnt_10_), 
	.A1(FE_PHN970_U_dsdc_init_cnt_11_));
   NOR2_X2 U_dsdc_U1501 (.ZN(U_dsdc_n481), 
	.A2(U_dsdc_init_cnt_12_), 
	.A1(U_dsdc_init_cnt_13_));
   NAND2_X2 U_dsdc_U1500 (.ZN(U_dsdc_n482), 
	.A2(U_dsdc_n481), 
	.A1(U_dsdc_n1679));
   AOI211_X2 U_dsdc_U1499 (.ZN(U_dsdc_n1475), 
	.C2(U_dsdc_n1473), 
	.C1(U_dsdc_n1474), 
	.B(U_dsdc_n1522), 
	.A(U_dsdc_n1521));
   AOI211_X2 U_dsdc_U1498 (.ZN(U_dsdc_n1504), 
	.C2(U_dsdc_n1675), 
	.C1(U_dsdc_n1526), 
	.B(U_dsdc_n1475), 
	.A(U_dsdc_n2064));
   AOI21_X2 U_dsdc_U1497 (.ZN(U_dsdc_n1477), 
	.B2(U_dsdc_n1476), 
	.B1(U_dsdc_n1489), 
	.A(U_dsdc_n1536));
   NAND3_X2 U_dsdc_U1496 (.ZN(U_dsdc_n1533), 
	.A3(U_dsdc_n1477), 
	.A2(U_dsdc_n1504), 
	.A1(U_dsdc_n1503));
   INV_X4 U_dsdc_U1495 (.ZN(U_dsdc_n1532), 
	.A(ctl_sd_in_sf_mode));
   OAI21_X2 U_dsdc_U1494 (.ZN(U_dsdc_n1523), 
	.B2(U_dsdc_n2056), 
	.B1(U_dsdc_n2057), 
	.A(U_dsdc_n1532));
   NAND2_X2 U_dsdc_U1493 (.ZN(U_dsdc_n1537), 
	.A2(U_dsdc_n1482), 
	.A1(U_dsdc_n1479));
   OAI22_X2 U_dsdc_U1492 (.ZN(U_dsdc_n1525), 
	.B2(U_dsdc_n1537), 
	.B1(n84), 
	.A2(U_dsdc_n2062), 
	.A1(U_dsdc_n2066));
   AOI221_X2 U_dsdc_U1491 (.ZN(U_dsdc_n1481), 
	.C2(U_dsdc_operation_cs_3_), 
	.C1(U_dsdc_n1523), 
	.B2(U_dsdc_operation_cs_3_), 
	.B1(U_dsdc_n1533), 
	.A(U_dsdc_n1525));
   NAND2_X2 U_dsdc_U1490 (.ZN(U_dsdc_n1480), 
	.A2(U_dsdc_n1433), 
	.A1(U_dsdc_n644));
   NAND4_X2 U_dsdc_U1489 (.ZN(U_dsdc_n2094), 
	.A4(U_dsdc_n1480), 
	.A3(U_dsdc_n1579), 
	.A2(U_dsdc_n1481), 
	.A1(FE_PHN771_U_dsdc_n1540));
   OAI22_X2 U_dsdc_U1488 (.ZN(U_dsdc_N4228), 
	.B2(FE_PHN931_U_dsdc_n2094), 
	.B1(U_dsdc_n2057), 
	.A2(U_dsdc_n1482), 
	.A1(U_dsdc_t_xp_cnt_0_));
   NAND3_X2 U_dsdc_U1487 (.ZN(U_dsdc_n1518), 
	.A3(U_dsdc_n1501), 
	.A2(U_dsdc_n1502), 
	.A1(U_dsdc_n1503));
   AOI211_X2 U_dsdc_U1486 (.ZN(U_dsdc_n1520), 
	.C2(U_dsdc_n2063), 
	.C1(U_dsdc_n2064), 
	.B(U_dsdc_n1518), 
	.A(U_dsdc_n1519));
   OAI21_X2 U_dsdc_U1485 (.ZN(U_dsdc_n1542), 
	.B2(U_dsdc_n1521), 
	.B1(U_dsdc_n1522), 
	.A(U_dsdc_n1520));
   NOR3_X2 U_dsdc_U1484 (.ZN(U_dsdc_n1530), 
	.A3(U_dsdc_n1542), 
	.A2(U_dsdc_n1523), 
	.A1(U_dsdc_n1524));
   NOR2_X2 U_dsdc_U1483 (.ZN(U_dsdc_n2061), 
	.A2(U_dsdc_n1675), 
	.A1(U_dsdc_n2065));
   OAI21_X2 U_dsdc_U1482 (.ZN(U_dsdc_n1618), 
	.B2(U_dsdc_n1505), 
	.B1(FE_PHN791_U_dsdc_n1491), 
	.A(U_dsdc_n2058));
   AOI211_X2 U_dsdc_U1481 (.ZN(U_dsdc_n1507), 
	.C2(U_dsdc_n1519), 
	.C1(U_dsdc_n1430), 
	.B(U_dsdc_n1493), 
	.A(ctl_init_done));
   NOR4_X2 U_dsdc_U1480 (.ZN(U_dsdc_n1528), 
	.A4(U_dsdc_n1527), 
	.A3(U_dsdc_n1618), 
	.A2(U_dsdc_n2061), 
	.A1(U_dsdc_n1581));
   OAI211_X2 U_dsdc_U1479 (.ZN(U_dsdc_n2096), 
	.C2(U_dsdc_n343), 
	.C1(U_dsdc_n1530), 
	.B(U_dsdc_n1528), 
	.A(U_dsdc_n1529));
   OAI21_X2 U_dsdc_U1478 (.ZN(U_dsdc_n1588), 
	.B2(U_dsdc_n1575), 
	.B1(U_dsdc_n2064), 
	.A(U_dsdc_n2063));
   NOR2_X2 U_dsdc_U1477 (.ZN(U_dsdc_n1667), 
	.A2(U_dsdc_n1509), 
	.A1(U_dsdc_n1510));
   NOR3_X2 U_dsdc_U1476 (.ZN(U_dsdc_n1580), 
	.A3(U_dsdc_n2063), 
	.A2(U_dsdc_n2051), 
	.A1(U_dsdc_n1564));
   INV_X4 U_dsdc_U1475 (.ZN(U_dsdc_n573), 
	.A(U_dsdc_n1576));
   NAND2_X2 U_dsdc_U1474 (.ZN(U_dsdc_n1578), 
	.A2(U_dsdc_n1728), 
	.A1(U_dsdc_n1536));
   OAI22_X2 U_dsdc_U1472 (.ZN(U_dsdc_rcar_cnt1_nxt[0]), 
	.B2(FE_PHN1052_U_cr_n127), 
	.B1(U_dsdc_n1590), 
	.A2(U_dsdc_n1588), 
	.A1(U_dsdc_rcar_cnt1_0_));
   OAI22_X2 U_dsdc_U1471 (.ZN(U_dsdc_N4229), 
	.B2(U_dsdc_n239), 
	.B1(U_dsdc_n474), 
	.A2(FE_PHN931_U_dsdc_n2094), 
	.A1(U_dsdc_n2057));
   NAND3_X2 U_dsdc_U1470 (.ZN(U_dsdc_n1497), 
	.A3(U_dsdc_n1434), 
	.A2(U_dsdc_n1430), 
	.A1(U_dsdc_n645));
   AOI21_X2 U_dsdc_U1469 (.ZN(U_dsdc_n1676), 
	.B2(cr_do_initialize), 
	.B1(U_dsdc_n1499), 
	.A(U_dsdc_n1498));
   AOI21_X2 U_dsdc_U1468 (.ZN(U_dsdc_n1544), 
	.B2(U_dsdc_n2056), 
	.B1(U_dsdc_n1534), 
	.A(U_dsdc_n1527));
   AOI211_X2 U_dsdc_U1467 (.ZN(U_dsdc_n1514), 
	.C2(U_dsdc_n1435), 
	.C1(U_dsdc_n1512), 
	.B(U_dsdc_n1667), 
	.A(U_dsdc_n1511));
   NOR2_X2 U_dsdc_U1466 (.ZN(U_dsdc_n1429), 
	.A2(cr_do_self_ref_rp), 
	.A1(U_dsdc_n2052));
   NAND3_X2 U_dsdc_U1465 (.ZN(U_dsdc_n1513), 
	.A3(U_cr_n61), 
	.A2(cr_exn_mode_reg_update), 
	.A1(U_dsdc_n1429));
   NAND4_X2 U_dsdc_U1464 (.ZN(U_dsdc_n1515), 
	.A4(U_dsdc_n1513), 
	.A3(U_dsdc_n1579), 
	.A2(U_dsdc_n1514), 
	.A1(U_dsdc_n1544));
   AOI221_X2 U_dsdc_U1463 (.ZN(U_dsdc_n1517), 
	.C2(U_dsdc_operation_cs_0_), 
	.C1(U_dsdc_n1516), 
	.B2(U_dsdc_operation_cs_0_), 
	.B1(U_dsdc_n1518), 
	.A(U_dsdc_n1515));
   NAND4_X2 U_dsdc_U1462 (.ZN(U_dsdc_n2097), 
	.A4(U_dsdc_n1517), 
	.A3(U_dsdc_n1676), 
	.A2(U_dsdc_n1733), 
	.A1(FE_PHN771_U_dsdc_n1540));
   AOI21_X2 U_dsdc_U1461 (.ZN(U_dsdc_n1582), 
	.B2(U_dsdc_rcar_cnt1_1_), 
	.B1(U_dsdc_rcar_cnt1_0_), 
	.A(U_dsdc_n1583));
   NOR2_X2 U_dsdc_U1459 (.ZN(U_dsdc_n1328), 
	.A2(U_dsdc_n1325), 
	.A1(U_dsdc_n1326));
   AOI21_X2 U_dsdc_U1458 (.ZN(U_dsdc_n1333), 
	.B2(cr_t_rp[0]), 
	.B1(U_dsdc_n1327), 
	.A(U_dsdc_n1336));
   NOR2_X2 U_dsdc_U1457 (.ZN(U_dsdc_n1334), 
	.A2(cr_t_rp[0]), 
	.A1(U_dsdc_n1328));
   NOR2_X2 U_dsdc_U1456 (.ZN(U_dsdc_n1331), 
	.A2(cr_t_rp[1]), 
	.A1(FE_PHN3514_U_cr_n148));
   NOR2_X2 U_dsdc_U1455 (.ZN(U_dsdc_n1421), 
	.A2(U_dsdc_n1425), 
	.A1(U_dsdc_n1357));
   AOI21_X2 U_dsdc_U1454 (.ZN(U_dsdc_n1335), 
	.B2(U_dsdc_n1629), 
	.B1(U_dsdc_n1421), 
	.A(U_dsdc_n1426));
   AOI22_X2 U_dsdc_U1453 (.ZN(U_dsdc_n1332), 
	.B2(U_dsdc_n1330), 
	.B1(U_dsdc_n1335), 
	.A2(U_dsdc_n1331), 
	.A1(U_dsdc_n1334));
   OAI21_X2 U_dsdc_U1452 (.ZN(U_dsdc_rp_cnt2_nxt[1]), 
	.B2(FE_PHN3012_U_cr_n147), 
	.B1(U_dsdc_n1333), 
	.A(U_dsdc_n1332));
   INV_X4 U_dsdc_U1451 (.ZN(U_dsdc_n1397), 
	.A(U_dsdc_n1349));
   NAND2_X2 U_dsdc_U1450 (.ZN(U_dsdc_n1805), 
	.A2(U_dsdc_n1414), 
	.A1(FE_PHN671_U_dsdc_n1637));
   NAND2_X2 U_dsdc_U1449 (.ZN(U_dsdc_n1803), 
	.A2(U_dsdc_n652), 
	.A1(U_dsdc_n915));
   NAND2_X2 U_dsdc_U1448 (.ZN(U_dsdc_n2074), 
	.A2(U_dsdc_n1803), 
	.A1(U_dsdc_n1804));
   NOR2_X2 U_dsdc_U1447 (.ZN(U_dsdc_n1398), 
	.A2(U_dsdc_n360), 
	.A1(U_dsdc_n2074));
   AOI21_X2 U_dsdc_U1446 (.ZN(U_dsdc_n730), 
	.B2(U_dsdc_n736), 
	.B1(U_dsdc_n740), 
	.A(U_dsdc_n728));
   OAI21_X2 U_dsdc_U1445 (.ZN(U_dsdc_n731), 
	.B2(U_dsdc_n440), 
	.B1(U_dsdc_n730), 
	.A(U_dsdc_n729));
   AOI21_X2 U_dsdc_U1444 (.ZN(U_dsdc_n732), 
	.B2(U_dsdc_n1415), 
	.B1(U_dsdc_n1805), 
	.A(U_dsdc_n731));
   OAI211_X2 U_dsdc_U1443 (.ZN(U_dsdc_n734), 
	.C2(U_dsdc_n733), 
	.C1(U_dsdc_n1397), 
	.B(U_dsdc_n732), 
	.A(U_dsdc_n1398));
   NOR2_X2 U_dsdc_U1442 (.ZN(U_dsdc_n329), 
	.A2(U_dsdc_n734), 
	.A1(hiu_terminate));
   NAND2_X2 U_dsdc_U1440 (.ZN(U_dsdc_n1812), 
	.A2(FE_PHN1416_U_dsdc_r_col_addr_1_), 
	.A1(U_dsdc_n619));
   NAND3_X2 U_dsdc_U1439 (.ZN(U_dsdc_n1670), 
	.A3(U_dsdc_n1497), 
	.A2(U_dsdc_n646), 
	.A1(U_dsdc_n1480));
   AOI21_X2 U_dsdc_U1433 (.ZN(U_dsdc_n1307), 
	.B2(U_dsdc_n1294), 
	.B1(U_dsdc_n1295), 
	.A(U_dsdc_n1293));
   AOI21_X2 U_dsdc_U1432 (.ZN(U_dsdc_n1303), 
	.B2(U_dsdc_n1297), 
	.B1(U_dsdc_wr_cnt_2_), 
	.A(U_dsdc_n1296));
   AOI21_X2 U_dsdc_U1431 (.ZN(U_dsdc_n1301), 
	.B2(U_dsdc_n1299), 
	.B1(U_dsdc_n1300), 
	.A(U_dsdc_n1298));
   NOR2_X2 U_dsdc_U1430 (.ZN(U_dsdc_n1304), 
	.A2(U_dsdc_n1309), 
	.A1(U_dsdc_n1301));
   NAND3_X2 U_dsdc_U1429 (.ZN(U_dsdc_n1302), 
	.A3(cr_t_wr[1]), 
	.A2(cr_t_wr[0]), 
	.A1(U_dsdc_n1304));
   OAI21_X2 U_dsdc_U1428 (.ZN(U_dsdc_wr_cnt_nxt[2]), 
	.B2(U_dsdc_n1303), 
	.B1(U_dsdc_n1307), 
	.A(U_dsdc_n1302));
   OAI21_X2 U_dsdc_U1406 (.ZN(U_dsdc_n1338), 
	.B2(cr_t_rp[2]), 
	.B1(cr_t_rp[1]), 
	.A(U_dsdc_n1334));
   AOI22_X2 U_dsdc_U1405 (.ZN(U_dsdc_n1337), 
	.B2(U_dsdc_n171), 
	.B1(U_dsdc_n1335), 
	.A2(cr_t_rp[0]), 
	.A1(U_dsdc_n1336));
   NAND2_X2 U_dsdc_U1404 (.ZN(U_dsdc_rp_cnt2_nxt[0]), 
	.A2(U_dsdc_n1337), 
	.A1(U_dsdc_n1338));
   NAND2_X2 U_dsdc_U1400 (.ZN(U_dsdc_n1123), 
	.A2(U_dsdc_oldest_bank_0_), 
	.A1(U_dsdc_n1003));
   INV_X4 U_dsdc_U1398 (.ZN(U_dsdc_n1308), 
	.A(U_dsdc_n1304));
   OAI22_X2 U_dsdc_U1397 (.ZN(U_dsdc_wr_cnt_nxt[1]), 
	.B2(U_dsdc_n1305), 
	.B1(U_dsdc_n1307), 
	.A2(U_dsdc_n1306), 
	.A1(U_dsdc_n1308));
   OAI22_X2 U_dsdc_U1396 (.ZN(U_dsdc_wr_cnt_nxt[0]), 
	.B2(U_dsdc_n1307), 
	.B1(U_dsdc_wr_cnt_0_), 
	.A2(cr_t_wr[0]), 
	.A1(U_dsdc_n1308));
   AOI221_X2 U_dsdc_U1395 (.ZN(U_dsdc_n1778), 
	.C2(U_dsdc_n1791), 
	.C1(U_dsdc_row_cnt_1_), 
	.B2(U_dsdc_n1791), 
	.B1(U_dsdc_row_cnt_0_), 
	.A(U_dsdc_n1800));
   NAND2_X2 U_dsdc_U1394 (.ZN(U_dsdc_n1774), 
	.A2(U_dsdc_n577), 
	.A1(U_dsdc_n1778));
   NOR4_X2 U_dsdc_U1393 (.ZN(U_dsdc_N4241), 
	.A4(U_cr_n42), 
	.A3(FE_PHN1064_cr_row_addr_width_3_), 
	.A2(cr_row_addr_width[0]), 
	.A1(FE_PHN3054_cr_row_addr_width_2_));
   NOR4_X2 U_dsdc_U1392 (.ZN(U_dsdc_N4240), 
	.A4(U_cr_n21), 
	.A3(FE_PHN1064_cr_row_addr_width_3_), 
	.A2(FE_PHN3054_cr_row_addr_width_2_), 
	.A1(cr_row_addr_width[1]));
   INV_X4 U_dsdc_U1391 (.ZN(U_dsdc_n1757), 
	.A(U_dsdc_n1578));
   AOI22_X2 U_dsdc_U1390 (.ZN(U_dsdc_n1801), 
	.B2(cr_ref_all_after_sr), 
	.B1(U_dsdc_n1757), 
	.A2(cr_ref_all_before_sr), 
	.A1(U_dsdc_n1758));
   INV_X4 U_dsdc_U1389 (.ZN(U_dsdc_n1797), 
	.A(U_dsdc_n1801));
   AOI22_X2 U_dsdc_U1388 (.ZN(U_dsdc_n1775), 
	.B2(U_dsdc_n1797), 
	.B1(U_dsdc_num_row[3]), 
	.A2(U_dsdc_row_cnt_3_), 
	.A1(U_dsdc_n1774));
   NAND2_X2 U_dsdc_U1387 (.ZN(U_dsdc_n582), 
	.A2(U_dsdc_n574), 
	.A1(U_dsdc_n1791));
   NAND2_X2 U_dsdc_U1386 (.ZN(U_dsdc_n375), 
	.A2(U_dsdc_n582), 
	.A1(U_dsdc_n1775));
   NAND2_X2 U_dsdc_U1385 (.ZN(U_dsdc_write_start_nxt), 
	.A2(U_dsdc_n1314), 
	.A1(U_dsdc_n1052));
   AOI21_X2 U_dsdc_U1383 (.ZN(U_dsdc_n1872), 
	.B2(U_dsdc_n1633), 
	.B1(U_dsdc_n1629), 
	.A(U_dsdc_n1632));
   OAI22_X2 U_dsdc_U1382 (.ZN(U_dsdc_n2070), 
	.B2(U_dsdc_n1629), 
	.B1(U_dsdc_n1423), 
	.A2(U_dsdc_n1633), 
	.A1(U_dsdc_n1424));
   NAND2_X2 U_dsdc_U1381 (.ZN(U_dsdc_n705), 
	.A2(U_dsdc_n2070), 
	.A1(U_dsdc_n1632));
   AOI21_X2 U_dsdc_U1379 (.ZN(U_dsdc_n1285), 
	.B2(U_dsdc_n1284), 
	.B1(hiu_wrapped_burst), 
	.A(U_dsdc_n1438));
   AOI211_X2 U_dsdc_U1378 (.ZN(U_dsdc_n1291), 
	.C2(U_dsdc_n1383), 
	.C1(U_dsdc_access_cs_4_), 
	.B(U_dsdc_n1287), 
	.A(U_dsdc_n1288));
   NAND3_X2 U_dsdc_U1377 (.ZN(U_dsdc_n[2088]), 
	.A3(U_dsdc_n1289), 
	.A2(U_dsdc_n1290), 
	.A1(U_dsdc_n1291));
   NAND2_X2 U_dsdc_U1376 (.ZN(U_dsdc_n1390), 
	.A2(U_dsdc_oldest_bank_1_), 
	.A1(U_dsdc_n1003));
   OAI21_X2 U_dsdc_U1375 (.ZN(U_dsdc_close_bank_addr_1_), 
	.B2(U_dsdc_n1130), 
	.B1(U_dsdc_n1391), 
	.A(U_dsdc_n1390));
   NAND2_X2 U_dsdc_U1372 (.ZN(U_dsdc_n766), 
	.A2(U_cr_n58), 
	.A1(U_dsdc_n1152));
   NAND2_X2 U_dsdc_U1371 (.ZN(U_dsdc_n1359), 
	.A2(U_dsdc_n766), 
	.A1(U_dsdc_n1344));
   NOR4_X2 U_dsdc_U1370 (.ZN(U_dsdc_n1369), 
	.A4(U_dsdc_n1363), 
	.A3(U_dsdc_n1364), 
	.A2(U_dsdc_n1365), 
	.A1(U_dsdc_n1366));
   NAND2_X2 U_dsdc_U1369 (.ZN(U_dsdc_n1368), 
	.A2(U_dsdc_n766), 
	.A1(U_dsdc_n767));
   NAND2_X2 U_dsdc_U1368 (.ZN(U_dsdc_n1387), 
	.A2(U_dsdc_n1367), 
	.A1(U_dsdc_n1805));
   NAND4_X2 U_dsdc_U1367 (.ZN(U_dsdc_n1371), 
	.A4(U_dsdc_n1387), 
	.A3(U_dsdc_n1368), 
	.A2(U_dsdc_n1369), 
	.A1(U_dsdc_n1370));
   AOI21_X2 U_dsdc_U1366 (.ZN(U_dsdc_n1377), 
	.B2(U_dsdc_n1372), 
	.B1(U_dsdc_n1373), 
	.A(U_dsdc_n1371));
   NAND2_X2 U_dsdc_U1365 (.ZN(U_dsdc_n1375), 
	.A2(U_dsdc_n983), 
	.A1(U_dsdc_n899));
   NAND3_X2 U_dsdc_U1364 (.ZN(U_dsdc_n[2092]), 
	.A3(U_dsdc_n1375), 
	.A2(U_dsdc_n1376), 
	.A1(U_dsdc_n1377));
   OAI22_X2 U_dsdc_U1363 (.ZN(U_dsdc_bm_close_bank_1_), 
	.B2(U_dsdc_n1123), 
	.B1(U_dsdc_oldest_bank_1_), 
	.A2(U_dsdc_n600), 
	.A1(U_dsdc_n1391));
   OAI21_X2 U_dsdc_U1362 (.ZN(U_dsdc_n1178), 
	.B2(U_dsdc_n1174), 
	.B1(U_dsdc_bm_rc_cnt_0__3_), 
	.A(n83));
   AOI21_X2 U_dsdc_U1361 (.ZN(U_dsdc_n1177), 
	.B2(U_dsdc_bm_rc_cnt_0__1_), 
	.B1(U_dsdc_bm_rc_cnt_0__0_), 
	.A(U_dsdc_n1176));
   OAI22_X2 U_dsdc_U1359 (.ZN(U_dsdc_N4333), 
	.B2(U_cr_n106), 
	.B1(n83), 
	.A2(FE_PHN3247_U_dsdc_n1177), 
	.A1(U_dsdc_n1178));
   OAI22_X2 U_dsdc_U1357 (.ZN(U_dsdc_N4332), 
	.B2(n83), 
	.B1(FE_OFN23_U_cr_n64), 
	.A2(U_dsdc_bm_rc_cnt_0__0_), 
	.A1(U_dsdc_n1178));
   OAI22_X2 U_dsdc_U1356 (.ZN(U_dsdc_n300), 
	.B2(U_dsdc_n1089), 
	.B1(U_dsdc_n1393), 
	.A2(FE_PHN2036_U_dsdc_cas_latency_cnt_0_), 
	.A1(U_dsdc_n1090));
   AOI21_X2 U_dsdc_U1355 (.ZN(U_dsdc_n1251), 
	.B2(U_dsdc_n1037), 
	.B1(U_dsdc_n1038), 
	.A(U_dsdc_n1293));
   AOI21_X2 U_dsdc_U1351 (.ZN(U_dsdc_n1851), 
	.B2(U_dsdc_n1847), 
	.B1(U_dsdc_n1867), 
	.A(U_dsdc_n1961));
   OAI221_X2 U_dsdc_U1350 (.ZN(U_dsdc_n1853), 
	.C2(U_dsdc_n1859), 
	.C1(FE_PHN958_U_dsdc_n353), 
	.B2(U_dsdc_n1860), 
	.B1(U_dsdc_bm_bank_age_2__0_), 
	.A(U_dsdc_n1851));
   OAI21_X2 U_dsdc_U1349 (.ZN(U_dsdc_n1854), 
	.B2(U_dsdc_n1853), 
	.B1(U_dsdc_n178), 
	.A(U_dsdc_n1852));
   OAI21_X2 U_dsdc_U1348 (.ZN(U_dsdc_n210), 
	.B2(U_dsdc_n1856), 
	.B1(U_dsdc_n1859), 
	.A(U_dsdc_n1854));
   OAI21_X2 U_dsdc_U1347 (.ZN(U_dsdc_bm_close_bank_0_), 
	.B2(U_dsdc_n572), 
	.B1(U_dsdc_n1391), 
	.A(U_dsdc_n1001));
   OAI21_X2 U_dsdc_U1346 (.ZN(U_dsdc_n1233), 
	.B2(U_dsdc_n1227), 
	.B1(U_dsdc_bm_rc_cnt_3__3_), 
	.A(U_dsdc_n313));
   AOI21_X2 U_dsdc_U1345 (.ZN(U_dsdc_n1231), 
	.B2(U_dsdc_bm_rc_cnt_3__1_), 
	.B1(U_dsdc_bm_rc_cnt_3__0_), 
	.A(U_dsdc_n1229));
   OAI22_X2 U_dsdc_U1344 (.ZN(U_dsdc_N4474), 
	.B2(U_cr_n106), 
	.B1(U_dsdc_n313), 
	.A2(FE_PHN3371_U_dsdc_n1231), 
	.A1(U_dsdc_n1233));
   OAI22_X2 U_dsdc_U1343 (.ZN(U_dsdc_N4473), 
	.B2(U_dsdc_n313), 
	.B1(FE_OFN23_U_cr_n64), 
	.A2(U_dsdc_bm_rc_cnt_3__0_), 
	.A1(U_dsdc_n1233));
   INV_X4 U_dsdc_U1342 (.ZN(U_dsdc_n289), 
	.A(U_dsdc_n763));
   AOI21_X2 U_dsdc_U1341 (.ZN(U_dsdc_n1785), 
	.B2(U_dsdc_n1788), 
	.B1(U_dsdc_n1791), 
	.A(U_dsdc_n1800));
   NAND2_X2 U_dsdc_U1340 (.ZN(U_dsdc_n1781), 
	.A2(U_dsdc_n578), 
	.A1(U_dsdc_n1785));
   NAND2_X2 U_dsdc_U1339 (.ZN(U_dsdc_n1662), 
	.A2(cr_row_addr_width[0]), 
	.A1(cr_row_addr_width[1]));
   NAND2_X2 U_dsdc_U1338 (.ZN(U_dsdc_n1653), 
	.A2(FE_PHN3054_cr_row_addr_width_2_), 
	.A1(U_dsdc_n1652));
   NAND2_X2 U_dsdc_U1336 (.ZN(U_dsdc_n1656), 
	.A2(U_cr_n70), 
	.A1(U_dsdc_n1653));
   NAND2_X2 U_dsdc_U1335 (.ZN(U_dsdc_n1661), 
	.A2(U_dsdc_n1656), 
	.A1(U_dsdc_n1657));
   NOR2_X2 U_dsdc_U1334 (.ZN(U_dsdc_N4253), 
	.A2(U_dsdc_n1661), 
	.A1(U_dsdc_n1658));
   NOR2_X2 U_dsdc_U1333 (.ZN(U_dsdc_N4252), 
	.A2(U_dsdc_n1661), 
	.A1(U_dsdc_n1659));
   NOR2_X2 U_dsdc_U1332 (.ZN(U_dsdc_N4250), 
	.A2(U_dsdc_n1661), 
	.A1(U_dsdc_n1662));
   NOR4_X2 U_dsdc_U1331 (.ZN(U_dsdc_N4248), 
	.A4(U_cr_n70), 
	.A3(U_cr_n21), 
	.A2(FE_PHN3054_cr_row_addr_width_2_), 
	.A1(cr_row_addr_width[1]));
   NOR2_X2 U_dsdc_U1330 (.ZN(U_dsdc_N4246), 
	.A2(U_dsdc_n1653), 
	.A1(FE_PHN1064_cr_row_addr_width_3_));
   NAND2_X2 U_dsdc_U1329 (.ZN(U_dsdc_n1655), 
	.A2(U_dsdc_n1654), 
	.A1(U_dsdc_n1657));
   NOR2_X2 U_dsdc_U1328 (.ZN(U_dsdc_N4244), 
	.A2(U_dsdc_n1655), 
	.A1(U_dsdc_n1659));
   NOR2_X2 U_dsdc_U1327 (.ZN(U_dsdc_N4242), 
	.A2(U_dsdc_n1656), 
	.A1(U_dsdc_n1662));
   NOR2_X2 U_dsdc_U1326 (.ZN(U_dsdc_n614), 
	.A2(U_dsdc_n613), 
	.A1(U_dsdc_N4242));
   NAND2_X2 U_dsdc_U1325 (.ZN(U_dsdc_n1660), 
	.A2(U_cr_n21), 
	.A1(U_cr_n42));
   NAND2_X2 U_dsdc_U1324 (.ZN(U_dsdc_n615), 
	.A2(U_dsdc_n345), 
	.A1(U_dsdc_n614));
   NOR2_X2 U_dsdc_U1323 (.ZN(U_dsdc_n616), 
	.A2(U_dsdc_n615), 
	.A1(U_dsdc_N4244));
   NAND2_X2 U_dsdc_U1322 (.ZN(U_dsdc_n617), 
	.A2(U_dsdc_n346), 
	.A1(U_dsdc_n616));
   NOR2_X2 U_dsdc_U1321 (.ZN(U_dsdc_n618), 
	.A2(U_dsdc_n617), 
	.A1(U_dsdc_N4246));
   NAND2_X2 U_dsdc_U1320 (.ZN(U_dsdc_n606), 
	.A2(U_dsdc_n358), 
	.A1(U_dsdc_n618));
   NOR2_X2 U_dsdc_U1319 (.ZN(U_dsdc_n607), 
	.A2(U_dsdc_n606), 
	.A1(U_dsdc_N4248));
   NAND2_X2 U_dsdc_U1318 (.ZN(U_dsdc_n608), 
	.A2(U_dsdc_n357), 
	.A1(U_dsdc_n607));
   NOR2_X2 U_dsdc_U1317 (.ZN(U_dsdc_n609), 
	.A2(U_dsdc_n608), 
	.A1(U_dsdc_N4250));
   NAND2_X2 U_dsdc_U1316 (.ZN(U_dsdc_n610), 
	.A2(U_dsdc_n399), 
	.A1(U_dsdc_n609));
   NOR2_X2 U_dsdc_U1315 (.ZN(U_dsdc_n611), 
	.A2(U_dsdc_n610), 
	.A1(U_dsdc_N4252));
   AOI22_X2 U_dsdc_U1314 (.ZN(U_dsdc_n1782), 
	.B2(U_dsdc_n1797), 
	.B1(U_dsdc_num_row[15]), 
	.A2(U_dsdc_n1781), 
	.A1(U_dsdc_row_cnt_15_));
   NOR3_X2 U_dsdc_U1313 (.ZN(U_dsdc_n1862), 
	.A3(U_dsdc_n1856), 
	.A2(U_dsdc_n1859), 
	.A1(U_dsdc_bm_bank_age_2__2_));
   OAI21_X2 U_dsdc_U1312 (.ZN(U_dsdc_n1863), 
	.B2(U_dsdc_n1862), 
	.B1(U_dsdc_n1868), 
	.A(U_dsdc_n459));
   OAI21_X2 U_dsdc_U1311 (.ZN(U_dsdc_n212), 
	.B2(U_dsdc_n459), 
	.B1(U_dsdc_n1864), 
	.A(U_dsdc_n1863));
   AOI21_X2 U_dsdc_U1310 (.ZN(U_dsdc_n1891), 
	.B2(U_dsdc_n1888), 
	.B1(U_dsdc_n1907), 
	.A(U_dsdc_n1961));
   OAI221_X2 U_dsdc_U1309 (.ZN(U_dsdc_n1893), 
	.C2(U_dsdc_n1899), 
	.C1(U_dsdc_n304), 
	.B2(U_dsdc_n1900), 
	.B1(U_dsdc_bm_bank_age_3__0_), 
	.A(U_dsdc_n1891));
   OAI21_X2 U_dsdc_U1308 (.ZN(U_dsdc_n1894), 
	.B2(U_dsdc_n1893), 
	.B1(U_dsdc_n302), 
	.A(U_dsdc_n1892));
   OAI21_X2 U_dsdc_U1307 (.ZN(U_dsdc_n219), 
	.B2(U_dsdc_n1896), 
	.B1(U_dsdc_n1899), 
	.A(U_dsdc_n1894));
   AOI21_X2 U_dsdc_U1306 (.ZN(U_dsdc_n1921), 
	.B2(U_dsdc_n1918), 
	.B1(U_dsdc_n1937), 
	.A(U_dsdc_n1961));
   OAI221_X2 U_dsdc_U1305 (.ZN(U_dsdc_n1923), 
	.C2(U_dsdc_n1929), 
	.C1(FE_PHN897_U_dsdc_n352), 
	.B2(U_dsdc_n1930), 
	.B1(U_dsdc_bm_bank_age_1__0_), 
	.A(U_dsdc_n1921));
   OAI21_X2 U_dsdc_U1304 (.ZN(U_dsdc_n1924), 
	.B2(U_dsdc_n1923), 
	.B1(U_dsdc_n335), 
	.A(U_dsdc_n1922));
   OAI21_X2 U_dsdc_U1303 (.ZN(U_dsdc_n224), 
	.B2(U_dsdc_n1926), 
	.B1(U_dsdc_n1929), 
	.A(FE_PHN3467_U_dsdc_n1924));
   NOR2_X2 U_dsdc_U1302 (.ZN(U_dsdc_n704), 
	.A2(U_dsdc_n2071), 
	.A1(U_dsdc_n994));
   NOR2_X2 U_dsdc_U1301 (.ZN(U_dsdc_n901), 
	.A2(U_dsdc_n704), 
	.A1(U_dsdc_n1367));
   NOR3_X2 U_dsdc_U1300 (.ZN(U_dsdc_n1932), 
	.A3(U_dsdc_n1926), 
	.A2(U_dsdc_n1929), 
	.A1(U_dsdc_bm_bank_age_1__2_));
   OAI21_X2 U_dsdc_U1299 (.ZN(U_dsdc_n1933), 
	.B2(U_dsdc_n1932), 
	.B1(U_dsdc_n1938), 
	.A(FE_PHN3077_U_dsdc_n460));
   OAI21_X2 U_dsdc_U1298 (.ZN(U_dsdc_n226), 
	.B2(FE_PHN3077_U_dsdc_n460), 
	.B1(U_dsdc_n1934), 
	.A(U_dsdc_n1933));
   OAI21_X2 U_dsdc_U1297 (.ZN(U_dsdc_n1206), 
	.B2(U_dsdc_n1202), 
	.B1(U_dsdc_bm_rc_cnt_2__3_), 
	.A(U_dsdc_n310));
   OAI22_X2 U_dsdc_U1296 (.ZN(U_dsdc_N4426), 
	.B2(U_dsdc_n310), 
	.B1(FE_OFN23_U_cr_n64), 
	.A2(FE_PHN3509_U_dsdc_bm_rc_cnt_2__0_), 
	.A1(U_dsdc_n1206));
   OAI21_X2 U_dsdc_U1295 (.ZN(U_dsdc_n1192), 
	.B2(U_dsdc_n1188), 
	.B1(U_dsdc_bm_rc_cnt_1__3_), 
	.A(U_dsdc_n620));
   AOI21_X2 U_dsdc_U1294 (.ZN(U_dsdc_n1191), 
	.B2(U_dsdc_bm_rc_cnt_1__1_), 
	.B1(FE_PHN3508_U_dsdc_bm_rc_cnt_1__0_), 
	.A(U_dsdc_n1190));
   OAI22_X2 U_dsdc_U1293 (.ZN(U_dsdc_N4380), 
	.B2(U_cr_n106), 
	.B1(U_dsdc_n620), 
	.A2(FE_PHN3252_U_dsdc_n1191), 
	.A1(U_dsdc_n1192));
   AOI21_X2 U_dsdc_U1292 (.ZN(U_dsdc_n1205), 
	.B2(U_dsdc_bm_rc_cnt_2__1_), 
	.B1(FE_PHN3509_U_dsdc_bm_rc_cnt_2__0_), 
	.A(U_dsdc_n1204));
   OAI22_X2 U_dsdc_U1291 (.ZN(U_dsdc_N4427), 
	.B2(U_cr_n106), 
	.B1(U_dsdc_n310), 
	.A2(FE_PHN3259_U_dsdc_n1205), 
	.A1(U_dsdc_n1206));
   OAI22_X2 U_dsdc_U1290 (.ZN(U_dsdc_N4379), 
	.B2(U_dsdc_n620), 
	.B1(FE_OFN23_U_cr_n64), 
	.A2(FE_PHN3508_U_dsdc_bm_rc_cnt_1__0_), 
	.A1(U_dsdc_n1192));
   OAI22_X2 U_dsdc_U1286 (.ZN(U_dsdc_wtr_cnt_nxt[0]), 
	.B2(U_dsdc_n1251), 
	.B1(U_dsdc_wtr_cnt_0_), 
	.A2(cr_t_wtr[0]), 
	.A1(U_dsdc_n1252));
   NAND2_X2 U_dsdc_U1285 (.ZN(U_dsdc_n1185), 
	.A2(U_dsdc_n1181), 
	.A1(n83));
   AOI21_X2 U_dsdc_U1284 (.ZN(U_dsdc_n1184), 
	.B2(U_dsdc_bm_ras_cnt_0__1_), 
	.B1(FE_PHN3511_U_dsdc_bm_ras_cnt_0__0_), 
	.A(U_dsdc_n1183));
   OAI22_X2 U_dsdc_U1282 (.ZN(U_dsdc_N4320), 
	.B2(U_cr_n120), 
	.B1(n83), 
	.A2(FE_PHN3258_U_dsdc_n1184), 
	.A1(U_dsdc_n1185));
   OAI22_X2 U_dsdc_U1280 (.ZN(U_dsdc_N4319), 
	.B2(n95), 
	.B1(n83), 
	.A2(FE_PHN3511_U_dsdc_bm_ras_cnt_0__0_), 
	.A1(U_dsdc_n1185));
   OAI22_X2 U_dsdc_U1279 (.ZN(U_dsdc_wtr_cnt_nxt[1]), 
	.B2(U_dsdc_n1246), 
	.B1(U_dsdc_n1251), 
	.A2(U_dsdc_n1247), 
	.A1(U_dsdc_n1252));
   NAND2_X2 U_dsdc_U1278 (.ZN(U_dsdc_n1250), 
	.A2(cr_t_wtr[0]), 
	.A1(cr_t_wtr[1]));
   AOI21_X2 U_dsdc_U1277 (.ZN(U_dsdc_n1249), 
	.B2(U_dsdc_n1248), 
	.B1(U_dsdc_wtr_cnt_2_), 
	.A(U_dsdc_n1284));
   OAI22_X2 U_dsdc_U1276 (.ZN(U_dsdc_wtr_cnt_nxt[2]), 
	.B2(U_dsdc_n1249), 
	.B1(U_dsdc_n1251), 
	.A2(U_dsdc_n1250), 
	.A1(U_dsdc_n1252));
   NAND2_X2 U_dsdc_U1275 (.ZN(U_dsdc_n1243), 
	.A2(U_dsdc_n1237), 
	.A1(U_dsdc_n313));
   AOI21_X2 U_dsdc_U1274 (.ZN(U_dsdc_n1241), 
	.B2(U_dsdc_bm_ras_cnt_3__1_), 
	.B1(FE_PHN3513_U_dsdc_bm_ras_cnt_3__0_), 
	.A(U_dsdc_n1239));
   AOI22_X2 U_dsdc_U1273 (.ZN(U_dsdc_n1777), 
	.B2(U_dsdc_n204), 
	.B1(U_dsdc_n325), 
	.A2(U_dsdc_n1797), 
	.A1(U_dsdc_num_row[2]));
   OAI21_X2 U_dsdc_U1272 (.ZN(U_dsdc_n374), 
	.B2(U_dsdc_n204), 
	.B1(U_dsdc_n1778), 
	.A(U_dsdc_n1777));
   NOR3_X2 U_dsdc_U1271 (.ZN(U_dsdc_n1972), 
	.A3(U_dsdc_n384), 
	.A2(U_dsdc_n1941), 
	.A1(U_dsdc_r_bm_open_bank[0]));
   NOR3_X2 U_dsdc_U1270 (.ZN(U_dsdc_n2081), 
	.A3(U_dsdc_n1942), 
	.A2(U_dsdc_n384), 
	.A1(U_dsdc_r_bm_close_bank_0_));
   INV_X4 U_dsdc_U1269 (.ZN(U_dsdc_n1965), 
	.A(U_dsdc_n2081));
   NAND2_X2 U_dsdc_U1268 (.ZN(U_dsdc_n480), 
	.A2(U_dsdc_n478), 
	.A1(U_dsdc_n479));
   NOR2_X2 U_dsdc_U1267 (.ZN(U_dsdc_n1947), 
	.A2(U_dsdc_n480), 
	.A1(U_dsdc_n1945));
   OAI21_X2 U_dsdc_U1263 (.ZN(U_dsdc_n2083), 
	.B2(U_dsdc_n2080), 
	.B1(U_dsdc_n1965), 
	.A(U_dsdc_n1956));
   AOI221_X2 U_dsdc_U1262 (.ZN(U_dsdc_n1958), 
	.C2(FE_PHN3235_U_dsdc_n201), 
	.C1(U_dsdc_n1972), 
	.B2(U_dsdc_bm_bank_age_0__0_), 
	.B1(U_dsdc_n2081), 
	.A(U_dsdc_n2083));
   NAND3_X2 U_dsdc_U1261 (.ZN(U_dsdc_n1962), 
	.A3(U_dsdc_n2080), 
	.A2(FE_PHN3235_U_dsdc_n201), 
	.A1(U_dsdc_n435));
   OAI221_X2 U_dsdc_U1260 (.ZN(U_dsdc_n228), 
	.C2(U_dsdc_n1958), 
	.C1(U_dsdc_n435), 
	.B2(U_dsdc_n1959), 
	.B1(U_dsdc_bm_bank_age_0__1_), 
	.A(U_dsdc_n1957));
   NOR2_X2 U_dsdc_U1259 (.ZN(U_dsdc_n1612), 
	.A2(U_dsdc_n1483), 
	.A1(U_dsdc_n939));
   NAND2_X2 U_dsdc_U1258 (.ZN(U_dsdc_n1601), 
	.A2(U_dsdc_n651), 
	.A1(U_dsdc_n1343));
   NOR3_X2 U_dsdc_U1257 (.ZN(U_dsdc_n1389), 
	.A3(U_dsdc_n1495), 
	.A2(U_dsdc_n1336), 
	.A1(U_dsdc_n1311));
   NOR3_X2 U_dsdc_U1256 (.ZN(U_dsdc_n1417), 
	.A3(U_dsdc_n1592), 
	.A2(U_dsdc_n659), 
	.A1(U_dsdc_n1383));
   NAND2_X2 U_dsdc_U1255 (.ZN(U_dsdc_n1213), 
	.A2(U_dsdc_n1209), 
	.A1(U_dsdc_n310));
   OAI22_X2 U_dsdc_U1254 (.ZN(U_dsdc_N4413), 
	.B2(n95), 
	.B1(U_dsdc_n310), 
	.A2(FE_PHN3510_U_dsdc_bm_ras_cnt_2__0_), 
	.A1(U_dsdc_n1213));
   AOI21_X2 U_dsdc_U1253 (.ZN(U_dsdc_n1212), 
	.B2(U_dsdc_bm_ras_cnt_2__1_), 
	.B1(FE_PHN3510_U_dsdc_bm_ras_cnt_2__0_), 
	.A(U_dsdc_n1211));
   OAI22_X2 U_dsdc_U1252 (.ZN(U_dsdc_N4414), 
	.B2(U_cr_n120), 
	.B1(U_dsdc_n310), 
	.A2(FE_PHN3260_U_dsdc_n1212), 
	.A1(U_dsdc_n1213));
   NAND2_X2 U_dsdc_U1251 (.ZN(U_dsdc_n1199), 
	.A2(U_dsdc_n1195), 
	.A1(U_dsdc_n620));
   OAI22_X2 U_dsdc_U1250 (.ZN(U_dsdc_N4366), 
	.B2(FE_OFN365_n95), 
	.B1(U_dsdc_n620), 
	.A2(FE_PHN3507_U_dsdc_bm_ras_cnt_1__0_), 
	.A1(U_dsdc_n1199));
   AOI21_X2 U_dsdc_U1249 (.ZN(U_dsdc_n1198), 
	.B2(U_dsdc_bm_ras_cnt_1__1_), 
	.B1(FE_PHN3507_U_dsdc_bm_ras_cnt_1__0_), 
	.A(U_dsdc_n1197));
   OAI22_X2 U_dsdc_U1248 (.ZN(U_dsdc_N4367), 
	.B2(U_cr_n120), 
	.B1(U_dsdc_n620), 
	.A2(FE_PHN3256_U_dsdc_n1198), 
	.A1(U_dsdc_n1199));
   NOR3_X2 U_dsdc_U1247 (.ZN(U_dsdc_n1541), 
	.A3(U_dsdc_n2055), 
	.A2(U_dsdc_n1533), 
	.A1(U_dsdc_n1534));
   AOI211_X2 U_dsdc_U1246 (.ZN(U_dsdc_n1539), 
	.C2(U_dsdc_n1621), 
	.C1(U_dsdc_n1431), 
	.B(U_dsdc_n1538), 
	.A(U_dsdc_n1757));
   NAND2_X2 U_dsdc_U1245 (.ZN(U_dsdc_n1792), 
	.A2(U_dsdc_n590), 
	.A1(U_dsdc_n1799));
   AOI22_X2 U_dsdc_U1244 (.ZN(U_dsdc_n1793), 
	.B2(U_dsdc_n1797), 
	.B1(U_dsdc_num_row[11]), 
	.A2(U_dsdc_n1792), 
	.A1(U_dsdc_row_cnt_11_));
   NAND2_X2 U_dsdc_U1243 (.ZN(U_dsdc_n368), 
	.A2(U_dsdc_n584), 
	.A1(U_dsdc_n1793));
   NAND2_X2 U_dsdc_U1242 (.ZN(U_dsdc_n1763), 
	.A2(U_dsdc_n583), 
	.A1(U_dsdc_n1767));
   AOI22_X2 U_dsdc_U1241 (.ZN(U_dsdc_n1764), 
	.B2(U_dsdc_n1797), 
	.B1(U_dsdc_num_row[7]), 
	.A2(U_dsdc_n1763), 
	.A1(U_dsdc_row_cnt_7_));
   NAND2_X2 U_dsdc_U1240 (.ZN(U_dsdc_n587), 
	.A2(U_dsdc_n579), 
	.A1(U_dsdc_n1791));
   NAND2_X2 U_dsdc_U1239 (.ZN(U_dsdc_n379), 
	.A2(U_dsdc_n587), 
	.A1(U_dsdc_n1764));
   NAND2_X2 U_dsdc_U1238 (.ZN(U_dsdc_n1786), 
	.A2(U_dsdc_n576), 
	.A1(U_dsdc_n1790));
   AOI22_X2 U_dsdc_U1237 (.ZN(U_dsdc_n1787), 
	.B2(U_dsdc_n1797), 
	.B1(U_dsdc_num_row[13]), 
	.A2(U_dsdc_n1786), 
	.A1(U_dsdc_row_cnt_13_));
   NAND2_X2 U_dsdc_U1236 (.ZN(U_dsdc_n588), 
	.A2(U_dsdc_n585), 
	.A1(U_dsdc_n1791));
   NAND2_X2 U_dsdc_U1235 (.ZN(U_dsdc_n370), 
	.A2(U_dsdc_n588), 
	.A1(U_dsdc_n1787));
   NAND2_X2 U_dsdc_U1234 (.ZN(U_dsdc_n1768), 
	.A2(U_dsdc_n591), 
	.A1(U_dsdc_n1773));
   AOI22_X2 U_dsdc_U1233 (.ZN(U_dsdc_n1769), 
	.B2(U_dsdc_n1797), 
	.B1(U_dsdc_num_row[5]), 
	.A2(U_dsdc_n1768), 
	.A1(U_dsdc_row_cnt_5_));
   NAND2_X2 U_dsdc_U1232 (.ZN(U_dsdc_n586), 
	.A2(U_dsdc_n581), 
	.A1(U_dsdc_n1791));
   NAND2_X2 U_dsdc_U1231 (.ZN(U_dsdc_n377), 
	.A2(U_dsdc_n586), 
	.A1(U_dsdc_n1769));
   NAND2_X2 U_dsdc_U1230 (.ZN(U_dsdc_n1759), 
	.A2(U_dsdc_n592), 
	.A1(U_dsdc_n1762));
   AOI22_X2 U_dsdc_U1229 (.ZN(U_dsdc_n1760), 
	.B2(U_dsdc_n1797), 
	.B1(U_dsdc_num_row[9]), 
	.A2(U_dsdc_n1759), 
	.A1(U_dsdc_row_cnt_9_));
   NAND2_X2 U_dsdc_U1228 (.ZN(U_dsdc_n381), 
	.A2(U_dsdc_n589), 
	.A1(U_dsdc_n1760));
   INV_X4 U_dsdc_U1227 (.ZN(U_dsdc_n1722), 
	.A(U_dsdc_n1676));
   AOI21_X2 U_dsdc_U1226 (.ZN(U_dsdc_n1717), 
	.B2(U_dsdc_n1722), 
	.B1(cr_t_init[2]), 
	.A(U_dsdc_n1716));
   OAI21_X2 U_dsdc_U1225 (.ZN(U_dsdc_n405), 
	.B2(U_dsdc_n1718), 
	.B1(U_dsdc_n468), 
	.A(U_dsdc_n1717));
   AOI21_X2 U_dsdc_U1224 (.ZN(U_dsdc_n1780), 
	.B2(U_dsdc_n1791), 
	.B1(U_dsdc_row_cnt_0_), 
	.A(U_dsdc_n1800));
   AOI21_X2 U_dsdc_U1223 (.ZN(U_dsdc_n1779), 
	.B2(U_dsdc_n1797), 
	.B1(U_dsdc_n598), 
	.A(U_dsdc_n325));
   OAI21_X2 U_dsdc_U1222 (.ZN(U_dsdc_n373), 
	.B2(U_dsdc_n465), 
	.B1(U_dsdc_n1780), 
	.A(U_dsdc_n1779));
   OAI211_X2 U_dsdc_U1221 (.ZN(U_dsdc_n1324), 
	.C2(U_dsdc_n1322), 
	.C1(U_dsdc_n1326), 
	.B(U_dsdc_n1321), 
	.A(cr_t_rp[2]));
   NAND2_X2 U_dsdc_U1220 (.ZN(U_dsdc_rp_cnt2_nxt[2]), 
	.A2(U_dsdc_n1323), 
	.A1(U_dsdc_n1324));
   NOR3_X2 U_dsdc_U1219 (.ZN(U_dsdc_n1902), 
	.A3(U_dsdc_n1896), 
	.A2(U_dsdc_n1899), 
	.A1(U_dsdc_bm_bank_age_3__2_));
   OAI21_X2 U_dsdc_U1218 (.ZN(U_dsdc_n1903), 
	.B2(U_dsdc_n1902), 
	.B1(U_dsdc_n1908), 
	.A(U_dsdc_n284));
   OAI21_X2 U_dsdc_U1217 (.ZN(U_dsdc_n221), 
	.B2(U_dsdc_n284), 
	.B1(U_dsdc_n1904), 
	.A(U_dsdc_n1903));
   AOI22_X2 U_dsdc_U1216 (.ZN(U_dsdc_n1798), 
	.B2(U_dsdc_n208), 
	.B1(U_dsdc_n1796), 
	.A2(U_dsdc_n1797), 
	.A1(U_dsdc_num_row[10]));
   OAI21_X2 U_dsdc_U1215 (.ZN(U_dsdc_n367), 
	.B2(U_dsdc_n208), 
	.B1(U_dsdc_n1799), 
	.A(U_dsdc_n1798));
   AOI22_X2 U_dsdc_U1214 (.ZN(U_dsdc_n1766), 
	.B2(U_dsdc_n206), 
	.B1(U_dsdc_n593), 
	.A2(U_dsdc_n1797), 
	.A1(U_dsdc_num_row[6]));
   OAI21_X2 U_dsdc_U1213 (.ZN(U_dsdc_n378), 
	.B2(U_dsdc_n206), 
	.B1(U_dsdc_n1767), 
	.A(U_dsdc_n1766));
   AOI22_X2 U_dsdc_U1212 (.ZN(U_dsdc_n1761), 
	.B2(U_dsdc_n205), 
	.B1(U_dsdc_n595), 
	.A2(U_dsdc_n1797), 
	.A1(U_dsdc_num_row[8]));
   OAI21_X2 U_dsdc_U1211 (.ZN(U_dsdc_n380), 
	.B2(U_dsdc_n205), 
	.B1(U_dsdc_n1762), 
	.A(U_dsdc_n1761));
   AOI22_X2 U_dsdc_U1210 (.ZN(U_dsdc_n1772), 
	.B2(U_dsdc_n207), 
	.B1(U_dsdc_n1771), 
	.A2(U_dsdc_n1797), 
	.A1(U_dsdc_num_row[4]));
   OAI21_X2 U_dsdc_U1209 (.ZN(U_dsdc_n376), 
	.B2(U_dsdc_n207), 
	.B1(U_dsdc_n1773), 
	.A(U_dsdc_n1772));
   AOI22_X2 U_dsdc_U1208 (.ZN(U_dsdc_n1784), 
	.B2(U_dsdc_n202), 
	.B1(U_dsdc_n1783), 
	.A2(U_dsdc_n1797), 
	.A1(U_dsdc_num_row[14]));
   OAI21_X2 U_dsdc_U1207 (.ZN(U_dsdc_n371), 
	.B2(U_dsdc_n202), 
	.B1(U_dsdc_n1785), 
	.A(U_dsdc_n1784));
   AOI22_X2 U_dsdc_U1206 (.ZN(U_dsdc_n1789), 
	.B2(U_dsdc_n203), 
	.B1(U_dsdc_n594), 
	.A2(U_dsdc_n1797), 
	.A1(U_dsdc_num_row[12]));
   OAI21_X2 U_dsdc_U1205 (.ZN(U_dsdc_n369), 
	.B2(U_dsdc_n203), 
	.B1(U_dsdc_n1790), 
	.A(U_dsdc_n1789));
   NAND2_X2 U_dsdc_U1204 (.ZN(U_dsdc_n1160), 
	.A2(U_dsdc_n1152), 
	.A1(U_dsdc_n1159));
   OAI21_X2 U_dsdc_U1203 (.ZN(U_dsdc_N4282), 
	.B2(U_dsdc_n1158), 
	.B1(U_dsdc_n1160), 
	.A(U_dsdc_n1157));
   NAND2_X2 U_dsdc_U1202 (.ZN(U_dsdc_n1154), 
	.A2(U_dsdc_bm_ras_cnt_max_2_), 
	.A1(U_dsdc_n1158));
   OAI21_X2 U_dsdc_U1201 (.ZN(U_dsdc_N4283), 
	.B2(U_dsdc_n1160), 
	.B1(FE_PHN1200_U_dsdc_n1161), 
	.A(U_dsdc_n1155));
   OAI221_X2 U_dsdc_U1200 (.ZN(U_dsdc_n220), 
	.C2(U_dsdc_n1898), 
	.C1(U_dsdc_n303), 
	.B2(U_dsdc_n1901), 
	.B1(U_dsdc_bm_bank_age_3__2_), 
	.A(U_dsdc_n1897));
   AOI22_X2 U_dsdc_U1199 (.ZN(U_dsdc_n1710), 
	.B2(U_dsdc_n1722), 
	.B1(cr_t_init[4]), 
	.A2(U_dsdc_n1709), 
	.A1(U_dsdc_init_cnt_4_));
   AOI22_X2 U_dsdc_U1198 (.ZN(U_dsdc_n1696), 
	.B2(U_dsdc_n1722), 
	.B1(cr_t_init[8]), 
	.A2(U_dsdc_n1695), 
	.A1(U_dsdc_init_cnt_8_));
   AOI22_X2 U_dsdc_U1197 (.ZN(U_dsdc_n1689), 
	.B2(U_dsdc_n1722), 
	.B1(cr_t_init[10]), 
	.A2(U_dsdc_n1688), 
	.A1(FE_PHN3268_U_dsdc_init_cnt_10_));
   AOI22_X2 U_dsdc_U1196 (.ZN(U_dsdc_n1703), 
	.B2(U_dsdc_n1722), 
	.B1(cr_t_init[6]), 
	.A2(U_dsdc_n1702), 
	.A1(U_dsdc_init_cnt_6_));
   OAI221_X2 U_dsdc_U1195 (.ZN(U_dsdc_n211), 
	.C2(U_dsdc_n1858), 
	.C1(U_dsdc_n336), 
	.B2(U_dsdc_n1861), 
	.B1(U_dsdc_bm_bank_age_2__2_), 
	.A(U_dsdc_n1857));
   OAI221_X2 U_dsdc_U1194 (.ZN(U_dsdc_n225), 
	.C2(U_dsdc_n1928), 
	.C1(U_dsdc_n337), 
	.B2(U_dsdc_n1931), 
	.B1(U_dsdc_bm_bank_age_1__2_), 
	.A(U_dsdc_n1927));
   INV_X4 U_dsdc_U1193 (.ZN(U_dsdc_n1966), 
	.A(U_dsdc_n1972));
   AOI21_X2 U_dsdc_U1192 (.ZN(U_dsdc_n1960), 
	.B2(U_dsdc_bm_bank_age_0__0_), 
	.B1(U_dsdc_bm_bank_age_0__1_), 
	.A(U_dsdc_n1966));
   AOI211_X2 U_dsdc_U1191 (.ZN(U_dsdc_n1964), 
	.C2(U_dsdc_n1962), 
	.C1(U_dsdc_n2081), 
	.B(U_dsdc_n1960), 
	.A(U_dsdc_n1961));
   OAI221_X2 U_dsdc_U1190 (.ZN(U_dsdc_n1971), 
	.C2(U_dsdc_n1965), 
	.C1(U_dsdc_n334), 
	.B2(U_dsdc_n1966), 
	.B1(U_dsdc_bm_bank_age_0__2_), 
	.A(U_dsdc_n1964));
   NAND3_X2 U_dsdc_U1189 (.ZN(U_dsdc_n1967), 
	.A3(U_dsdc_n1972), 
	.A2(U_dsdc_bm_bank_age_0__0_), 
	.A1(U_dsdc_bm_bank_age_0__1_));
   NOR2_X2 U_dsdc_U1188 (.ZN(U_dsdc_n1973), 
	.A2(U_dsdc_n1967), 
	.A1(U_dsdc_n334));
   NAND3_X2 U_dsdc_U1187 (.ZN(U_dsdc_n410), 
	.A3(U_dsdc_n1698), 
	.A2(U_dsdc_n1699), 
	.A1(U_dsdc_n1700));
   NAND3_X2 U_dsdc_U1186 (.ZN(U_dsdc_n412), 
	.A3(U_dsdc_n1691), 
	.A2(U_dsdc_n1692), 
	.A1(U_dsdc_n1693));
   NAND3_X2 U_dsdc_U1185 (.ZN(U_dsdc_n408), 
	.A3(U_dsdc_n1705), 
	.A2(U_dsdc_n1706), 
	.A1(U_dsdc_n1707));
   OAI211_X2 U_dsdc_U1184 (.ZN(U_dsdc_n1713), 
	.C2(U_dsdc_n1711), 
	.C1(U_dsdc_init_cnt_2_), 
	.B(U_dsdc_n1715), 
	.A(FE_PHN1062_U_dsdc_init_cnt_3_));
   NAND3_X2 U_dsdc_U1183 (.ZN(U_dsdc_n406), 
	.A3(U_dsdc_n1712), 
	.A2(U_dsdc_n1713), 
	.A1(U_dsdc_n1714));
   NOR3_X2 U_dsdc_U1182 (.ZN(U_dsdc_n1968), 
	.A3(U_dsdc_n1962), 
	.A2(U_dsdc_n1965), 
	.A1(U_dsdc_bm_bank_age_0__2_));
   OAI221_X2 U_dsdc_U1181 (.ZN(U_dsdc_n229), 
	.C2(U_dsdc_n1964), 
	.C1(U_dsdc_n334), 
	.B2(U_dsdc_n1967), 
	.B1(U_dsdc_bm_bank_age_0__2_), 
	.A(U_dsdc_n1963));
   OAI221_X2 U_dsdc_U1180 (.ZN(U_dsdc_n223), 
	.C2(U_dsdc_n1921), 
	.C1(FE_PHN897_U_dsdc_n352), 
	.B2(U_dsdc_n1919), 
	.B1(U_dsdc_bm_bank_age_1__0_), 
	.A(FE_PHN4246_U_dsdc_n356));
   OAI221_X2 U_dsdc_U1179 (.ZN(U_dsdc_n218), 
	.C2(U_dsdc_n1891), 
	.C1(U_dsdc_n304), 
	.B2(U_dsdc_n1889), 
	.B1(U_dsdc_bm_bank_age_3__0_), 
	.A(FE_PHN4075_U_dsdc_n185));
   OAI21_X2 U_dsdc_U1178 (.ZN(U_dsdc_n1969), 
	.B2(U_dsdc_n1968), 
	.B1(U_dsdc_n1973), 
	.A(U_dsdc_n458));
   OAI21_X2 U_dsdc_U1177 (.ZN(U_dsdc_n230), 
	.B2(U_dsdc_n458), 
	.B1(U_dsdc_n1970), 
	.A(U_dsdc_n1969));
   OAI221_X2 U_dsdc_U1176 (.ZN(U_dsdc_n209), 
	.C2(U_dsdc_n1851), 
	.C1(FE_PHN958_U_dsdc_n353), 
	.B2(U_dsdc_n1848), 
	.B1(U_dsdc_bm_bank_age_2__0_), 
	.A(U_dsdc_n164));
   OAI221_X2 U_dsdc_U1175 (.ZN(U_dsdc_n283), 
	.C2(U_dsdc_n2084), 
	.C1(FE_PHN3235_U_dsdc_n201), 
	.B2(U_dsdc_n2085), 
	.B1(U_dsdc_bm_bank_age_0__0_), 
	.A(U_dsdc_n168));
   AOI22_X2 U_dsdc_U1174 (.ZN(U_dsdc_n1681), 
	.B2(U_dsdc_n1722), 
	.B1(cr_t_init[12]), 
	.A2(U_dsdc_n1680), 
	.A1(U_dsdc_init_cnt_12_));
   INV_X4 U_dsdc_U1173 (.ZN(U_dsdc_n287), 
	.A(U_dsdc_n765));
   AOI21_X2 U_dsdc_U1170 (.ZN(U_dsdc_n1339), 
	.B2(hiu_burst_size[0]), 
	.B1(U_dsdc_n1270), 
	.A(U_dsdc_n1261));
   NAND2_X2 U_dsdc_U1169 (.ZN(U_dsdc_n1282), 
	.A2(FE_PHN1335_U_dsdc_n1281), 
	.A1(FE_PHN1161_U_dsdc_n1339));
   OAI21_X2 U_dsdc_U1168 (.ZN(U_dsdc_n1279), 
	.B2(U_dsdc_n1263), 
	.B1(U_dsdc_n1266), 
	.A(U_dsdc_n1262));
   NOR2_X2 U_dsdc_U1167 (.ZN(U_dsdc_n1278), 
	.A2(U_dsdc_n1279), 
	.A1(U_dsdc_n1282));
   NAND2_X2 U_dsdc_U1166 (.ZN(U_dsdc_n1273), 
	.A2(FE_PHN1343_U_dsdc_n1276), 
	.A1(U_dsdc_n1278));
   OAI21_X2 U_dsdc_U1165 (.ZN(U_dsdc_n1274), 
	.B2(U_dmc_n16), 
	.B1(U_dsdc_n1266), 
	.A(U_dsdc_n1264));
   NOR2_X2 U_dsdc_U1164 (.ZN(U_dsdc_n1272), 
	.A2(U_dsdc_n1274), 
	.A1(U_dsdc_n1273));
   NOR2_X2 U_dsdc_U1163 (.ZN(U_dsdc_cas_cnt_nxt[5]), 
	.A2(U_dsdc_n1340), 
	.A1(U_dsdc_n1271));
   AOI21_X2 U_dsdc_U1162 (.ZN(U_dsdc_n1275), 
	.B2(U_dsdc_n1273), 
	.B1(U_dsdc_n1274), 
	.A(U_dsdc_n1272));
   NOR2_X2 U_dsdc_U1161 (.ZN(U_dsdc_cas_cnt_nxt[4]), 
	.A2(U_dsdc_n1340), 
	.A1(FE_PHN1101_U_dsdc_n1275));
   OAI22_X2 U_dsdc_U1160 (.ZN(U_dsdc_N4281), 
	.B2(n95), 
	.B1(U_dsdc_n1159), 
	.A2(FE_PHN2034_U_dsdc_bm_ras_cnt_max_0_), 
	.A1(U_dsdc_n1160));
   AOI21_X2 U_dsdc_U1159 (.ZN(U_dsdc_n1721), 
	.B2(U_dsdc_init_cnt_0_), 
	.B1(U_dsdc_init_cnt_1_), 
	.A(U_dsdc_n1719));
   NAND2_X2 U_dsdc_U1158 (.ZN(U_dsdc_n1720), 
	.A2(U_dsdc_n1722), 
	.A1(cr_t_init[1]));
   NAND2_X2 U_dsdc_U1157 (.ZN(U_dsdc_n1723), 
	.A2(U_dsdc_n1722), 
	.A1(FE_PHN3041_cr_t_init_0_));
   NOR3_X2 U_dsdc_U1154 (.ZN(ctl_mode_reg_done), 
	.A3(U_dsdc_n1521), 
	.A2(U_dsdc_n1490), 
	.A1(FE_PHN791_U_dsdc_n1491));
   NOR3_X2 U_dsdc_U1153 (.ZN(ctl_ext_mode_reg_done), 
	.A3(U_dsdc_n1521), 
	.A2(U_dsdc_n1506), 
	.A1(FE_PHN791_U_dsdc_n1491));
   NOR2_X2 U_dsdc_U1152 (.ZN(U_dsdc_cas_cnt_nxt[3]), 
	.A2(U_dsdc_n1340), 
	.A1(U_dsdc_n1277));
   AOI21_X2 U_dsdc_U1151 (.ZN(U_dsdc_n1280), 
	.B2(U_dsdc_n1282), 
	.B1(U_dsdc_n1279), 
	.A(U_dsdc_n1278));
   NOR2_X2 U_dsdc_U1150 (.ZN(U_dsdc_cas_cnt_nxt[2]), 
	.A2(U_dsdc_n1340), 
	.A1(U_dsdc_n1280));
   AOI21_X2 U_dsdc_U1149 (.ZN(U_dsdc_n1630), 
	.B2(U_dsdc_n1419), 
	.B1(U_dsdc_n1414), 
	.A(U_dsdc_n1629));
   AOI211_X2 U_dsdc_U1148 (.ZN(U_dsdc_n1635), 
	.C2(U_dsdc_n1420), 
	.C1(U_dsdc_n1632), 
	.B(U_dsdc_n1630), 
	.A(U_dsdc_n1631));
   NOR3_X2 U_dsdc_U1147 (.ZN(U_dsdc_n1648), 
	.A3(U_dsdc_n1632), 
	.A2(U_dsdc_n1633), 
	.A1(U_dsdc_n1414));
   OAI21_X2 U_dsdc_U1146 (.ZN(U_dsdc_n1639), 
	.B2(U_dsdc_n1635), 
	.B1(U_dsdc_n1424), 
	.A(U_dsdc_n1634));
   NAND2_X2 U_dsdc_U1145 (.ZN(U_dsdc_n1636), 
	.A2(U_dsdc_n1872), 
	.A1(U_dsdc_n1414));
   INV_X4 U_dsdc_U1144 (.ZN(U_dsdc_n1642), 
	.A(U_dsdc_n1636));
   NOR2_X2 U_dsdc_U1143 (.ZN(U_dsdc_n1646), 
	.A2(U_dsdc_n1642), 
	.A1(U_dsdc_n1639));
   AOI22_X2 U_dsdc_U1142 (.ZN(U_dsdc_n1643), 
	.B2(U_dsdc_n1639), 
	.B1(U_dsdc_n1640), 
	.A2(U_dsdc_n1641), 
	.A1(U_dsdc_n1642));
   OAI21_X2 U_dsdc_U1141 (.ZN(U_dsdc_n1647), 
	.B2(U_dsdc_n200), 
	.B1(U_dsdc_n1646), 
	.A(U_dsdc_n1643));
   NOR2_X2 U_dsdc_U1140 (.ZN(U_dsdc_n1379), 
	.A2(U_dsdc_n1359), 
	.A1(U_dsdc_n1876));
   NOR3_X2 U_dsdc_U1137 (.ZN(U_dsdc_n1649), 
	.A3(U_dsdc_n1636), 
	.A2(U_dsdc_n1640), 
	.A1(U_dsdc_n1444));
   OAI21_X2 U_dsdc_U1136 (.ZN(U_dsdc_n2073), 
	.B2(U_dsdc_n2069), 
	.B1(U_dsdc_n1419), 
	.A(U_dsdc_n1398));
   INV_X4 U_dsdc_U1135 (.ZN(U_dsdc_n708), 
	.A(U_dsdc_n901));
   NOR2_X2 U_dsdc_U1134 (.ZN(U_dsdc_n1875), 
	.A2(U_dsdc_n1416), 
	.A1(U_dsdc_n708));
   NOR2_X2 U_dsdc_U1133 (.ZN(U_dsdc_n1880), 
	.A2(U_dsdc_n1881), 
	.A1(U_dsdc_n461));
   AOI21_X2 U_dsdc_U1132 (.ZN(U_dsdc_n2072), 
	.B2(U_dsdc_n1871), 
	.B1(U_dsdc_n1425), 
	.A(U_dsdc_n2073));
   OAI21_X2 U_dsdc_U1129 (.ZN(U_dsdc_n1879), 
	.B2(U_dsdc_n1875), 
	.B1(U_dsdc_delta_delay_0_), 
	.A(U_dsdc_n183));
   AOI21_X2 U_dsdc_U1128 (.ZN(U_dsdc_n1878), 
	.B2(U_dsdc_n464), 
	.B1(U_dsdc_n1874), 
	.A(U_dsdc_n1879));
   NAND2_X2 U_dsdc_U1127 (.ZN(U_dsdc_n1877), 
	.A2(U_dsdc_n1880), 
	.A1(U_dsdc_delta_delay_1_));
   AOI22_X2 U_dsdc_U1126 (.ZN(U_dsdc_n214), 
	.B2(U_dsdc_n467), 
	.B1(U_dsdc_n1877), 
	.A2(U_dsdc_n1878), 
	.A1(U_dsdc_delta_delay_2_));
   AOI211_X2 U_dsdc_U1125 (.ZN(U_dsdc_n1488), 
	.C2(U_dsdc_operation_cs_0_), 
	.C1(U_dsdc_n1487), 
	.B(U_dsdc_n1486), 
	.A(U_dsdc_n1429));
   AOI21_X2 U_dsdc_U1124 (.ZN(U_dsdc_n1645), 
	.B2(U_dsdc_n1639), 
	.B1(U_dsdc_n1638), 
	.A(U_dsdc_n1649));
   NOR2_X2 U_dsdc_U1123 (.ZN(U_dsdc_n770), 
	.A2(U_dsdc_n1414), 
	.A1(U_dsdc_n1359));
   AOI211_X2 U_dsdc_U1121 (.ZN(U_dsdc_n1976), 
	.C2(U_dsdc_n1975), 
	.C1(U_dsdc_n1427), 
	.B(U_dsdc_n1974), 
	.A(U_dsdc_n1425));
   NAND3_X2 U_dsdc_U1120 (.ZN(U_dsdc_n713), 
	.A3(U_dsdc_n1976), 
	.A2(U_dsdc_n1397), 
	.A1(U_dsdc_n869));
   NOR2_X2 U_dsdc_U1119 (.ZN(U_dsdc_n1396), 
	.A2(U_dsdc_n1802), 
	.A1(U_dsdc_n713));
   INV_X4 U_dsdc_U1118 (.ZN(U_dsdc_n718), 
	.A(U_dsdc_n956));
   NAND2_X2 U_dsdc_U1117 (.ZN(U_dsdc_n2067), 
	.A2(U_dsdc_n718), 
	.A1(U_dsdc_n1396));
   NOR2_X2 U_dsdc_U1116 (.ZN(U_dsdc_n1395), 
	.A2(U_dsdc_n1411), 
	.A1(U_dsdc_n2067));
   NAND2_X2 U_dsdc_U1115 (.ZN(U_dsdc_n280), 
	.A2(U_dsdc_n1346), 
	.A1(U_dsdc_n1347));
   AOI22_X2 U_dsdc_U1114 (.ZN(U_dsdc_n773), 
	.B2(U_dsdc_n770), 
	.B1(U_dsdc_r_cas_latency_3_), 
	.A2(U_dsdc_n1379), 
	.A1(U_dsdc_N2002));
   NAND2_X2 U_dsdc_U1113 (.ZN(U_dsdc_n772), 
	.A2(U_dsdc_N1990), 
	.A1(n89));
   OAI211_X2 U_dsdc_U1112 (.ZN(U_dsdc_n774), 
	.C2(U_dsdc_n1644), 
	.C1(U_dsdc_n1645), 
	.B(U_dsdc_n772), 
	.A(U_dsdc_n773));
   AOI21_X2 U_dsdc_U1111 (.ZN(U_dsdc_n775), 
	.B2(U_dsdc_term_cnt_3_), 
	.B1(U_dsdc_n1647), 
	.A(U_dsdc_n774));
   INV_X4 U_dsdc_U1110 (.ZN(U_dsdc_term_cnt_nxt[3]), 
	.A(U_dsdc_n775));
   NAND2_X2 U_dsdc_U1109 (.ZN(U_dsdc_n418), 
	.A2(U_dsdc_n1673), 
	.A1(U_dsdc_n1674));
   NAND2_X2 U_dsdc_U1108 (.ZN(U_dsdc_n717), 
	.A2(U_dsdc_n759), 
	.A1(U_dsdc_n879));
   NOR2_X2 U_dsdc_U1081 (.ZN(U_dsdc_cas_cnt_nxt[0]), 
	.A2(U_dsdc_n1340), 
	.A1(U_dsdc_n1341));
   NAND3_X2 U_dsdc_U1080 (.ZN(U_dsdc_n676), 
	.A3(U_dsdc_n674), 
	.A2(U_dsdc_n675), 
	.A1(U_dsdc_n717));
   AOI22_X2 U_dsdc_U1076 (.ZN(U_dsdc_n1742), 
	.B2(U_dsdc_n1754), 
	.B1(cr_t_xsr[4]), 
	.A2(U_dsdc_n1741), 
	.A1(U_dsdc_xsr_cnt_4_));
   OAI21_X2 U_dsdc_U1075 (.ZN(U_dsdc_n390), 
	.B2(U_dsdc_n1744), 
	.B1(U_dsdc_xsr_cnt_4_), 
	.A(U_dsdc_n1742));
   AOI22_X2 U_dsdc_U1070 (.ZN(U_dsdc_n1813), 
	.B2(U_dsdc_n1817), 
	.B1(U_dsdc_n354), 
	.A2(U_dsdc_n1815), 
	.A1(debug_ad_col_addr_1_));
   NAND2_X2 U_dsdc_U1069 (.ZN(U_dsdc_n319), 
	.A2(U_dsdc_n1812), 
	.A1(U_dsdc_n1813));
   NOR2_X2 U_dsdc_U1061 (.ZN(U_dsdc_n1747), 
	.A2(FE_PHN1033_U_dsdc_xsr_cnt_1_), 
	.A1(U_dsdc_xsr_cnt_0_));
   NAND2_X2 U_dsdc_U1060 (.ZN(U_dsdc_n1751), 
	.A2(U_dsdc_n1750), 
	.A1(U_dsdc_n1747));
   NOR2_X2 U_dsdc_U1059 (.ZN(U_dsdc_n1748), 
	.A2(U_dsdc_n1756), 
	.A1(U_dsdc_n1747));
   AOI22_X2 U_dsdc_U1058 (.ZN(U_dsdc_n1749), 
	.B2(U_dsdc_n1754), 
	.B1(cr_t_xsr[2]), 
	.A2(U_dsdc_n1748), 
	.A1(U_dsdc_xsr_cnt_2_));
   OAI21_X2 U_dsdc_U1057 (.ZN(U_dsdc_n388), 
	.B2(U_dsdc_n1751), 
	.B1(U_dsdc_xsr_cnt_2_), 
	.A(U_dsdc_n1749));
   AOI22_X2 U_dsdc_U1046 (.ZN(U_dsdc_n2025), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_11_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[11]));
   INV_X4 U_dsdc_U1045 (.ZN(U_dsdc_n257), 
	.A(U_dsdc_n2025));
   AOI22_X2 U_dsdc_U1044 (.ZN(U_dsdc_n2024), 
	.B2(U_dsdc_n2038), 
	.B1(FE_PHN1148_U_dsdc_r_row_addr_10_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[10]));
   INV_X4 U_dsdc_U1043 (.ZN(U_dsdc_n256), 
	.A(U_dsdc_n2024));
   AOI22_X2 U_dsdc_U1042 (.ZN(U_dsdc_n2023), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_0_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[0]));
   INV_X4 U_dsdc_U1041 (.ZN(U_dsdc_n255), 
	.A(U_dsdc_n2023));
   AOI22_X2 U_dsdc_U1040 (.ZN(U_dsdc_n2029), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_15_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[15]));
   INV_X4 U_dsdc_U1039 (.ZN(U_dsdc_n261), 
	.A(U_dsdc_n2029));
   AOI22_X2 U_dsdc_U1038 (.ZN(U_dsdc_n2030), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_1_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[1]));
   INV_X4 U_dsdc_U1037 (.ZN(U_dsdc_n262), 
	.A(U_dsdc_n2030));
   AOI22_X2 U_dsdc_U1036 (.ZN(U_dsdc_n2031), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_2_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[2]));
   INV_X4 U_dsdc_U1035 (.ZN(U_dsdc_n263), 
	.A(U_dsdc_n2031));
   AOI22_X2 U_dsdc_U1034 (.ZN(U_dsdc_n2032), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_3_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[3]));
   INV_X4 U_dsdc_U1033 (.ZN(U_dsdc_n264), 
	.A(U_dsdc_n2032));
   AOI22_X2 U_dsdc_U1032 (.ZN(U_dsdc_n2033), 
	.B2(U_dsdc_n2038), 
	.B1(FE_PHN1147_U_dsdc_r_row_addr_4_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[4]));
   INV_X4 U_dsdc_U1031 (.ZN(U_dsdc_n265), 
	.A(U_dsdc_n2033));
   AOI22_X2 U_dsdc_U1030 (.ZN(U_dsdc_n2028), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_14_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[14]));
   INV_X4 U_dsdc_U1029 (.ZN(U_dsdc_n260), 
	.A(U_dsdc_n2028));
   AOI22_X2 U_dsdc_U1028 (.ZN(U_dsdc_n2035), 
	.B2(U_dsdc_n2038), 
	.B1(FE_PHN1146_U_dsdc_r_row_addr_6_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[6]));
   INV_X4 U_dsdc_U1027 (.ZN(U_dsdc_n267), 
	.A(U_dsdc_n2035));
   AOI22_X2 U_dsdc_U1026 (.ZN(U_dsdc_n2037), 
	.B2(U_dsdc_n2038), 
	.B1(FE_PHN1151_U_dsdc_r_row_addr_8_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[8]));
   INV_X4 U_dsdc_U1025 (.ZN(U_dsdc_n269), 
	.A(U_dsdc_n2037));
   AOI22_X2 U_dsdc_U1024 (.ZN(U_dsdc_n2040), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_9_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[9]));
   INV_X4 U_dsdc_U1023 (.ZN(U_dsdc_n270), 
	.A(U_dsdc_n2040));
   AOI22_X2 U_dsdc_U1022 (.ZN(U_dsdc_n2026), 
	.B2(FE_OFN303_U_dsdc_n2038), 
	.B1(FE_PHN1149_U_dsdc_r_row_addr_12_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[12]));
   INV_X4 U_dsdc_U1021 (.ZN(U_dsdc_n258), 
	.A(U_dsdc_n2026));
   AOI22_X2 U_dsdc_U1020 (.ZN(U_dsdc_n2034), 
	.B2(U_dsdc_n2038), 
	.B1(FE_PHN1152_U_dsdc_r_row_addr_5_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[5]));
   INV_X4 U_dsdc_U1019 (.ZN(U_dsdc_n266), 
	.A(U_dsdc_n2034));
   AOI22_X2 U_dsdc_U1018 (.ZN(U_dsdc_n2027), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_13_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[13]));
   INV_X4 U_dsdc_U1017 (.ZN(U_dsdc_n259), 
	.A(U_dsdc_n2027));
   AOI22_X2 U_dsdc_U1016 (.ZN(U_dsdc_n2036), 
	.B2(U_dsdc_n2038), 
	.B1(U_dsdc_r_row_addr_7_), 
	.A2(U_dsdc_n2039), 
	.A1(debug_ad_row_addr[7]));
   INV_X4 U_dsdc_U1015 (.ZN(U_dsdc_n268), 
	.A(U_dsdc_n2036));
   AOI22_X2 U_dsdc_U1014 (.ZN(U_dsdc_n216), 
	.B2(U_dsdc_n461), 
	.B1(U_dsdc_n1881), 
	.A2(U_dsdc_n183), 
	.A1(U_dsdc_delta_delay_0_));
   NOR3_X2 U_dsdc_U1013 (.ZN(U_dsdc_n2075), 
	.A3(U_dsdc_n2070), 
	.A2(U_dsdc_n1412), 
	.A1(U_dsdc_n1416));
   NAND2_X2 U_dsdc_U1012 (.ZN(U_dsdc_n2049), 
	.A2(U_dsdc_n1396), 
	.A1(U_dsdc_n2041));
   NOR4_X2 U_dsdc_U1011 (.ZN(U_dsdc_N4174), 
	.A4(U_dsdc_n1670), 
	.A3(FE_PHN1081_U_dsdc_n1671), 
	.A2(U_dsdc_n1430), 
	.A1(U_dsdc_mrd_cnt_0_));
   AOI211_X2 U_dsdc_U1010 (.ZN(U_dsdc_n1672), 
	.C2(U_dsdc_mrd_cnt_0_), 
	.C1(U_dsdc_mrd_cnt_1_), 
	.B(U_dsdc_n1670), 
	.A(FE_PHN1081_U_dsdc_n1671));
   INV_X4 U_dsdc_U1009 (.ZN(U_dsdc_n423), 
	.A(U_dsdc_n1672));
   AOI22_X2 U_dsdc_U1008 (.ZN(U_dsdc_n279), 
	.B2(U_dsdc_n2068), 
	.B1(FE_PHN1887_U_dsdc_n166), 
	.A2(U_dsdc_n1438), 
	.A1(U_dsdc_n1395));
   NAND3_X2 U_dsdc_U1007 (.ZN(U_dsdc_n389), 
	.A3(U_dsdc_n1744), 
	.A2(U_dsdc_n1745), 
	.A1(U_dsdc_n1746));
   NAND2_X2 U_dsdc_U1006 (.ZN(U_dsdc_n391), 
	.A2(U_dsdc_n1738), 
	.A1(U_dsdc_n1739));
   OAI21_X2 U_dsdc_U1005 (.ZN(U_dsdc_n282), 
	.B2(U_dsdc_n2078), 
	.B1(U_dsdc_n2079), 
	.A(U_dsdc_n2077));
   NAND3_X2 U_dsdc_U1004 (.ZN(U_dsdc_n387), 
	.A3(U_dsdc_n1751), 
	.A2(U_dsdc_n1752), 
	.A1(U_dsdc_n1753));
   NAND2_X2 U_dsdc_U1003 (.ZN(U_dsdc_n1734), 
	.A2(U_dsdc_n1750), 
	.A1(U_dsdc_n1729));
   NAND2_X2 U_dsdc_U1002 (.ZN(U_dsdc_n392), 
	.A2(U_dsdc_n1734), 
	.A1(U_dsdc_n1735));
   NOR2_X2 U_dsdc_U1001 (.ZN(U_dsdc_n1597), 
	.A2(U_dsdc_n1591), 
	.A1(U_dsdc_n1592));
   INV_X4 U_dsdc_U1000 (.ZN(U_dsdc_n1609), 
	.A(U_dsdc_n1597));
   NAND2_X2 U_dsdc_U999 (.ZN(U_dsdc_n1615), 
	.A2(U_dsdc_n1609), 
	.A1(U_dsdc_rcar_cnt2_3_));
   NAND2_X2 U_dsdc_U998 (.ZN(U_dsdc_n1603), 
	.A2(FE_PHN1482_U_cr_n151), 
	.A1(FE_PHN1052_U_cr_n127));
   NAND2_X2 U_dsdc_U997 (.ZN(U_dsdc_n1593), 
	.A2(FE_PHN1407_U_cr_n104), 
	.A1(FE_PHN1482_U_cr_n151));
   OAI21_X2 U_dsdc_U996 (.ZN(U_dsdc_n1596), 
	.B2(U_dsdc_n1593), 
	.B1(cr_t_rcar[3]), 
	.A(U_dsdc_n1612));
   INV_X4 U_dsdc_U995 (.ZN(U_dsdc_n1602), 
	.A(U_dsdc_n1596));
   AOI21_X2 U_dsdc_U994 (.ZN(U_dsdc_n1610), 
	.B2(U_dsdc_n1602), 
	.B1(U_dsdc_n1603), 
	.A(U_dsdc_n1601));
   AOI21_X2 U_dsdc_U993 (.ZN(U_dsdc_n1614), 
	.B2(FE_PHN3240_cr_t_rcar_2_), 
	.B1(U_dsdc_n1612), 
	.A(U_dsdc_n1611));
   OAI22_X2 U_dsdc_U992 (.ZN(U_dsdc_rcar_cnt2_nxt[3]), 
	.B2(U_cr_n72), 
	.B1(U_dsdc_n1614), 
	.A2(U_dsdc_n1615), 
	.A1(U_dsdc_n1616));
   NAND2_X2 U_dsdc_U991 (.ZN(U_dsdc_n1573), 
	.A2(U_dsdc_n1580), 
	.A1(U_dsdc_n1568));
   NOR3_X2 U_dsdc_U990 (.ZN(U_dsdc_n1666), 
	.A3(U_dsdc_n2063), 
	.A2(FE_PHN843_U_dsdc_num_init_ref_cnt_1_), 
	.A1(U_dsdc_num_init_ref_cnt_0_));
   AOI22_X2 U_dsdc_U989 (.ZN(U_dsdc_n1572), 
	.B2(cr_num_init_ref[2]), 
	.B1(U_dsdc_n1667), 
	.A2(U_dsdc_n1571), 
	.A1(U_dsdc_num_init_ref_cnt_2_));
   OAI21_X2 U_dsdc_U988 (.ZN(U_dsdc_num_init_ref_cnt_nxt[2]), 
	.B2(U_dsdc_n1573), 
	.B1(U_dsdc_num_init_ref_cnt_2_), 
	.A(U_dsdc_n1572));
   NOR2_X2 U_dsdc_U987 (.ZN(U_dsdc_n1604), 
	.A2(U_dsdc_rcar_cnt2_0_), 
	.A1(U_dsdc_rcar_cnt2_1_));
   OAI221_X2 U_dsdc_U986 (.ZN(U_dsdc_rcar_cnt2_nxt[2]), 
	.C2(U_dsdc_n1610), 
	.C1(FE_PHN1407_U_cr_n104), 
	.B2(U_dsdc_n1608), 
	.B1(FE_PHN3240_cr_t_rcar_2_), 
	.A(U_dsdc_n1606));
   AOI21_X2 U_dsdc_U985 (.ZN(U_dsdc_n1668), 
	.B2(U_dsdc_n473), 
	.B1(U_dsdc_n1666), 
	.A(U_dsdc_n2051));
   AOI22_X2 U_dsdc_U984 (.ZN(U_dsdc_n1669), 
	.B2(cr_num_init_ref[3]), 
	.B1(U_dsdc_n1667), 
	.A2(U_dsdc_n1668), 
	.A1(U_dsdc_num_init_ref_cnt_3_));
   INV_X4 U_dsdc_U983 (.ZN(U_dsdc_n431), 
	.A(U_dsdc_n1669));
   AOI22_X2 U_dsdc_U982 (.ZN(U_dsdc_n1594), 
	.B2(FE_PHN1052_U_cr_n127), 
	.B1(U_dsdc_n1602), 
	.A2(U_dsdc_n1601), 
	.A1(cr_t_rcar[0]));
   OAI221_X2 U_dsdc_U981 (.ZN(U_dsdc_n1598), 
	.C2(U_dsdc_rcar_cnt2_1_), 
	.C1(U_dsdc_n1604), 
	.B2(U_dsdc_rcar_cnt2_0_), 
	.B1(U_dsdc_n1604), 
	.A(U_dsdc_n1609));
   OAI211_X2 U_dsdc_U980 (.ZN(U_dsdc_rcar_cnt2_nxt[1]), 
	.C2(FE_PHN1482_U_cr_n151), 
	.C1(U_dsdc_n1600), 
	.B(U_dsdc_n1598), 
	.A(U_dsdc_n1608));
   OAI21_X2 U_dsdc_U979 (.ZN(U_dsdc_num_init_ref_cnt_nxt[0]), 
	.B2(U_dsdc_n1567), 
	.B1(U_dsdc_num_init_ref_cnt_0_), 
	.A(U_dsdc_n1566));
   NAND2_X2 U_dsdc_U978 (.ZN(U_dsdc_n394), 
	.A2(U_dsdc_n1725), 
	.A1(U_dsdc_n1726));
   NAND3_X2 U_dsdc_U977 (.ZN(U_dsdc_num_init_ref_cnt_nxt[1]), 
	.A3(U_dsdc_n1569), 
	.A2(U_dsdc_n1573), 
	.A1(U_dsdc_n1570));
   INV_X4 U_dsdc_U976 (.ZN(U_dsdc_n1622), 
	.A(U_dsdc_n1618));
   NOR2_X2 U_dsdc_U975 (.ZN(U_dsdc_n1624), 
	.A2(FE_PHN3313_U_dsdc_rp_cnt1_0_), 
	.A1(U_dsdc_rp_cnt1_1_));
   AOI21_X2 U_dsdc_U974 (.ZN(U_dsdc_n1620), 
	.B2(U_dsdc_rp_cnt1_1_), 
	.B1(FE_PHN3313_U_dsdc_rp_cnt1_0_), 
	.A(U_dsdc_n1624));
   OAI22_X2 U_dsdc_U973 (.ZN(U_dsdc_rp_cnt1_nxt[1]), 
	.B2(U_dsdc_n1619), 
	.B1(U_dsdc_n1620), 
	.A2(FE_PHN3012_U_cr_n147), 
	.A1(U_dsdc_n1622));
   NAND2_X2 U_dsdc_U972 (.ZN(U_dsdc_n1623), 
	.A2(U_dsdc_n1621), 
	.A1(U_dsdc_rp_cnt1_2_));
   OAI22_X2 U_dsdc_U971 (.ZN(U_dsdc_rp_cnt1_nxt[2]), 
	.B2(FE_PHN3514_U_cr_n148), 
	.B1(U_dsdc_n1622), 
	.A2(U_dsdc_n1623), 
	.A1(U_dsdc_n1624));
   OAI22_X2 U_dsdc_U970 (.ZN(U_dsdc_rp_cnt1_nxt[0]), 
	.B2(FE_PHN3505_U_cr_n45), 
	.B1(U_dsdc_n1622), 
	.A2(U_dsdc_n1619), 
	.A1(FE_PHN3313_U_dsdc_rp_cnt1_0_));
   NOR2_X2 U_dsdc_U969 (.ZN(U_dsdc_n1445), 
	.A2(U_dsdc_access_cs_1_), 
	.A1(U_dsdc_access_cs_3_));
   NOR2_X2 U_dsdc_U968 (.ZN(U_dsdc_n998), 
	.A2(debug_ad_bank_addr[0]), 
	.A1(debug_ad_bank_addr[1]));
   OAI21_X2 U_dsdc_U967 (.ZN(U_dsdc_n1473), 
	.B2(debug_ref_req), 
	.B1(U_dsdc_n1428), 
	.A(U_dsdc_n2056));
   AOI222_X1 U_dsdc_U965 (.ZN(U_dsdc_n1920), 
	.C2(U_dsdc_n1954), 
	.C1(U_dsdc_n349), 
	.B2(U_dsdc_n1954), 
	.B1(U_dsdc_n1917), 
	.A2(U_dsdc_n349), 
	.A1(U_dsdc_n1917));
   NAND2_X2 U_dsdc_U964 (.ZN(U_dsdc_n1315), 
	.A2(U_dsdc_n1411), 
	.A1(U_dsdc_n903));
   NOR2_X1 U_dsdc_U963 (.ZN(U_dsdc_n883), 
	.A2(hiu_rw), 
	.A1(U_dsdc_n1557));
   INV_X1 U_dsdc_U962 (.ZN(U_dsdc_n885), 
	.A(U_dsdc_n884));
   NAND3_X1 U_dsdc_U959 (.ZN(U_dsdc_n1008), 
	.A3(U_dsdc_n180), 
	.A2(U_dsdc_bm_num_open_bank_0_), 
	.A1(U_dsdc_n1166));
   OAI22_X2 U_dsdc_U958 (.ZN(U_dsdc_n1493), 
	.B2(U_dsdc_n2063), 
	.B1(U_dsdc_n1492), 
	.A2(U_dsdc_n1537), 
	.A1(debug_ref_req));
   OAI21_X2 U_dsdc_U957 (.ZN(U_dsdc_n1527), 
	.B2(U_dsdc_n432), 
	.B1(U_dsdc_n1508), 
	.A(U_dsdc_n1507));
   INV_X1 U_dsdc_U955 (.ZN(U_dsdc_n1373), 
	.A(U_dsdc_n1286));
   NOR4_X2 U_dsdc_U954 (.ZN(U_dsdc_n1716), 
	.A4(U_dsdc_n1724), 
	.A3(U_dsdc_init_cnt_2_), 
	.A2(U_dsdc_init_cnt_1_), 
	.A1(U_dsdc_init_cnt_0_));
   INV_X1 U_dsdc_U953 (.ZN(U_dsdc_n1686), 
	.A(U_dsdc_n1679));
   AOI22_X2 U_dsdc_U952 (.ZN(U_dsdc_n1264), 
	.B2(U_dsdc_n1269), 
	.B1(FE_PHN1888_U_dsdc_r_burst_size_4_), 
	.A2(U_dsdc_cas_cnt_4_), 
	.A1(U_dsdc_n1268));
   NAND2_X2 U_dsdc_U949 (.ZN(U_dsdc_n974), 
	.A2(U_dsdc_n1412), 
	.A1(U_dsdc_n891));
   OAI222_X2 U_dsdc_U929 (.ZN(U_dsdc_DP_OP_1642_126_2028_I5_0_), 
	.C2(U_dsdc_n1253), 
	.C1(U_dsdc_n1546), 
	.B2(U_dsdc_n601), 
	.B1(U_dsdc_n347), 
	.A2(U_dsdc_n1258), 
	.A1(U_dsdc_n182));
   INV_X1 U_dsdc_U928 (.ZN(U_dsdc_n572), 
	.A(U_dsdc_n998));
   AOI21_X1 U_dsdc_U924 (.ZN(U_dsdc_n848), 
	.B2(U_dsdc_n976), 
	.B1(U_dsdc_n910), 
	.A(U_dsdc_n836));
   INV_X1 U_dsdc_U923 (.ZN(U_dsdc_n574), 
	.A(U_dsdc_n1776));
   INV_X1 U_dsdc_U922 (.ZN(U_dsdc_n1130), 
	.A(debug_ad_bank_addr[1]));
   INV_X1 U_dsdc_U921 (.ZN(U_dsdc_n580), 
	.A(U_dsdc_n1794));
   INV_X1 U_dsdc_U920 (.ZN(U_dsdc_n579), 
	.A(U_dsdc_n1765));
   INV_X1 U_dsdc_U919 (.ZN(U_dsdc_n581), 
	.A(U_dsdc_n1770));
   INV_X1 U_dsdc_U918 (.ZN(U_dsdc_n575), 
	.A(U_dsdc_n1795));
   NOR2_X2 U_dsdc_U917 (.ZN(U_dsdc_n2041), 
	.A2(U_dsdc_n676), 
	.A1(U_dsdc_n716));
   NAND2_X1 U_dsdc_U915 (.ZN(U_dsdc_n666), 
	.A2(U_dsdc_n1445), 
	.A1(U_dsdc_n167));
   NAND2_X2 U_dsdc_U914 (.ZN(U_dsdc_n1136), 
	.A2(U_dsdc_n1384), 
	.A1(U_dsdc_n1422));
   INV_X4 U_dsdc_U913 (.ZN(U_dsdc_n619), 
	.A(U_dsdc_n184));
   OAI21_X2 U_dsdc_U911 (.ZN(U_dsdc_n1671), 
	.B2(U_dsdc_n1509), 
	.B1(U_dsdc_n643), 
	.A(U_dsdc_n1513));
   NOR4_X2 U_dsdc_U910 (.ZN(U_dsdc_n1804), 
	.A4(U_dsdc_n1802), 
	.A3(U_dsdc_n1418), 
	.A2(U_dsdc_n1427), 
	.A1(U_dsdc_n1411));
   NOR4_X1 U_dsdc_U908 (.ZN(U_dsdc_N4239), 
	.A4(FE_PHN1064_cr_row_addr_width_3_), 
	.A3(FE_PHN3054_cr_row_addr_width_2_), 
	.A2(cr_row_addr_width[0]), 
	.A1(cr_row_addr_width[1]));
   OAI22_X1 U_dsdc_U907 (.ZN(U_dsdc_bm_close_bank_3_), 
	.B2(U_dsdc_n1390), 
	.B1(U_dsdc_n999), 
	.A2(U_dsdc_n987), 
	.A1(U_dsdc_n1391));
   OAI22_X1 U_dsdc_U906 (.ZN(U_dsdc_bm_close_bank_2_), 
	.B2(U_dsdc_n1390), 
	.B1(U_dsdc_oldest_bank_0_), 
	.A2(U_dsdc_n599), 
	.A1(U_dsdc_n1391));
   AOI21_X1 U_dsdc_U905 (.ZN(U_dsdc_n1799), 
	.B2(U_dsdc_n1795), 
	.B1(U_dsdc_n1791), 
	.A(U_dsdc_n1800));
   AOI21_X1 U_dsdc_U904 (.ZN(U_dsdc_n1767), 
	.B2(U_dsdc_n1770), 
	.B1(U_dsdc_n1791), 
	.A(U_dsdc_n1800));
   AOI21_X1 U_dsdc_U903 (.ZN(U_dsdc_n1790), 
	.B2(U_dsdc_n1794), 
	.B1(U_dsdc_n1791), 
	.A(U_dsdc_n1800));
   AOI21_X1 U_dsdc_U902 (.ZN(U_dsdc_n1773), 
	.B2(U_dsdc_n1776), 
	.B1(U_dsdc_n1791), 
	.A(U_dsdc_n1800));
   AOI21_X1 U_dsdc_U901 (.ZN(U_dsdc_n1762), 
	.B2(U_dsdc_n1765), 
	.B1(U_dsdc_n1791), 
	.A(U_dsdc_n1800));
   INV_X4 U_dsdc_U900 (.ZN(U_dsdc_n1715), 
	.A(U_dsdc_n1724));
   AOI21_X2 U_dsdc_U899 (.ZN(U_dsdc_n2039), 
	.B2(U_dsdc_n2013), 
	.B1(FE_OFN304_U_dsdc_n2014), 
	.A(U_dsdc_n2067));
   OAI21_X2 U_dsdc_U898 (.ZN(U_dsdc_n2038), 
	.B2(U_dsdc_n1309), 
	.B1(U_dsdc_n891), 
	.A(U_dsdc_n720));
   OAI221_X2 U_dsdc_U897 (.ZN(U_dsdc_n1606), 
	.C2(U_dsdc_n1605), 
	.C1(U_dsdc_n1616), 
	.B2(U_dsdc_rcar_cnt2_2_), 
	.B1(U_dsdc_n1616), 
	.A(U_dsdc_n1609));
   NOR2_X2 U_dsdc_U895 (.ZN(U_dsdc_n1412), 
	.A2(U_dsdc_n666), 
	.A1(U_dsdc_n667));
   NAND2_X2 U_dsdc_U894 (.ZN(U_dsdc_n501), 
	.A2(U_dsdc_bm_row_addr_0__6_), 
	.A1(U_dsdc_n998));
   NOR2_X2 U_dsdc_U893 (.ZN(U_dsdc_n891), 
	.A2(U_dsdc_n759), 
	.A1(U_dsdc_n903));
   NOR2_X1 U_dsdc_U892 (.ZN(U_dsdc_n1416), 
	.A2(U_dsdc_access_cs_0_), 
	.A1(U_dsdc_n741));
   NAND4_X2 U_dsdc_U891 (.ZN(U_dsdc_n1633), 
	.A4(U_dsdc_n1445), 
	.A3(U_dsdc_access_cs_0_), 
	.A2(U_dsdc_access_cs_2_), 
	.A1(U_dsdc_n167));
   NAND3_X1 U_dsdc_U890 (.ZN(U_dsdc_n2062), 
	.A3(U_dsdc_n1577), 
	.A2(U_dsdc_n1478), 
	.A1(cr_do_self_ref_rp));
   AOI22_X2 U_dsdc_U889 (.ZN(U_dsdc_n2085), 
	.B2(U_dsdc_n2080), 
	.B1(U_dsdc_n2081), 
	.A2(U_dsdc_n2082), 
	.A1(U_dsdc_bm_bank_status_0_));
   AOI22_X2 U_dsdc_U887 (.ZN(U_dsdc_n1739), 
	.B2(U_dsdc_n1754), 
	.B1(cr_t_xsr[5]), 
	.A2(U_dsdc_n1750), 
	.A1(U_dsdc_n1736));
   NAND2_X1 U_dsdc_U886 (.ZN(U_dsdc_n2014), 
	.A2(U_dsdc_n167), 
	.A1(U_dsdc_n964));
   AOI21_X2 U_dsdc_U884 (.ZN(U_dsdc_n977), 
	.B2(U_dsdc_n988), 
	.B1(U_dsdc_n976), 
	.A(U_dsdc_n1546));
   NAND2_X1 U_dsdc_U883 (.ZN(U_dsdc_n641), 
	.A2(U_dsdc_n432), 
	.A1(U_dsdc_n196));
   AOI21_X1 U_dsdc_U882 (.ZN(U_dsdc_n1319), 
	.B2(U_dsdc_access_cs_3_), 
	.B1(U_dsdc_n1318), 
	.A(U_dsdc_n1317));
   NAND2_X2 U_dsdc_U881 (.ZN(U_dsdc_n1724), 
	.A2(U_dsdc_n1675), 
	.A1(U_dsdc_n1676));
   AOI22_X2 U_dsdc_U880 (.ZN(U_dsdc_n1889), 
	.B2(U_dsdc_n1890), 
	.B1(U_dsdc_n1907), 
	.A2(U_dsdc_n2082), 
	.A1(U_dsdc_bm_bank_status_3_));
   AOI21_X2 U_dsdc_U879 (.ZN(U_dsdc_n2048), 
	.B2(U_dsdc_n2014), 
	.B1(U_dsdc_n1977), 
	.A(U_dsdc_n2012));
   NOR2_X2 U_dsdc_U877 (.ZN(U_dsdc_n1411), 
	.A2(U_dsdc_n711), 
	.A1(U_dsdc_n692));
   OAI21_X2 U_dsdc_U875 (.ZN(U_dsdc_close_bank_addr_0_), 
	.B2(U_dsdc_n1127), 
	.B1(U_dsdc_n1391), 
	.A(U_dsdc_n1123));
   NAND2_X2 U_dsdc_U874 (.ZN(U_dsdc_n1712), 
	.A2(U_dsdc_n1715), 
	.A1(U_dsdc_n1708));
   NAND2_X2 U_dsdc_U873 (.ZN(U_dsdc_n1705), 
	.A2(U_dsdc_n1715), 
	.A1(U_dsdc_n1701));
   NOR2_X1 U_dsdc_U871 (.ZN(U_dsdc_n871), 
	.A2(U_dsdc_n170), 
	.A1(U_dsdc_n712));
   NAND2_X1 U_dsdc_U870 (.ZN(U_dsdc_n1650), 
	.A2(U_dsdc_n355), 
	.A1(U_dsdc_n871));
   NAND2_X2 U_dsdc_U869 (.ZN(U_dsdc_n789), 
	.A2(U_dsdc_bm_row_addr_1__11_), 
	.A1(U_dsdc_n604));
   NAND2_X2 U_dsdc_U868 (.ZN(U_dsdc_n782), 
	.A2(U_dsdc_bm_row_addr_1__15_), 
	.A1(U_dsdc_n604));
   NOR2_X1 U_dsdc_U867 (.ZN(U_dsdc_n1059), 
	.A2(U_dsdc_n935), 
	.A1(U_dsdc_n936));
   NAND3_X1 U_dsdc_U866 (.ZN(U_dsdc_n660), 
	.A3(U_dsdc_access_cs_1_), 
	.A2(U_dsdc_n167), 
	.A1(U_dsdc_n173));
   NAND2_X2 U_dsdc_U865 (.ZN(U_dsdc_n792), 
	.A2(U_dsdc_bm_row_addr_1__5_), 
	.A1(U_dsdc_n604));
   NAND2_X2 U_dsdc_U864 (.ZN(U_dsdc_n500), 
	.A2(U_dsdc_bm_row_addr_1__6_), 
	.A1(U_dsdc_n604));
   AOI22_X2 U_dsdc_U863 (.ZN(U_dsdc_n1919), 
	.B2(U_dsdc_n1920), 
	.B1(U_dsdc_n1937), 
	.A2(U_dsdc_n2082), 
	.A1(FE_PHN1593_U_dsdc_bm_bank_status_1_));
   AOI222_X1 U_dsdc_U862 (.ZN(U_dsdc_n752), 
	.C2(hiu_burst_size[1]), 
	.C1(U_dsdc_n983), 
	.B2(U_dsdc_r_burst_size_1_), 
	.B1(U_dsdc_n751), 
	.A2(U_dsdc_data_cnt_1_), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n85));
   NAND2_X2 U_dsdc_U861 (.ZN(U_dsdc_n1546), 
	.A2(U_dsdc_n1038), 
	.A1(U_dsdc_n670));
   INV_X4 U_dsdc_U860 (.ZN(U_dsdc_n601), 
	.A(U_dsdc_RSOP_1683_C2_CONTROL1));
   AOI22_X1 U_dsdc_U859 (.ZN(U_dsdc_n748), 
	.B2(FE_PHN1888_U_dsdc_r_burst_size_4_), 
	.B1(U_dsdc_n751), 
	.A2(U_dsdc_data_cnt_4_), 
	.A1(U_dsdc_RSOP_1683_C2_CONTROL1));
   NAND2_X2 U_dsdc_U858 (.ZN(U_dsdc_n1326), 
	.A2(U_dsdc_n1004), 
	.A1(U_dsdc_n1391));
   NAND2_X2 U_dsdc_U857 (.ZN(U_dsdc_n1391), 
	.A2(U_dsdc_n980), 
	.A1(U_dsdc_n981));
   NAND2_X1 U_dsdc_U855 (.ZN(U_dsdc_n1386), 
	.A2(U_dsdc_n991), 
	.A1(U_dsdc_n992));
   NAND2_X2 U_dsdc_U852 (.ZN(U_dsdc_n738), 
	.A2(U_dsdc_n1312), 
	.A1(U_dsdc_n936));
   NAND2_X1 U_dsdc_U851 (.ZN(U_dsdc_n933), 
	.A2(U_dsdc_n181), 
	.A1(U_dsdc_n1558));
   NAND2_X1 U_dsdc_U850 (.ZN(U_dsdc_n1651), 
	.A2(U_dsdc_n1558), 
	.A1(U_dsdc_n1410));
   NOR3_X1 U_dsdc_U849 (.ZN(U_dsdc_n1563), 
	.A3(U_dsdc_n1556), 
	.A2(U_dsdc_n1557), 
	.A1(U_dsdc_n1558));
   AOI211_X1 U_dsdc_U848 (.ZN(U_dsdc_n727), 
	.C2(U_dsdc_n724), 
	.C1(U_dsdc_n1558), 
	.B(U_dsdc_n722), 
	.A(U_dsdc_n723));
   NOR2_X1 U_dsdc_U847 (.ZN(U_dsdc_n1413), 
	.A2(U_dsdc_n165), 
	.A1(U_dsdc_n1558));
   AOI22_X2 U_dsdc_U846 (.ZN(U_dsdc_DP_OP_1642_126_2028_n4), 
	.B2(U_dsdc_DP_OP_1642_126_2028_n19), 
	.B1(U_dsdc_DP_OP_1642_126_2028_n60), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n14), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n5));
   AOI22_X2 U_dsdc_U845 (.ZN(U_dsdc_DP_OP_1642_126_2028_n6), 
	.B2(U_dsdc_DP_OP_1642_126_2028_n20), 
	.B1(U_dsdc_DP_OP_1642_126_2028_n59), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n15), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n7));
   AOI22_X2 U_dsdc_U844 (.ZN(U_dsdc_DP_OP_1642_126_2028_n2), 
	.B2(U_dsdc_DP_OP_1642_126_2028_n85), 
	.B1(U_dsdc_DP_OP_1642_126_2028_n61), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n3), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n13));
   XNOR2_X2 U_dsdc_U843 (.ZN(U_dsdc_n162), 
	.B(U_dsdc_DP_OP_1642_126_2028_n85), 
	.A(U_dsdc_DP_OP_1642_126_2028_n86));
   XNOR2_X2 U_dsdc_U842 (.ZN(U_dsdc_DP_OP_1642_126_2028_n11), 
	.B(U_dsdc_DP_OP_1642_126_2028_n85), 
	.A(U_dsdc_n162));
   INV_X2 U_dsdc_U841 (.ZN(U_dsdc_n1484), 
	.A(s_rd_ready));
   NAND2_X1 U_dsdc_U840 (.ZN(U_dsdc_n1156), 
	.A2(FE_PHN1158_U_dsdc_bm_ras_cnt_max_1_), 
	.A1(FE_PHN2034_U_dsdc_bm_ras_cnt_max_0_));
   NOR3_X2 U_dsdc_U839 (.ZN(U_dsdc_n1512), 
	.A3(U_dsdc_n432), 
	.A2(U_dsdc_operation_cs_2_), 
	.A1(U_dsdc_operation_cs_3_));
   NAND3_X2 U_dsdc_U836 (.ZN(U_dsdc_n692), 
	.A3(U_dsdc_access_cs_3_), 
	.A2(U_dsdc_n167), 
	.A1(U_dsdc_n298));
   NOR2_X2 U_dsdc_U834 (.ZN(U_dsdc_n1458), 
	.A2(U_dsdc_n170), 
	.A1(U_dsdc_n355));
   NOR2_X1 U_dsdc_U833 (.ZN(U_dsdc_n1568), 
	.A2(FE_PHN843_U_dsdc_num_init_ref_cnt_1_), 
	.A1(U_dsdc_num_init_ref_cnt_0_));
   NAND2_X1 U_dsdc_U832 (.ZN(U_dsdc_n739), 
	.A2(U_dsdc_data_flag), 
	.A1(U_dsdc_n306));
   OR2_X1 U_dsdc_U831 (.ZN(U_dsdc_n1644), 
	.A2(U_dsdc_term_cnt_2_), 
	.A1(U_dsdc_term_cnt_3_));
   OR4_X2 U_dsdc_U830 (.ZN(U_dsdc_n1446), 
	.A4(U_dsdc_cas_cnt_1_), 
	.A3(U_dsdc_cas_cnt_4_), 
	.A2(U_dsdc_cas_cnt_3_), 
	.A1(U_dsdc_cas_cnt_5_));
   NAND3_X2 U_dsdc_U829 (.ZN(U_dsdc_n712), 
	.A3(U_dsdc_access_cs_1_), 
	.A2(U_dsdc_access_cs_3_), 
	.A1(U_dsdc_n167));
   OR4_X2 U_dsdc_U828 (.ZN(U_dsdc_n1846), 
	.A4(U_dsdc_r_bm_close_bank_3_), 
	.A3(U_dsdc_r_bm_close_bank_1_), 
	.A2(U_dsdc_r_bm_close_bank_0_), 
	.A1(U_dsdc_r_bm_close_bank_2_));
   NAND2_X2 U_dsdc_U825 (.ZN(U_dsdc_n667), 
	.A2(U_dsdc_access_cs_2_), 
	.A1(U_dsdc_n170));
   NOR3_X2 U_dsdc_U824 (.ZN(U_dsdc_n1616), 
	.A3(U_dsdc_rcar_cnt2_0_), 
	.A2(U_dsdc_rcar_cnt2_1_), 
	.A1(U_dsdc_rcar_cnt2_2_));
   NAND2_X2 U_dsdc_U820 (.ZN(U_dsdc_n711), 
	.A2(U_dsdc_n170), 
	.A1(U_dsdc_n355));
   NAND2_X2 U_dsdc_U819 (.ZN(U_dsdc_n1522), 
	.A2(U_dsdc_operation_cs_0_), 
	.A1(U_dsdc_operation_cs_1_));
   OR4_X2 U_dsdc_U818 (.ZN(U_dsdc_n1776), 
	.A4(U_dsdc_row_cnt_3_), 
	.A3(U_dsdc_row_cnt_2_), 
	.A2(U_dsdc_row_cnt_1_), 
	.A1(U_dsdc_row_cnt_0_));
   NAND3_X2 U_dsdc_U815 (.ZN(U_dsdc_n1485), 
	.A3(U_dsdc_n432), 
	.A2(U_dsdc_operation_cs_2_), 
	.A1(U_dsdc_operation_cs_3_));
   NAND2_X2 U_dsdc_U814 (.ZN(U_dsdc_n1490), 
	.A2(U_dsdc_n344), 
	.A1(U_dsdc_n343));
   NOR2_X2 U_dsdc_U813 (.ZN(U_dsdc_n1435), 
	.A2(U_dsdc_n344), 
	.A1(U_dsdc_operation_cs_1_));
   NAND2_X2 U_dsdc_U812 (.ZN(U_dsdc_n1455), 
	.A2(U_dsdc_n344), 
	.A1(U_dsdc_operation_cs_1_));
   NAND3_X2 U_dsdc_U811 (.ZN(U_dsdc_n1451), 
	.A3(U_dsdc_n341), 
	.A2(U_dsdc_n432), 
	.A1(U_dsdc_operation_cs_3_));
   XNOR2_X1 U_dsdc_U810 (.ZN(U_dsdc_n1305), 
	.B(U_dsdc_wr_cnt_0_), 
	.A(U_dsdc_n195));
   AND2_X2 U_dsdc_U808 (.ZN(U_dsdc_n308), 
	.A2(U_dsdc_bm_bank_age_0__2_), 
	.A1(U_dsdc_n1842));
   INV_X1 U_dsdc_U807 (.ZN(U_dsdc_n1585), 
	.A(U_dsdc_n1583));
   INV_X1 U_dsdc_U806 (.ZN(U_dsdc_n1190), 
	.A(U_dsdc_n1189));
   OAI21_X1 U_dsdc_U805 (.ZN(U_dsdc_n1330), 
	.B2(U_dsdc_n309), 
	.B1(U_dsdc_n171), 
	.A(U_dsdc_n1329));
   INV_X2 U_dsdc_U804 (.ZN(U_dsdc_n1431), 
	.A(U_dsdc_n1509));
   INV_X1 U_dsdc_U802 (.ZN(U_dsdc_n1158), 
	.A(U_dsdc_n1153));
   INV_X1 U_dsdc_U801 (.ZN(U_dsdc_n1197), 
	.A(FE_PHN1154_U_dsdc_n1196));
   INV_X2 U_dsdc_U800 (.ZN(U_dsdc_n642), 
	.A(U_dsdc_n1522));
   INV_X1 U_dsdc_U799 (.ZN(U_dsdc_n1743), 
	.A(U_dsdc_n1747));
   INV_X2 U_dsdc_U798 (.ZN(U_dsdc_n476), 
	.A(U_dsdc_n1841));
   NAND2_X1 U_dsdc_U797 (.ZN(U_dsdc_n1460), 
	.A2(s_cas_latency[1]), 
	.A1(FE_PHN787_n90));
   OR4_X2 U_dsdc_U796 (.ZN(U_dsdc_n357), 
	.A4(U_cr_n70), 
	.A3(U_cr_n42), 
	.A2(cr_row_addr_width[0]), 
	.A1(FE_PHN3054_cr_row_addr_width_2_));
   INV_X1 U_dsdc_U795 (.ZN(U_dsdc_n657), 
	.A(U_dsdc_n692));
   NAND3_X1 U_dsdc_U794 (.ZN(U_dsdc_n688), 
	.A3(U_dsdc_n301), 
	.A2(U_dsdc_n172), 
	.A1(U_dsdc_n687));
   INV_X2 U_dsdc_U793 (.ZN(U_dsdc_n661), 
	.A(U_dsdc_n1455));
   INV_X1 U_dsdc_U792 (.ZN(U_dsdc_n1711), 
	.A(U_dsdc_n1719));
   INV_X1 U_dsdc_U791 (.ZN(U_dsdc_n1211), 
	.A(FE_PHN1155_U_dsdc_n1210));
   INV_X1 U_dsdc_U790 (.ZN(U_dsdc_n645), 
	.A(U_dsdc_n1490));
   NOR2_X2 U_dsdc_U789 (.ZN(U_dsdc_n1427), 
	.A2(U_dsdc_access_cs_1_), 
	.A1(U_dsdc_n649));
   INV_X1 U_dsdc_U788 (.ZN(U_dsdc_n1087), 
	.A(U_dsdc_n1082));
   NAND2_X1 U_dsdc_U787 (.ZN(U_dsdc_n1641), 
	.A2(FE_PHN671_U_dsdc_n1637), 
	.A1(U_dsdc_n1638));
   INV_X1 U_dsdc_U786 (.ZN(U_dsdc_n1204), 
	.A(U_dsdc_n1203));
   INV_X2 U_dsdc_U785 (.ZN(U_dsdc_n1632), 
	.A(U_dsdc_n1419));
   INV_X1 U_dsdc_U784 (.ZN(U_dsdc_n915), 
	.A(U_dsdc_n712));
   INV_X1 U_dsdc_U783 (.ZN(U_dsdc_n652), 
	.A(U_dsdc_n711));
   INV_X2 U_dsdc_U782 (.ZN(U_dsdc_n658), 
	.A(U_dsdc_n1458));
   INV_X1 U_dsdc_U781 (.ZN(U_dsdc_n654), 
	.A(U_dsdc_n660));
   INV_X2 U_dsdc_U780 (.ZN(U_dsdc_n1465), 
	.A(FE_PHN2909_U_dsdc_n1436));
   INV_X1 U_dsdc_U779 (.ZN(U_dsdc_n1176), 
	.A(FE_PHN945_U_dsdc_n1175));
   INV_X1 U_dsdc_U778 (.ZN(U_dsdc_n1229), 
	.A(U_dsdc_n1228));
   INV_X2 U_dsdc_U777 (.ZN(U_dsdc_n1605), 
	.A(U_dsdc_n1604));
   NAND2_X1 U_dsdc_U776 (.ZN(U_dsdc_n1658), 
	.A2(U_cr_n21), 
	.A1(cr_row_addr_width[1]));
   OR3_X2 U_dsdc_U775 (.ZN(U_dsdc_n1770), 
	.A3(U_dsdc_n1776), 
	.A2(U_dsdc_row_cnt_4_), 
	.A1(U_dsdc_row_cnt_5_));
   INV_X1 U_dsdc_U774 (.ZN(U_dsdc_n1487), 
	.A(U_dsdc_n1485));
   INV_X2 U_dsdc_U773 (.ZN(U_dsdc_n1652), 
	.A(U_dsdc_n1662));
   OR4_X2 U_dsdc_U772 (.ZN(U_dsdc_n358), 
	.A4(U_cr_n70), 
	.A3(FE_PHN3054_cr_row_addr_width_2_), 
	.A2(cr_row_addr_width[0]), 
	.A1(cr_row_addr_width[1]));
   INV_X1 U_dsdc_U771 (.ZN(U_dsdc_n1239), 
	.A(FE_PHN1497_U_dsdc_n1238));
   NOR2_X1 U_dsdc_U770 (.ZN(U_dsdc_n714), 
	.A2(n84), 
	.A1(U_dsdc_n1040));
   NAND2_X1 U_dsdc_U769 (.ZN(U_dsdc_n1659), 
	.A2(U_cr_n42), 
	.A1(cr_row_addr_width[0]));
   INV_X1 U_dsdc_U768 (.ZN(U_dsdc_n1183), 
	.A(FE_PHN1156_U_dsdc_n1182));
   OAI22_X1 U_dsdc_U767 (.ZN(U_dsdc_n1162), 
	.B2(U_dsdc_n174), 
	.B1(U_dsdc_n326), 
	.A2(U_dsdc_n1165), 
	.A1(U_dsdc_n1163));
   NOR2_X1 U_dsdc_U765 (.ZN(U_dsdc_n1245), 
	.A2(FE_PHN1333_U_dsdc_n382), 
	.A1(U_dsdc_n1244));
   NOR2_X1 U_dsdc_U764 (.ZN(U_dsdc_n1187), 
	.A2(FE_PHN1337_U_dsdc_n363), 
	.A1(U_dsdc_n1186));
   OAI21_X1 U_dsdc_U760 (.ZN(U_dsdc_n1832), 
	.B2(U_dsdc_n304), 
	.B1(U_dsdc_n1841), 
	.A(U_dsdc_n1831));
   OAI21_X1 U_dsdc_U759 (.ZN(U_dsdc_n1830), 
	.B2(U_dsdc_n302), 
	.B1(U_dsdc_n1841), 
	.A(U_dsdc_n1829));
   AOI21_X1 U_dsdc_U758 (.ZN(U_dsdc_n1508), 
	.B2(U_dsdc_n1506), 
	.B1(U_dsdc_operation_cs_2_), 
	.A(U_dsdc_operation_cs_3_));
   INV_X1 U_dsdc_U757 (.ZN(U_dsdc_n662), 
	.A(U_dsdc_n1454));
   INV_X1 U_dsdc_U756 (.ZN(U_dsdc_n1956), 
	.A(U_dsdc_n1961));
   INV_X1 U_dsdc_U755 (.ZN(U_dsdc_n1037), 
	.A(U_dsdc_n1284));
   NOR2_X1 U_dsdc_U754 (.ZN(U_dsdc_n1164), 
	.A2(U_dsdc_rcd_cnt_0_), 
	.A1(U_dsdc_n1163));
   XNOR2_X1 U_dsdc_U753 (.ZN(U_dsdc_n1088), 
	.B(s_cas_latency[2]), 
	.A(U_dsdc_n1460));
   INV_X2 U_dsdc_U752 (.ZN(U_dsdc_n1461), 
	.A(FE_PHN894_U_dsdc_n1464));
   NAND2_X1 U_dsdc_U751 (.ZN(U_dsdc_n1081), 
	.A2(s_cas_latency[2]), 
	.A1(U_dsdc_n1460));
   INV_X2 U_dsdc_U750 (.ZN(U_dsdc_n1452), 
	.A(U_dsdc_n1536));
   NAND2_X2 U_dsdc_U749 (.ZN(U_dsdc_n1558), 
	.A2(FE_PHN1035_U_dsdc_n327), 
	.A1(U_dsdc_n663));
   INV_X1 U_dsdc_U747 (.ZN(U_dsdc_n1420), 
	.A(U_dsdc_n1633));
   NAND2_X2 U_dsdc_U746 (.ZN(U_dsdc_n966), 
	.A2(U_dsdc_access_cs_0_), 
	.A1(U_dsdc_n1427));
   NOR2_X1 U_dsdc_U745 (.ZN(U_dsdc_n612), 
	.A2(U_dsdc_N4239), 
	.A1(U_dsdc_N4240));
   NOR2_X1 U_dsdc_U744 (.ZN(U_dsdc_n1215), 
	.A2(FE_PHN1334_U_dsdc_n365), 
	.A1(U_dsdc_n1214));
   AOI21_X1 U_dsdc_U743 (.ZN(U_dsdc_n1586), 
	.B2(U_dsdc_n1585), 
	.B1(U_dsdc_rcar_cnt1_2_), 
	.A(U_dsdc_n1584));
   NOR2_X1 U_dsdc_U742 (.ZN(U_dsdc_n1201), 
	.A2(FE_PHN1336_U_dsdc_n364), 
	.A1(U_dsdc_n1200));
   NAND2_X1 U_dsdc_U741 (.ZN(U_dsdc_n1589), 
	.A2(U_dsdc_n1587), 
	.A1(U_dsdc_rcar_cnt1_3_));
   OR3_X2 U_dsdc_U740 (.ZN(U_dsdc_n1765), 
	.A3(U_dsdc_n1770), 
	.A2(U_dsdc_row_cnt_6_), 
	.A1(U_dsdc_row_cnt_7_));
   INV_X1 U_dsdc_U739 (.ZN(U_dsdc_n1348), 
	.A(U_dsdc_n1427));
   INV_X1 U_dsdc_U738 (.ZN(U_dsdc_n1360), 
	.A(U_dsdc_n1426));
   NAND2_X1 U_dsdc_U737 (.ZN(U_dsdc_n1628), 
	.A2(U_dsdc_r_rw), 
	.A1(U_dsdc_n1425));
   INV_X2 U_dsdc_U736 (.ZN(U_dsdc_n710), 
	.A(U_dsdc_n1418));
   NAND2_X1 U_dsdc_U735 (.ZN(U_dsdc_n1531), 
	.A2(U_dsdc_n343), 
	.A1(U_dsdc_n1434));
   INV_X2 U_dsdc_U734 (.ZN(U_dsdc_n1300), 
	.A(U_dsdc_n1312));
   OAI21_X1 U_dsdc_U733 (.ZN(U_dsdc_n1357), 
	.B2(U_dsdc_n667), 
	.B1(U_dsdc_n692), 
	.A(U_dsdc_n653));
   INV_X2 U_dsdc_U732 (.ZN(U_dsdc_n1152), 
	.A(U_dsdc_n1437));
   NAND2_X1 U_dsdc_U731 (.ZN(U_dsdc_n937), 
	.A2(U_dsdc_n1415), 
	.A1(U_dsdc_n904));
   NAND2_X1 U_dsdc_U729 (.ZN(U_dsdc_n828), 
	.A2(U_dsdc_n940), 
	.A1(U_dsdc_n988));
   NAND2_X1 U_dsdc_U728 (.ZN(U_dsdc_n674), 
	.A2(U_dsdc_n1412), 
	.A1(U_dsdc_n904));
   NOR2_X1 U_dsdc_U727 (.ZN(U_dsdc_n1365), 
	.A2(U_dsdc_n1803), 
	.A1(U_dsdc_n1362));
   OR3_X2 U_dsdc_U726 (.ZN(U_dsdc_n1795), 
	.A3(U_dsdc_n1765), 
	.A2(U_dsdc_row_cnt_8_), 
	.A1(U_dsdc_row_cnt_9_));
   INV_X2 U_dsdc_U725 (.ZN(U_dsdc_n668), 
	.A(U_dsdc_n904));
   NAND2_X1 U_dsdc_U724 (.ZN(U_dsdc_n868), 
	.A2(U_dsdc_n866), 
	.A1(U_dsdc_n867));
   INV_X1 U_dsdc_U723 (.ZN(U_dsdc_n659), 
	.A(U_dsdc_n1292));
   NAND2_X1 U_dsdc_U722 (.ZN(U_dsdc_n852), 
	.A2(U_dsdc_n1384), 
	.A1(U_dsdc_n1362));
   NAND2_X1 U_dsdc_U721 (.ZN(U_dsdc_n648), 
	.A2(U_dsdc_n1577), 
	.A1(U_dsdc_n1564));
   INV_X2 U_dsdc_U720 (.ZN(U_dsdc_n643), 
	.A(U_dsdc_n1432));
   OAI21_X2 U_dsdc_U719 (.ZN(U_dsdc_n1754), 
	.B2(cr_do_self_ref_rp), 
	.B1(U_dsdc_n1532), 
	.A(U_dsdc_n1497));
   INV_X2 U_dsdc_U718 (.ZN(U_dsdc_n684), 
	.A(U_dsdc_n1424));
   INV_X2 U_dsdc_U717 (.ZN(U_dsdc_n1438), 
	.A(hiu_rw));
   INV_X2 U_dsdc_U716 (.ZN(U_dsdc_n736), 
	.A(U_dsdc_n741));
   INV_X2 U_dsdc_U715 (.ZN(U_dsdc_n1524), 
	.A(U_dsdc_n1510));
   INV_X2 U_dsdc_U714 (.ZN(U_dsdc_n1079), 
	.A(U_dsdc_n1414));
   INV_X1 U_dsdc_U713 (.ZN(U_dsdc_n1471), 
	.A(U_dsdc_n1479));
   NAND2_X1 U_dsdc_U712 (.ZN(U_dsdc_n1469), 
	.A2(FE_PHN2909_U_dsdc_n1436), 
	.A1(U_dsdc_n1428));
   INV_X4 U_dsdc_U711 (.ZN(U_dsdc_n703), 
	.A(U_dsdc_n1558));
   NAND2_X1 U_dsdc_U710 (.ZN(U_dsdc_n735), 
	.A2(U_cr_n58), 
	.A1(U_dsdc_n1414));
   INV_X2 U_dsdc_U709 (.ZN(U_dsdc_n1631), 
	.A(U_dsdc_n1628));
   INV_X2 U_dsdc_U708 (.ZN(U_dsdc_n1470), 
	.A(U_dsdc_n1499));
   INV_X2 U_dsdc_U704 (.ZN(U_dsdc_n837), 
	.A(U_dsdc_n1195));
   INV_X2 U_dsdc_U703 (.ZN(U_dsdc_n838), 
	.A(U_dsdc_n1181));
   INV_X2 U_dsdc_U702 (.ZN(U_dsdc_n841), 
	.A(U_dsdc_n1237));
   INV_X2 U_dsdc_U701 (.ZN(U_dsdc_n842), 
	.A(U_dsdc_n1209));
   NAND3_X1 U_dsdc_U700 (.ZN(U_dsdc_n1901), 
	.A3(U_dsdc_n1906), 
	.A2(U_dsdc_bm_bank_age_3__0_), 
	.A1(U_dsdc_bm_bank_age_3__1_));
   XNOR2_X1 U_dsdc_U698 (.ZN(U_dsdc_add_x_2600_1_n8), 
	.B(FE_PHN5064_s_read_pipe_0_), 
	.A(U_dsdc_n1088));
   INV_X2 U_dsdc_U697 (.ZN(U_dsdc_n751), 
	.A(U_dsdc_n1258));
   NAND2_X1 U_dsdc_U696 (.ZN(U_dsdc_n1447), 
	.A2(U_dsdc_n1437), 
	.A1(debug_ref_req));
   NAND2_X1 U_dsdc_U695 (.ZN(U_dsdc_n1959), 
	.A2(U_dsdc_n1972), 
	.A1(U_dsdc_bm_bank_age_0__0_));
   INV_X2 U_dsdc_U693 (.ZN(U_dsdc_n1061), 
	.A(U_dsdc_n903));
   NAND2_X1 U_dsdc_U692 (.ZN(U_dsdc_n856), 
	.A2(U_cr_n58), 
	.A1(U_dsdc_n1437));
   NOR2_X1 U_dsdc_U691 (.ZN(U_dsdc_n1115), 
	.A2(U_dsdc_n450), 
	.A1(U_dsdc_n1136));
   INV_X2 U_dsdc_U689 (.ZN(U_dsdc_n1109), 
	.A(U_dsdc_n1136));
   NOR2_X1 U_dsdc_U687 (.ZN(U_dsdc_n1132), 
	.A2(U_dsdc_n454), 
	.A1(U_dsdc_n1136));
   NOR2_X1 U_dsdc_U686 (.ZN(U_dsdc_n1134), 
	.A2(U_dsdc_n455), 
	.A1(U_dsdc_n1136));
   NOR2_X1 U_dsdc_U685 (.ZN(U_dsdc_n1137), 
	.A2(U_dsdc_n456), 
	.A1(U_dsdc_n1136));
   NAND2_X1 U_dsdc_U683 (.ZN(U_dsdc_n1044), 
	.A2(U_dsdc_n1413), 
	.A1(U_dsdc_n1410));
   NOR2_X1 U_dsdc_U682 (.ZN(U_dsdc_n1116), 
	.A2(U_dsdc_n451), 
	.A1(U_dsdc_n1136));
   XNOR2_X1 U_dsdc_U681 (.ZN(U_dsdc_n1091), 
	.B(s_read_pipe[2]), 
	.A(FE_PHN893_U_dsdc_n1092));
   INV_X1 U_dsdc_U680 (.ZN(U_dsdc_n1263), 
	.A(hiu_burst_size[2]));
   NAND2_X1 U_dsdc_U678 (.ZN(U_dsdc_n478), 
	.A2(U_dsdc_n334), 
	.A1(U_dsdc_n477));
   AOI21_X1 U_dsdc_U677 (.ZN(U_dsdc_n1946), 
	.B2(U_dsdc_bm_bank_age_0__1_), 
	.B1(U_dsdc_n1944), 
	.A(U_dsdc_bm_bank_age_0__0_));
   NOR2_X1 U_dsdc_U676 (.ZN(U_dsdc_n1913), 
	.A2(U_dsdc_n1953), 
	.A1(U_dsdc_bm_bank_age_1__3_));
   NOR2_X1 U_dsdc_U673 (.ZN(U_dsdc_n1117), 
	.A2(U_dsdc_n452), 
	.A1(U_dsdc_n1136));
   NOR2_X1 U_dsdc_U672 (.ZN(U_dsdc_n1122), 
	.A2(U_dsdc_n453), 
	.A1(U_dsdc_n1136));
   OAI21_X1 U_dsdc_U671 (.ZN(U_dsdc_n1892), 
	.B2(U_dsdc_n1900), 
	.B1(U_dsdc_n304), 
	.A(U_dsdc_n302));
   NOR2_X1 U_dsdc_U670 (.ZN(U_dsdc_n1883), 
	.A2(U_dsdc_n1953), 
	.A1(U_dsdc_bm_bank_age_3__3_));
   OAI21_X1 U_dsdc_U669 (.ZN(U_dsdc_n1852), 
	.B2(FE_PHN958_U_dsdc_n353), 
	.B1(U_dsdc_n1860), 
	.A(U_dsdc_n178));
   INV_X1 U_dsdc_U668 (.ZN(U_dsdc_n1729), 
	.A(FE_PHN969_U_dsdc_n1727));
   NAND2_X1 U_dsdc_U667 (.ZN(U_dsdc_n1726), 
	.A2(U_dsdc_n1754), 
	.A1(cr_t_xsr[8]));
   NOR2_X1 U_dsdc_U666 (.ZN(U_dsdc_n1538), 
	.A2(U_dsdc_n1537), 
	.A1(n84));
   OAI21_X1 U_dsdc_U665 (.ZN(U_dsdc_n1824), 
	.B2(U_dsdc_n436), 
	.B1(U_dsdc_n1825), 
	.A(FE_PHN773_U_dsdc_n1823));
   NAND2_X1 U_dsdc_U664 (.ZN(U_dsdc_n1385), 
	.A2(U_dsdc_n865), 
	.A1(U_dsdc_n1496));
   INV_X2 U_dsdc_U663 (.ZN(U_dsdc_n2069), 
	.A(U_dsdc_n1416));
   OR4_X2 U_dsdc_U661 (.ZN(U_dsdc_n1448), 
	.A4(hiu_burst_size[1]), 
	.A3(hiu_burst_size[2]), 
	.A2(hiu_burst_size[3]), 
	.A1(hiu_burst_size[5]));
   INV_X2 U_dsdc_U660 (.ZN(U_dsdc_n1511), 
	.A(U_dsdc_n2058));
   INV_X2 U_dsdc_U658 (.ZN(U_dsdc_n721), 
	.A(U_dsdc_n1805));
   NAND2_X1 U_dsdc_U657 (.ZN(U_dsdc_n737), 
	.A2(U_dsdc_n1419), 
	.A1(U_dsdc_n736));
   AND2_X2 U_dsdc_U656 (.ZN(U_dsdc_n362), 
	.A2(U_dsdc_n1433), 
	.A1(U_dsdc_n648));
   INV_X1 U_dsdc_U655 (.ZN(U_dsdc_n761), 
	.A(U_dsdc_n1876));
   INV_X1 U_dsdc_U654 (.ZN(U_dsdc_n1253), 
	.A(hiu_burst_size[0]));
   NOR2_X1 U_dsdc_U653 (.ZN(U_dsdc_n1069), 
	.A2(U_dsdc_n447), 
	.A1(U_dsdc_n1136));
   INV_X2 U_dsdc_U652 (.ZN(U_dsdc_n644), 
	.A(U_dsdc_n648));
   INV_X2 U_dsdc_U651 (.ZN(U_dsdc_n723), 
	.A(U_dsdc_n1315));
   INV_X2 U_dsdc_U650 (.ZN(U_dsdc_n1634), 
	.A(U_dsdc_n1648));
   NOR2_X1 U_dsdc_U648 (.ZN(U_dsdc_n1073), 
	.A2(U_dsdc_n448), 
	.A1(U_dsdc_n1136));
   INV_X2 U_dsdc_U646 (.ZN(U_dsdc_n675), 
	.A(U_dsdc_n881));
   NAND2_X1 U_dsdc_U645 (.ZN(U_dsdc_n1353), 
	.A2(U_dsdc_n1483), 
	.A1(U_dsdc_n1496));
   INV_X2 U_dsdc_U644 (.ZN(U_dsdc_n682), 
	.A(U_dsdc_n879));
   INV_X1 U_dsdc_U643 (.ZN(U_dsdc_n1361), 
	.A(U_dsdc_n1357));
   NOR2_X1 U_dsdc_U642 (.ZN(U_dsdc_n1095), 
	.A2(U_dsdc_n449), 
	.A1(U_dsdc_n1136));
   OR3_X2 U_dsdc_U641 (.ZN(U_dsdc_n1794), 
	.A3(U_dsdc_n1795), 
	.A2(U_dsdc_row_cnt_10_), 
	.A1(U_dsdc_row_cnt_11_));
   INV_X1 U_dsdc_U640 (.ZN(U_dsdc_n1259), 
	.A(U_dsdc_n1269));
   NOR2_X1 U_dsdc_U639 (.ZN(U_dsdc_n935), 
	.A2(U_dsdc_n933), 
	.A1(U_dsdc_n934));
   INV_X2 U_dsdc_U638 (.ZN(U_dsdc_n1592), 
	.A(U_dsdc_n852));
   NAND2_X1 U_dsdc_U637 (.ZN(U_dsdc_n1746), 
	.A2(U_dsdc_n1754), 
	.A1(cr_t_xsr[3]));
   INV_X2 U_dsdc_U636 (.ZN(U_dsdc_n1866), 
	.A(U_dsdc_n1860));
   NAND2_X1 U_dsdc_U635 (.ZN(U_dsdc_n1755), 
	.A2(U_dsdc_n1754), 
	.A1(cr_t_xsr[0]));
   INV_X2 U_dsdc_U634 (.ZN(U_dsdc_n1654), 
	.A(U_dsdc_n1656));
   NAND2_X1 U_dsdc_U633 (.ZN(U_dsdc_n1753), 
	.A2(U_dsdc_n1754), 
	.A1(FE_PHN4714_cr_t_xsr_1_));
   AOI21_X1 U_dsdc_U631 (.ZN(U_dsdc_n733), 
	.B2(U_dsdc_n440), 
	.B1(U_dsdc_n1805), 
	.A(U_dsdc_early_term_flag));
   AOI22_X1 U_dsdc_U630 (.ZN(U_dsdc_n1566), 
	.B2(cr_num_init_ref[0]), 
	.B1(U_dsdc_n1667), 
	.A2(U_dsdc_num_init_ref_cnt_0_), 
	.A1(U_dsdc_n1565));
   NAND2_X1 U_dsdc_U629 (.ZN(U_dsdc_n1575), 
	.A2(U_dsdc_n1574), 
	.A1(U_dsdc_n2051));
   OAI211_X1 U_dsdc_U628 (.ZN(U_dsdc_n1569), 
	.C2(U_dsdc_n2063), 
	.C1(U_dsdc_num_init_ref_cnt_0_), 
	.B(FE_PHN843_U_dsdc_num_init_ref_cnt_1_), 
	.A(U_dsdc_n1433));
   NAND2_X1 U_dsdc_U627 (.ZN(U_dsdc_n1570), 
	.A2(cr_num_init_ref[1]), 
	.A1(U_dsdc_n1667));
   NAND3_X1 U_dsdc_U626 (.ZN(U_dsdc_n1295), 
	.A3(U_dsdc_n1650), 
	.A2(U_dsdc_n2014), 
	.A1(U_dsdc_n1292));
   NAND2_X1 U_dsdc_U624 (.ZN(U_dsdc_n1837), 
	.A2(U_dsdc_n1911), 
	.A1(U_dsdc_bm_bank_age_2__2_));
   NOR2_X1 U_dsdc_U623 (.ZN(U_dsdc_n1474), 
	.A2(U_dsdc_n1483), 
	.A1(U_dsdc_n2014));
   OAI21_X1 U_dsdc_U622 (.ZN(U_dsdc_n993), 
	.B2(U_dsdc_n1650), 
	.B1(U_dsdc_n1496), 
	.A(U_dsdc_n1342));
   NAND2_X1 U_dsdc_U621 (.ZN(U_dsdc_n1476), 
	.A2(U_dsdc_n1728), 
	.A1(U_dsdc_n1430));
   NOR2_X1 U_dsdc_U619 (.ZN(U_dsdc_n836), 
	.A2(U_dsdc_n1353), 
	.A1(U_dsdc_n988));
   NAND2_X1 U_dsdc_U617 (.ZN(U_dsdc_n2078), 
	.A2(U_dsdc_n1397), 
	.A1(U_dsdc_n165));
   NAND2_X1 U_dsdc_U616 (.ZN(U_dsdc_n651), 
	.A2(U_dsdc_n1425), 
	.A1(U_dsdc_n1423));
   NOR2_X2 U_dsdc_U614 (.ZN(U_dsdc_n1478), 
	.A2(U_dsdc_n597), 
	.A1(U_dsdc_n1794));
   NAND3_X1 U_dsdc_U613 (.ZN(U_dsdc_n1350), 
	.A3(U_dsdc_n868), 
	.A2(U_dsdc_n869), 
	.A1(U_dsdc_n1385));
   NAND2_X1 U_dsdc_U610 (.ZN(U_dsdc_n1313), 
	.A2(U_dsdc_n1060), 
	.A1(U_dsdc_n879));
   NOR3_X1 U_dsdc_U608 (.ZN(U_dsdc_wrapped_pop_flag_nxt), 
	.A3(U_dsdc_n181), 
	.A2(U_dsdc_n1651), 
	.A1(cr_delayed_precharge));
   NOR2_X1 U_dsdc_U607 (.ZN(U_dsdc_n1730), 
	.A2(U_dsdc_n1754), 
	.A1(U_dsdc_n1729));
   OAI21_X1 U_dsdc_U606 (.ZN(U_dsdc_n1732), 
	.B2(U_dsdc_n1736), 
	.B1(FE_PHN816_U_dsdc_n359), 
	.A(U_dsdc_n1733));
   NAND2_X1 U_dsdc_U605 (.ZN(U_dsdc_n1915), 
	.A2(U_dsdc_n1911), 
	.A1(U_dsdc_bm_bank_age_1__2_));
   INV_X2 U_dsdc_U604 (.ZN(U_dsdc_n1951), 
	.A(U_dsdc_n1911));
   INV_X2 U_dsdc_U603 (.ZN(U_dsdc_n479), 
	.A(U_dsdc_n1946));
   NAND2_X1 U_dsdc_U602 (.ZN(U_dsdc_n1674), 
	.A2(U_dsdc_n1722), 
	.A1(cr_t_init[15]));
   INV_X2 U_dsdc_U601 (.ZN(U_dsdc_n1948), 
	.A(U_dsdc_n1943));
   NAND3_X1 U_dsdc_U600 (.ZN(U_dsdc_n1939), 
	.A3(U_dsdc_bm_bank_age_1__3_), 
	.A2(U_dsdc_n1938), 
	.A1(U_dsdc_n349));
   NAND2_X1 U_dsdc_U599 (.ZN(U_dsdc_n1693), 
	.A2(U_dsdc_n1722), 
	.A1(cr_t_init[9]));
   INV_X1 U_dsdc_U598 (.ZN(U_dsdc_n1567), 
	.A(U_dsdc_n1580));
   NAND2_X1 U_dsdc_U597 (.ZN(U_dsdc_n1700), 
	.A2(U_dsdc_n1722), 
	.A1(cr_t_init[7]));
   NAND2_X1 U_dsdc_U596 (.ZN(U_dsdc_n1707), 
	.A2(U_dsdc_n1722), 
	.A1(cr_t_init[5]));
   NAND2_X1 U_dsdc_U595 (.ZN(U_dsdc_n1714), 
	.A2(U_dsdc_n1722), 
	.A1(cr_t_init[3]));
   OR3_X2 U_dsdc_U594 (.ZN(U_dsdc_n1788), 
	.A3(U_dsdc_n1794), 
	.A2(U_dsdc_row_cnt_12_), 
	.A1(U_dsdc_row_cnt_13_));
   NOR2_X1 U_dsdc_U593 (.ZN(U_dsdc_n1571), 
	.A2(U_dsdc_n2051), 
	.A1(U_dsdc_n1666));
   INV_X2 U_dsdc_U592 (.ZN(U_dsdc_n1621), 
	.A(U_dsdc_n1535));
   OAI211_X1 U_dsdc_U591 (.ZN(U_dsdc_n2055), 
	.C2(U_dsdc_n1532), 
	.C1(U_cr_n39), 
	.B(U_dsdc_n1531), 
	.A(U_dsdc_n1535));
   OAI211_X1 U_dsdc_U590 (.ZN(U_dsdc_n1725), 
	.C2(FE_PHN969_U_dsdc_n1727), 
	.C1(U_dsdc_xsr_cnt_7_), 
	.B(U_dsdc_n1733), 
	.A(U_dsdc_xsr_cnt_8_));
   NAND2_X1 U_dsdc_U589 (.ZN(U_dsdc_n1885), 
	.A2(U_dsdc_n1911), 
	.A1(U_dsdc_bm_bank_age_3__2_));
   INV_X2 U_dsdc_U585 (.ZN(U_dsdc_n585), 
	.A(U_dsdc_n1788));
   INV_X4 U_dsdc_U581 (.ZN(U_dsdc_n1344), 
	.A(U_dsdc_n991));
   OAI211_X1 U_dsdc_U580 (.ZN(U_dsdc_n1745), 
	.C2(U_dsdc_n1743), 
	.C1(U_dsdc_xsr_cnt_2_), 
	.B(U_dsdc_n1750), 
	.A(FE_PHN1030_U_dsdc_xsr_cnt_3_));
   INV_X2 U_dsdc_U579 (.ZN(U_dsdc_n1619), 
	.A(U_dsdc_n1617));
   INV_X2 U_dsdc_U577 (.ZN(U_dsdc_n1502), 
	.A(U_dsdc_n1500));
   AOI22_X1 U_dsdc_U576 (.ZN(U_dsdc_n1731), 
	.B2(U_dsdc_n1754), 
	.B1(cr_t_xsr[7]), 
	.A2(U_dsdc_n1730), 
	.A1(U_dsdc_xsr_cnt_7_));
   OAI21_X1 U_dsdc_U574 (.ZN(U_dsdc_n1735), 
	.B2(U_dsdc_n1733), 
	.B1(cr_t_xsr[6]), 
	.A(U_dsdc_n1732));
   OAI211_X1 U_dsdc_U573 (.ZN(U_dsdc_n1738), 
	.C2(U_dsdc_n1737), 
	.C1(U_dsdc_xsr_cnt_4_), 
	.B(U_dsdc_n1750), 
	.A(U_dsdc_xsr_cnt_5_));
   INV_X2 U_dsdc_U572 (.ZN(U_dsdc_n1756), 
	.A(U_dsdc_n1750));
   NAND3_X1 U_dsdc_U571 (.ZN(U_dsdc_n1752), 
	.A3(U_dsdc_n1750), 
	.A2(FE_PHN1033_U_dsdc_xsr_cnt_1_), 
	.A1(U_dsdc_xsr_cnt_0_));
   NAND3_X1 U_dsdc_U570 (.ZN(U_dsdc_n1323), 
	.A3(U_dsdc_n1329), 
	.A2(U_dsdc_rp_cnt2_2_), 
	.A1(U_dsdc_n1335));
   INV_X2 U_dsdc_U568 (.ZN(U_dsdc_n669), 
	.A(U_dsdc_n760));
   INV_X2 U_dsdc_U567 (.ZN(U_dsdc_n1062), 
	.A(U_dsdc_n1059));
   NOR2_X1 U_dsdc_U565 (.ZN(U_dsdc_n1351), 
	.A2(U_dsdc_n1349), 
	.A1(U_dsdc_n1350));
   OAI211_X1 U_dsdc_U562 (.ZN(U_dsdc_n1363), 
	.C2(U_dsdc_n165), 
	.C1(U_dsdc_n1627), 
	.B(U_dsdc_n1342), 
	.A(U_dsdc_n1343));
   NAND2_X1 U_dsdc_U559 (.ZN(U_dsdc_n939), 
	.A2(debug_ref_req), 
	.A1(U_dsdc_n1038));
   OAI21_X1 U_dsdc_U558 (.ZN(U_dsdc_n1821), 
	.B2(U_dsdc_n437), 
	.B1(U_dsdc_n1822), 
	.A(U_dsdc_n1820));
   INV_X2 U_dsdc_U557 (.ZN(U_dsdc_n1031), 
	.A(U_dsdc_n891));
   INV_X1 U_dsdc_U556 (.ZN(U_dsdc_n1543), 
	.A(U_dsdc_n1429));
   INV_X2 U_dsdc_U555 (.ZN(U_dsdc_n2076), 
	.A(U_dsdc_n2075));
   INV_X2 U_dsdc_U554 (.ZN(U_dsdc_n1579), 
	.A(U_dsdc_n1758));
   NAND2_X1 U_dsdc_U553 (.ZN(U_dsdc_n864), 
	.A2(U_dsdc_n181), 
	.A1(U_dsdc_n1031));
   OAI21_X1 U_dsdc_U552 (.ZN(U_dsdc_n393), 
	.B2(U_dsdc_n1734), 
	.B1(U_dsdc_xsr_cnt_7_), 
	.A(U_dsdc_n1731));
   NOR2_X1 U_dsdc_U551 (.ZN(U_dsdc_n1741), 
	.A2(U_dsdc_n1756), 
	.A1(U_dsdc_n1740));
   NAND3_X1 U_dsdc_U549 (.ZN(U_dsdc_n1869), 
	.A3(U_dsdc_n350), 
	.A2(U_dsdc_n1868), 
	.A1(U_dsdc_bm_bank_age_2__3_));
   NAND2_X1 U_dsdc_U546 (.ZN(U_dsdc_n646), 
	.A2(cr_mode_reg_update), 
	.A1(U_dsdc_n1429));
   OR3_X2 U_dsdc_U544 (.ZN(U_dsdc_n1321), 
	.A3(cr_t_rp[0]), 
	.A2(cr_t_rp[1]), 
	.A1(U_dsdc_n1336));
   AOI22_X1 U_dsdc_U543 (.ZN(U_dsdc_n1063), 
	.B2(U_dsdc_n1060), 
	.B1(U_dsdc_n1410), 
	.A2(U_dsdc_n1061), 
	.A1(U_dsdc_n1062));
   INV_X2 U_dsdc_U542 (.ZN(U_dsdc_n806), 
	.A(debug_ad_row_addr[15]));
   OAI211_X1 U_dsdc_U541 (.ZN(U_dsdc_n1317), 
	.C2(U_dsdc_n1315), 
	.C1(U_dsdc_n1316), 
	.B(U_dsdc_n1313), 
	.A(U_dsdc_n1314));
   NOR2_X2 U_dsdc_U540 (.ZN(U_dsdc_n1791), 
	.A2(U_dsdc_n2063), 
	.A1(U_dsdc_n573));
   NAND2_X2 U_dsdc_U539 (.ZN(U_dsdc_n1268), 
	.A2(U_dsdc_n1063), 
	.A1(U_dsdc_n1403));
   OAI211_X1 U_dsdc_U536 (.ZN(U_dsdc_n1366), 
	.C2(U_dsdc_n1360), 
	.C1(U_dsdc_n1361), 
	.B(U_dsdc_n1358), 
	.A(U_dsdc_n1359));
   AND2_X2 U_dsdc_U535 (.ZN(U_dsdc_n1977), 
	.A2(U_dsdc_n1409), 
	.A1(U_dsdc_n2013));
   OAI21_X1 U_dsdc_U533 (.ZN(U_dsdc_n2077), 
	.B2(U_dsdc_n2076), 
	.B1(U_dsdc_n2079), 
	.A(U_dsdc_early_term_flag));
   OAI21_X1 U_dsdc_U531 (.ZN(U_dsdc_n957), 
	.B2(debug_ref_req), 
	.B1(U_dsdc_n1372), 
	.A(U_dsdc_n1038));
   NAND2_X1 U_dsdc_U529 (.ZN(U_dsdc_n992), 
	.A2(U_dsdc_n1412), 
	.A1(U_dsdc_n864));
   OR2_X2 U_dsdc_U526 (.ZN(U_dsdc_n1495), 
	.A2(U_dsdc_n1601), 
	.A1(U_dsdc_n1612));
   NAND2_X1 U_dsdc_U525 (.ZN(U_dsdc_n576), 
	.A2(U_dsdc_row_cnt_12_), 
	.A1(U_dsdc_n1791));
   NOR3_X1 U_dsdc_U524 (.ZN(U_dsdc_n1356), 
	.A3(U_dsdc_n1348), 
	.A2(U_dsdc_access_cs_4_), 
	.A1(U_dsdc_n1507));
   NAND2_X1 U_dsdc_U523 (.ZN(U_dsdc_n583), 
	.A2(U_dsdc_row_cnt_6_), 
	.A1(U_dsdc_n1791));
   NAND2_X1 U_dsdc_U520 (.ZN(U_dsdc_n590), 
	.A2(U_dsdc_row_cnt_10_), 
	.A1(U_dsdc_n1791));
   INV_X1 U_dsdc_U518 (.ZN(U_dsdc_n1874), 
	.A(U_dsdc_n1875));
   NAND2_X1 U_dsdc_U517 (.ZN(U_dsdc_n591), 
	.A2(U_dsdc_row_cnt_4_), 
	.A1(U_dsdc_n1791));
   AOI22_X1 U_dsdc_U516 (.ZN(U_dsdc_n1262), 
	.B2(U_dsdc_r_burst_size_2_), 
	.B1(U_dsdc_n1269), 
	.A2(FE_PHN1227_U_dsdc_cas_cnt_2_), 
	.A1(U_dsdc_n1268));
   NAND2_X1 U_dsdc_U514 (.ZN(U_dsdc_n578), 
	.A2(U_dsdc_row_cnt_14_), 
	.A1(U_dsdc_n1791));
   NAND2_X1 U_dsdc_U511 (.ZN(U_dsdc_n577), 
	.A2(U_dsdc_row_cnt_2_), 
	.A1(U_dsdc_n1791));
   OR2_X2 U_dsdc_U509 (.ZN(U_dsdc_N430), 
	.A2(U_dsdc_n1495), 
	.A1(U_dsdc_n1581));
   INV_X2 U_dsdc_U508 (.ZN(U_dsdc_n767), 
	.A(U_dsdc_n992));
   NOR2_X1 U_dsdc_U507 (.ZN(U_dsdc_n1680), 
	.A2(U_dsdc_n1722), 
	.A1(U_dsdc_n1679));
   OR2_X2 U_dsdc_U503 (.ZN(U_dsdc_n1608), 
	.A2(U_dsdc_n1596), 
	.A1(U_dsdc_n1603));
   NAND2_X1 U_dsdc_U502 (.ZN(U_dsdc_n592), 
	.A2(U_dsdc_row_cnt_8_), 
	.A1(U_dsdc_n1791));
   INV_X2 U_dsdc_U498 (.ZN(U_dsdc_n1783), 
	.A(U_dsdc_n588));
   INV_X1 U_dsdc_U497 (.ZN(U_dsdc_n1098), 
	.A(debug_ad_row_addr[6]));
   INV_X2 U_dsdc_U496 (.ZN(U_dsdc_n594), 
	.A(U_dsdc_n584));
   NAND2_X1 U_dsdc_U495 (.ZN(U_dsdc_n1318), 
	.A2(U_dsdc_n1650), 
	.A1(U_dsdc_n1417));
   INV_X1 U_dsdc_U493 (.ZN(U_dsdc_n1111), 
	.A(debug_ad_row_addr[4]));
   INV_X2 U_dsdc_U491 (.ZN(U_dsdc_n595), 
	.A(U_dsdc_n587));
   NAND4_X1 U_dsdc_U490 (.ZN(U_dsdc_n921), 
	.A4(U_dsdc_n1449), 
	.A3(U_dsdc_n1038), 
	.A2(U_dsdc_n1428), 
	.A1(FE_PHN2909_U_dsdc_n1436));
   OAI22_X1 U_dsdc_U489 (.ZN(U_dsdc_n1261), 
	.B2(U_dsdc_n182), 
	.B1(U_dsdc_n1259), 
	.A2(FE_PHN1035_U_dsdc_n327), 
	.A1(U_dsdc_n1260));
   INV_X2 U_dsdc_U488 (.ZN(U_dsdc_n800), 
	.A(debug_ad_row_addr[13]));
   OAI211_X1 U_dsdc_U486 (.ZN(U_dsdc_n1678), 
	.C2(U_dsdc_n1686), 
	.C1(U_dsdc_init_cnt_12_), 
	.B(U_dsdc_n1676), 
	.A(U_dsdc_init_cnt_13_));
   INV_X2 U_dsdc_U485 (.ZN(U_dsdc_n1771), 
	.A(U_dsdc_n582));
   AOI21_X1 U_dsdc_U484 (.ZN(U_dsdc_n1600), 
	.B2(U_dsdc_n1602), 
	.B1(cr_t_rcar[0]), 
	.A(U_dsdc_n1601));
   OR3_X2 U_dsdc_U483 (.ZN(U_dsdc_n1675), 
	.A3(U_dsdc_n482), 
	.A2(U_dsdc_init_cnt_14_), 
	.A1(U_dsdc_init_cnt_15_));
   INV_X1 U_dsdc_U482 (.ZN(U_dsdc_n1028), 
	.A(debug_ad_row_addr[10]));
   INV_X2 U_dsdc_U480 (.ZN(U_dsdc_n593), 
	.A(U_dsdc_n586));
   INV_X1 U_dsdc_U479 (.ZN(U_dsdc_n1076), 
	.A(debug_ad_row_addr[8]));
   OAI22_X1 U_dsdc_U478 (.ZN(U_dsdc_rcar_cnt1_nxt[3]), 
	.B2(U_dsdc_n1588), 
	.B1(U_dsdc_n1589), 
	.A2(U_cr_n72), 
	.A1(U_dsdc_n1590));
   INV_X2 U_dsdc_U477 (.ZN(U_dsdc_n1611), 
	.A(U_dsdc_n1610));
   INV_X4 U_dsdc_U476 (.ZN(U_dsdc_n1127), 
	.A(debug_ad_bank_addr[0]));
   OAI22_X1 U_dsdc_U475 (.ZN(U_dsdc_rcar_cnt1_nxt[2]), 
	.B2(U_dsdc_n1588), 
	.B1(U_dsdc_n1586), 
	.A2(FE_PHN1407_U_cr_n104), 
	.A1(U_dsdc_n1590));
   INV_X2 U_dsdc_U473 (.ZN(U_dsdc_n1000), 
	.A(U_dsdc_oldest_bank_1_));
   XNOR2_X1 U_dsdc_U472 (.ZN(U_dsdc_num_row[9]), 
	.B(U_dsdc_n358), 
	.A(U_dsdc_n618));
   INV_X1 U_dsdc_U471 (.ZN(U_dsdc_n1847), 
	.A(U_dsdc_n1849));
   OAI21_X1 U_dsdc_U470 (.ZN(U_dsdc_rcar_cnt2_nxt[0]), 
	.B2(U_dsdc_n1597), 
	.B1(U_dsdc_rcar_cnt2_0_), 
	.A(FE_PHN3463_U_dsdc_n1594));
   INV_X1 U_dsdc_U469 (.ZN(U_dsdc_n1888), 
	.A(U_dsdc_n1890));
   OAI22_X1 U_dsdc_U468 (.ZN(U_dsdc_rcar_cnt1_nxt[1]), 
	.B2(U_dsdc_n1588), 
	.B1(U_dsdc_n1582), 
	.A2(FE_PHN1482_U_cr_n151), 
	.A1(U_dsdc_n1590));
   INV_X2 U_dsdc_U467 (.ZN(U_dsdc_n1545), 
	.A(U_dsdc_n1542));
   INV_X1 U_dsdc_U465 (.ZN(U_dsdc_n1918), 
	.A(U_dsdc_n1920));
   AOI21_X1 U_dsdc_U464 (.ZN(U_dsdc_n1848), 
	.B2(U_dsdc_n1849), 
	.B1(U_dsdc_n1867), 
	.A(U_dsdc_n1850));
   OAI21_X1 U_dsdc_U459 (.ZN(U_dsdc_DP_OP_1642_126_2028_I5_2_), 
	.B2(U_dsdc_n1263), 
	.B1(U_dsdc_n1546), 
	.A(U_dsdc_n750));
   OAI21_X1 U_dsdc_U457 (.ZN(U_dsdc_DP_OP_1642_126_2028_I5_4_), 
	.B2(U_dmc_n16), 
	.B1(U_dsdc_n1546), 
	.A(U_dsdc_n748));
   NOR2_X1 U_dsdc_U456 (.ZN(U_dsdc_n1695), 
	.A2(U_dsdc_n1724), 
	.A1(U_dsdc_n1694));
   NOR2_X1 U_dsdc_U454 (.ZN(U_dsdc_n1702), 
	.A2(U_dsdc_n1724), 
	.A1(U_dsdc_n1701));
   NOR2_X1 U_dsdc_U453 (.ZN(U_dsdc_n1709), 
	.A2(U_dsdc_n1724), 
	.A1(U_dsdc_n1708));
   NOR2_X1 U_dsdc_U452 (.ZN(U_dsdc_n1688), 
	.A2(U_dsdc_n1724), 
	.A1(U_dsdc_n1687));
   OAI211_X2 U_dsdc_U451 (.ZN(U_dsdc_n2093), 
	.C2(U_dsdc_n432), 
	.C1(U_dsdc_n1545), 
	.B(U_dsdc_n1543), 
	.A(U_dsdc_n1544));
   OAI211_X1 U_dsdc_U450 (.ZN(U_dsdc_n416), 
	.C2(U_dsdc_n482), 
	.C1(U_dsdc_n1724), 
	.B(U_dsdc_n1677), 
	.A(U_dsdc_n1678));
   OAI21_X1 U_dsdc_U449 (.ZN(U_dsdc_n404), 
	.B2(U_dsdc_n1724), 
	.B1(U_dsdc_n1721), 
	.A(U_dsdc_n1720));
   OAI21_X1 U_dsdc_U448 (.ZN(U_dsdc_n403), 
	.B2(U_dsdc_n1724), 
	.B1(U_dsdc_init_cnt_0_), 
	.A(U_dsdc_n1723));
   INV_X2 U_dsdc_U444 (.ZN(U_dsdc_n1897), 
	.A(U_dsdc_n1902));
   INV_X2 U_dsdc_U443 (.ZN(U_dsdc_n2012), 
	.A(U_dsdc_n1396));
   INV_X2 U_dsdc_U442 (.ZN(U_dsdc_n754), 
	.A(U_dsdc_n753));
   OAI21_X1 U_dsdc_U441 (.ZN(U_dsdc_n1718), 
	.B2(U_dsdc_init_cnt_1_), 
	.B1(U_dsdc_init_cnt_0_), 
	.A(U_dsdc_n1715));
   INV_X2 U_dsdc_U440 (.ZN(U_dsdc_n2084), 
	.A(U_dsdc_n2083));
   OAI211_X1 U_dsdc_U439 (.ZN(U_dsdc_n1706), 
	.C2(U_dsdc_n1704), 
	.C1(U_dsdc_init_cnt_4_), 
	.B(U_dsdc_n1715), 
	.A(FE_PHN971_U_dsdc_init_cnt_5_));
   XNOR2_X1 U_dsdc_U438 (.ZN(U_dsdc_num_row[11]), 
	.B(U_dsdc_n357), 
	.A(U_dsdc_n607));
   INV_X2 U_dsdc_U437 (.ZN(U_dsdc_n1857), 
	.A(U_dsdc_n1862));
   OAI211_X1 U_dsdc_U436 (.ZN(U_dsdc_n1699), 
	.C2(U_dsdc_n1697), 
	.C1(U_dsdc_init_cnt_6_), 
	.B(U_dsdc_n1715), 
	.A(FE_PHN1031_U_dsdc_init_cnt_7_));
   OR2_X2 U_dsdc_U435 (.ZN(U_dsdc_n1957), 
	.A2(U_dsdc_n1962), 
	.A1(U_dsdc_n1965));
   NAND2_X1 U_dsdc_U434 (.ZN(U_dsdc_n1691), 
	.A2(U_dsdc_n1715), 
	.A1(U_dsdc_n1687));
   OAI211_X1 U_dsdc_U432 (.ZN(U_dsdc_n1692), 
	.C2(U_dsdc_n1690), 
	.C1(U_dsdc_init_cnt_8_), 
	.B(U_dsdc_n1715), 
	.A(FE_PHN1032_U_dsdc_init_cnt_9_));
   OAI211_X1 U_dsdc_U430 (.ZN(U_dsdc_n1685), 
	.C2(U_dsdc_n1683), 
	.C1(FE_PHN3268_U_dsdc_init_cnt_10_), 
	.B(U_dsdc_n1715), 
	.A(FE_PHN970_U_dsdc_init_cnt_11_));
   INV_X2 U_dsdc_U429 (.ZN(U_dsdc_n1927), 
	.A(U_dsdc_n1932));
   NAND2_X1 U_dsdc_U428 (.ZN(U_dsdc_n1682), 
	.A2(U_dsdc_n1715), 
	.A1(U_dsdc_n1679));
   INV_X2 U_dsdc_U426 (.ZN(U_dsdc_DP_OP_1642_126_2028_I5_3_), 
	.A(U_dsdc_n749));
   INV_X2 U_dsdc_U425 (.ZN(U_dsdc_n1864), 
	.A(U_dsdc_n1865));
   INV_X2 U_dsdc_U424 (.ZN(U_dsdc_n1963), 
	.A(U_dsdc_n1968));
   INV_X2 U_dsdc_U422 (.ZN(U_dsdc_DP_OP_1642_126_2028_I5_5_), 
	.A(U_dsdc_n747));
   INV_X2 U_dsdc_U420 (.ZN(U_dsdc_n1904), 
	.A(U_dsdc_n1905));
   INV_X2 U_dsdc_U416 (.ZN(U_dsdc_n1934), 
	.A(U_dsdc_n1935));
   OAI21_X1 U_dsdc_U415 (.ZN(U_dsdc_n415), 
	.B2(U_dsdc_n1682), 
	.B1(U_dsdc_init_cnt_12_), 
	.A(U_dsdc_n1681));
   OAI211_X1 U_dsdc_U414 (.ZN(U_dsdc_n1516), 
	.C2(U_dsdc_n1505), 
	.C1(U_dsdc_n1430), 
	.B(U_dsdc_n1504), 
	.A(U_dsdc_n2060));
   OAI21_X1 U_dsdc_U413 (.ZN(U_dsdc_n409), 
	.B2(U_dsdc_n1705), 
	.B1(U_dsdc_init_cnt_6_), 
	.A(U_dsdc_n1703));
   OAI211_X1 U_dsdc_U412 (.ZN(U_dsdc_n414), 
	.C2(U_dsdc_n1686), 
	.C1(U_dsdc_n1724), 
	.B(U_dsdc_n1684), 
	.A(U_dsdc_n1685));
   INV_X2 U_dsdc_U411 (.ZN(U_dsdc_n720), 
	.A(U_dsdc_n2067));
   OAI21_X1 U_dsdc_U410 (.ZN(U_dsdc_n413), 
	.B2(U_dsdc_n1691), 
	.B1(FE_PHN3268_U_dsdc_init_cnt_10_), 
	.A(U_dsdc_n1689));
   OAI21_X1 U_dsdc_U409 (.ZN(U_dsdc_n411), 
	.B2(U_dsdc_n1698), 
	.B1(U_dsdc_init_cnt_8_), 
	.A(U_dsdc_n1696));
   AOI22_X1 U_dsdc_U407 (.ZN(U_dsdc_n2047), 
	.B2(U_dsdc_n2048), 
	.B1(hiu_burst_size[5]), 
	.A2(FE_PHN1890_U_dsdc_r_burst_size_5_), 
	.A1(U_dsdc_n2049));
   AOI22_X1 U_dsdc_U406 (.ZN(U_dsdc_n2043), 
	.B2(U_dsdc_n2048), 
	.B1(hiu_burst_size[1]), 
	.A2(FE_PHN1896_U_dsdc_r_burst_size_1_), 
	.A1(U_dsdc_n2049));
   AOI22_X1 U_dsdc_U405 (.ZN(U_dsdc_n2045), 
	.B2(U_dsdc_n2048), 
	.B1(hiu_burst_size[3]), 
	.A2(FE_PHN1892_U_dsdc_r_burst_size_3_), 
	.A1(U_dsdc_n2049));
   AOI22_X1 U_dsdc_U404 (.ZN(U_dsdc_n2042), 
	.B2(U_dsdc_n2048), 
	.B1(hiu_burst_size[0]), 
	.A2(U_dsdc_r_burst_size_0_), 
	.A1(U_dsdc_n2049));
   AOI22_X1 U_dsdc_U403 (.ZN(U_dsdc_n2046), 
	.B2(U_dsdc_n2048), 
	.B1(hiu_burst_size[4]), 
	.A2(FE_PHN1888_U_dsdc_r_burst_size_4_), 
	.A1(U_dsdc_n2049));
   INV_X4 U_dsdc_U402 (.ZN(U_dsdc_n978), 
	.A(U_dsdc_n987));
   AOI22_X1 U_dsdc_U401 (.ZN(U_dsdc_n2050), 
	.B2(U_dsdc_n2048), 
	.B1(hiu_wrapped_burst), 
	.A2(U_dsdc_r_wrapped_burst), 
	.A1(U_dsdc_n2049));
   INV_X2 U_dsdc_U400 (.ZN(U_dsdc_n1970), 
	.A(U_dsdc_n1971));
   AOI22_X1 U_dsdc_U399 (.ZN(U_dsdc_n2044), 
	.B2(U_dsdc_n2048), 
	.B1(hiu_burst_size[2]), 
	.A2(U_dsdc_r_burst_size_2_), 
	.A1(U_dsdc_n2049));
   AND2_X2 U_dsdc_U397 (.ZN(U_dsdc_n176), 
	.A2(U_dsdc_n604), 
	.A1(U_dsdc_bm_row_addr_1__10_));
   INV_X2 U_dsdc_U396 (.ZN(U_dsdc_n1266), 
	.A(U_dsdc_n1270));
   OAI211_X1 U_dsdc_U395 (.ZN(U_dsdc_n1355), 
	.C2(U_dsdc_n1353), 
	.C1(U_dsdc_n1354), 
	.B(U_dsdc_n1351), 
	.A(U_dsdc_n1352));
   INV_X2 U_dsdc_U394 (.ZN(U_dsdc_n2068), 
	.A(U_dsdc_n1395));
   INV_X2 U_dsdc_U392 (.ZN(U_dsdc_n1341), 
	.A(FE_PHN1161_U_dsdc_n1339));
   NAND2_X1 U_dsdc_U391 (.ZN(U_dsdc_n797), 
	.A2(U_dsdc_bm_row_addr_3__7_), 
	.A1(U_dsdc_n978));
   OAI211_X1 U_dsdc_U390 (.ZN(U_dsdc_n2095), 
	.C2(U_dsdc_n341), 
	.C1(U_dsdc_n1541), 
	.B(U_dsdc_n1539), 
	.A(FE_PHN771_U_dsdc_n1540));
   INV_X2 U_dsdc_U389 (.ZN(U_dsdc_n275), 
	.A(U_dsdc_n2046));
   INV_X2 U_dsdc_U388 (.ZN(U_dsdc_n276), 
	.A(U_dsdc_n2047));
   INV_X2 U_dsdc_U387 (.ZN(U_dsdc_n277), 
	.A(U_dsdc_n2050));
   NAND2_X1 U_dsdc_U386 (.ZN(U_dsdc_n778), 
	.A2(U_dsdc_bm_row_addr_3__13_), 
	.A1(U_dsdc_n978));
   OAI21_X1 U_dsdc_U385 (.ZN(U_dsdc_n831), 
	.B2(U_dsdc_bm_rc_cnt_3__3_), 
	.B1(U_dsdc_bm_rc_cnt_3__2_), 
	.A(U_dsdc_n978));
   INV_X2 U_dsdc_U384 (.ZN(U_dsdc_n274), 
	.A(U_dsdc_n2045));
   INV_X2 U_dsdc_U383 (.ZN(U_dsdc_n273), 
	.A(U_dsdc_n2044));
   AOI22_X1 U_dsdc_U382 (.ZN(U_dsdc_n1991), 
	.B2(U_dsdc_n2048), 
	.B1(debug_ad_col_addr_1_), 
	.A2(FE_PHN1416_U_dsdc_r_col_addr_1_), 
	.A1(U_dsdc_n2007));
   INV_X2 U_dsdc_U381 (.ZN(U_dsdc_n272), 
	.A(U_dsdc_n2043));
   OAI21_X1 U_dsdc_U379 (.ZN(U_dsdc_n1346), 
	.B2(U_dsdc_n1483), 
	.B1(U_dsdc_n2068), 
	.A(U_dsdc_r_chip_slct_0_));
   INV_X2 U_dsdc_U378 (.ZN(U_dsdc_n271), 
	.A(U_dsdc_n2042));
   INV_X2 U_dsdc_U374 (.ZN(U_dsdc_n240), 
	.A(U_dsdc_n1991));
   INV_X1 U_dsdc_U373 (.ZN(U_dsdc_n1288), 
	.A(U_dsdc_n1283));
   AND4_X2 U_dsdc_U371 (.ZN(U_dsdc_n835), 
	.A4(U_dsdc_n829), 
	.A3(U_dsdc_n830), 
	.A2(U_dsdc_n831), 
	.A1(U_dsdc_n832));
   INV_X2 U_dsdc_U370 (.ZN(U_dsdc_n809), 
	.A(U_dsdc_n808));
   AND2_X2 U_dsdc_U369 (.ZN(U_dsdc_n333), 
	.A2(U_dsdc_n800), 
	.A1(U_dsdc_n785));
   OR3_X2 U_dsdc_U368 (.ZN(U_dsdc_n332), 
	.A3(U_dsdc_bm_row_addr_0__7_), 
	.A2(U_dsdc_n816), 
	.A1(U_dsdc_n602));
   AND2_X2 U_dsdc_U367 (.ZN(U_dsdc_n318), 
	.A2(debug_ad_row_addr[1]), 
	.A1(U_dsdc_n813));
   NAND2_X1 U_dsdc_U366 (.ZN(U_dsdc_n997), 
	.A2(FE_PHN1593_U_dsdc_bm_bank_status_1_), 
	.A1(FE_PHN683_U_dsdc_n1394));
   NAND2_X1 U_dsdc_U365 (.ZN(U_dsdc_n996), 
	.A2(U_dsdc_bm_bank_status_3_), 
	.A1(FE_PHN683_U_dsdc_n1394));
   NAND2_X1 U_dsdc_U364 (.ZN(U_dsdc_n1002), 
	.A2(U_dsdc_bm_bank_status_0_), 
	.A1(FE_PHN683_U_dsdc_n1394));
   NAND2_X1 U_dsdc_U363 (.ZN(U_dsdc_n1392), 
	.A2(U_dsdc_bm_bank_status_2_), 
	.A1(FE_PHN683_U_dsdc_n1394));
   INV_X2 U_dsdc_U362 (.ZN(U_dsdc_n1322), 
	.A(FE_PHN683_U_dsdc_n1394));
   AND2_X2 U_dsdc_U361 (.ZN(U_dsdc_n177), 
	.A2(U_dsdc_n425), 
	.A1(U_dsdc_n533));
   INV_X2 U_dsdc_U360 (.ZN(U_dsdc_n817), 
	.A(U_dsdc_n818));
   NAND3_X1 U_dsdc_U359 (.ZN(U_dsdc_n847), 
	.A3(U_dsdc_n982), 
	.A2(U_dsdc_n984), 
	.A1(U_dsdc_n986));
   NAND3_X1 U_dsdc_U358 (.ZN(U_dsdc_n985), 
	.A3(U_dsdc_n982), 
	.A2(U_dsdc_n983), 
	.A1(U_dsdc_n984));
   NAND2_X1 U_dsdc_U357 (.ZN(U_dsdc_n910), 
	.A2(U_dsdc_n828), 
	.A1(U_dsdc_n975));
   NAND3_X1 U_dsdc_U356 (.ZN(U_dsdc_n1001), 
	.A3(U_dsdc_n999), 
	.A2(U_dsdc_n1000), 
	.A1(U_dsdc_n1003));
   NAND2_X2 U_dsdc_U355 (.ZN(U_dsdc_n1112), 
	.A2(U_dsdc_n977), 
	.A1(U_dsdc_n1345));
   NAND2_X2 U_dsdc_U354 (.ZN(U_dsdc_n1166), 
	.A2(U_dsdc_n1136), 
	.A1(U_dsdc_n1112));
   INV_X2 U_dsdc_U352 (.ZN(U_dsdc_n1159), 
	.A(U_dsdc_n1166));
   INV_X2 U_dsdc_U351 (.ZN(U_dsdc_n1012), 
	.A(U_dsdc_n1020));
   NOR3_X1 U_dsdc_U350 (.ZN(U_dsdc_n1021), 
	.A3(U_dsdc_n338), 
	.A2(U_dsdc_n179), 
	.A1(U_dsdc_n1020));
   OAI21_X1 U_dsdc_U349 (.ZN(U_dsdc_N4449), 
	.B2(FE_PHN1893_U_dsdc_n1392), 
	.B1(U_dsdc_bm_close_bank_2_), 
	.A(U_dsdc_n310));
   OAI21_X1 U_dsdc_U347 (.ZN(U_dsdc_N4496), 
	.B2(FE_PHN1895_U_dsdc_n996), 
	.B1(U_dsdc_bm_close_bank_3_), 
	.A(U_dsdc_n313));
   INV_X2 U_dsdc_U346 (.ZN(U_dsdc_n894), 
	.A(U_dsdc_n960));
   INV_X2 U_dsdc_U345 (.ZN(U_dsdc_n1013), 
	.A(U_dsdc_n1017));
   INV_X1 U_dsdc_U343 (.ZN(U_dsdc_n1327), 
	.A(U_dsdc_n1328));
   NAND3_X1 U_dsdc_U340 (.ZN(U_dsdc_n[2089]), 
	.A3(U_dsdc_n1319), 
	.A2(U_dsdc_n1320), 
	.A1(U_dsdc_n1389));
   OR3_X2 U_dsdc_U338 (.ZN(U_dsdc_N429), 
	.A3(U_dsdc_n963), 
	.A2(U_dsdc_n1374), 
	.A1(hiu_terminate));
   INV_X1 U_dsdc_U337 (.ZN(U_dsdc_n1376), 
	.A(U_dsdc_n1374));
   INV_X2 U_dsdc_U336 (.ZN(U_dsdc_n1052), 
	.A(U_dsdc_n1051));
   OR2_X2 U_dsdc_U335 (.ZN(U_dsdc_n603), 
	.A2(U_dsdc_n1026), 
	.A1(U_dsdc_bm_num_open_bank_4_));
   NAND2_X2 U_dsdc_U331 (.ZN(U_dsdc_n649), 
	.A2(U_dsdc_n355), 
	.A1(U_dsdc_n173));
   NOR2_X1 U_dsdc_U330 (.ZN(U_dsdc_n1719), 
	.A2(U_dsdc_init_cnt_1_), 
	.A1(U_dsdc_init_cnt_0_));
   XNOR2_X1 U_dsdc_U328 (.ZN(U_dsdc_n1246), 
	.B(U_dsdc_wtr_cnt_0_), 
	.A(U_dsdc_n194));
   NOR2_X1 U_dsdc_U327 (.ZN(U_dsdc_n1583), 
	.A2(U_dsdc_rcar_cnt1_0_), 
	.A1(U_dsdc_rcar_cnt1_1_));
   NAND2_X2 U_dsdc_U326 (.ZN(U_dsdc_n690), 
	.A2(U_dsdc_access_cs_0_), 
	.A1(U_dsdc_n355));
   INV_X2 U_dsdc_U325 (.ZN(U_dsdc_n598), 
	.A(U_dsdc_N4239));
   INV_X2 U_dsdc_U324 (.ZN(U_dsdc_n1704), 
	.A(U_dsdc_n1708));
   INV_X2 U_dsdc_U322 (.ZN(U_dsdc_n1227), 
	.A(U_dsdc_n1234));
   INV_X2 U_dsdc_U321 (.ZN(U_dsdc_n1188), 
	.A(U_dsdc_n1193));
   INV_X2 U_dsdc_U320 (.ZN(U_dsdc_n1202), 
	.A(U_dsdc_n1207));
   INV_X2 U_dsdc_U319 (.ZN(U_dsdc_n1174), 
	.A(U_dsdc_n1179));
   NAND2_X1 U_dsdc_U318 (.ZN(U_dsdc_n1292), 
	.A2(U_dsdc_n657), 
	.A1(U_dsdc_n1458));
   NAND2_X1 U_dsdc_U317 (.ZN(U_dsdc_n1505), 
	.A2(U_dsdc_n1435), 
	.A1(U_dsdc_n1434));
   INV_X2 U_dsdc_U316 (.ZN(U_dsdc_n865), 
	.A(U_dsdc_n1650));
   NAND2_X1 U_dsdc_U315 (.ZN(U_dsdc_n1343), 
	.A2(U_dsdc_n1426), 
	.A1(U_dsdc_n360));
   NOR2_X1 U_dsdc_U314 (.ZN(U_dsdc_n1591), 
	.A2(U_dsdc_n1803), 
	.A1(U_dsdc_n1422));
   INV_X2 U_dsdc_U313 (.ZN(U_dsdc_n1697), 
	.A(U_dsdc_n1701));
   INV_X2 U_dsdc_U312 (.ZN(U_dsdc_n2065), 
	.A(U_dsdc_n1526));
   OAI21_X1 U_dsdc_U311 (.ZN(U_dsdc_n1922), 
	.B2(U_dsdc_n1930), 
	.B1(FE_PHN897_U_dsdc_n352), 
	.A(U_dsdc_n335));
   INV_X2 U_dsdc_U310 (.ZN(U_dsdc_n1060), 
	.A(U_dsdc_n933));
   INV_X2 U_dsdc_U309 (.ZN(U_dsdc_n869), 
	.A(U_dsdc_n945));
   INV_X2 U_dsdc_U308 (.ZN(U_dsdc_n1733), 
	.A(U_dsdc_n1754));
   INV_X2 U_dsdc_U307 (.ZN(U_dsdc_n1089), 
	.A(FE_PHN1249_U_dsdc_add_x_2600_1_n8));
   INV_X2 U_dsdc_U306 (.ZN(U_dsdc_n994), 
	.A(U_dsdc_n856));
   NAND3_X1 U_dsdc_U305 (.ZN(U_dsdc_n1861), 
	.A3(U_dsdc_bm_bank_age_2__0_), 
	.A2(U_dsdc_bm_bank_age_2__1_), 
	.A1(U_dsdc_n1866));
   NAND2_X1 U_dsdc_U304 (.ZN(U_dsdc_n1684), 
	.A2(U_dsdc_n1722), 
	.A1(cr_t_init[11]));
   NAND2_X1 U_dsdc_U303 (.ZN(U_dsdc_n1677), 
	.A2(U_dsdc_n1722), 
	.A1(cr_t_init[13]));
   NAND2_X1 U_dsdc_U302 (.ZN(U_dsdc_n672), 
	.A2(U_dsdc_n758), 
	.A1(U_dsdc_n1556));
   INV_X2 U_dsdc_U301 (.ZN(U_dsdc_n826), 
	.A(U_dsdc_n982));
   NAND2_X1 U_dsdc_U300 (.ZN(U_dsdc_n1909), 
	.A2(U_dsdc_n1908), 
	.A1(U_dsdc_bm_bank_age_3__3_));
   INV_X4 U_dsdc_U299 (.ZN(U_dsdc_n685), 
	.A(U_dsdc_n1629));
   INV_X2 U_dsdc_U298 (.ZN(U_dsdc_n1690), 
	.A(U_dsdc_n1694));
   NAND2_X1 U_dsdc_U297 (.ZN(U_dsdc_n1744), 
	.A2(U_dsdc_n1750), 
	.A1(U_dsdc_n1740));
   INV_X2 U_dsdc_U295 (.ZN(U_dsdc_n1683), 
	.A(U_dsdc_n1687));
   INV_X2 U_dsdc_U294 (.ZN(U_dsdc_n755), 
	.A(U_dsdc_DP_OP_1642_126_2028_I4));
   OAI21_X1 U_dsdc_U291 (.ZN(U_dsdc_n386), 
	.B2(U_dsdc_n1756), 
	.B1(U_dsdc_xsr_cnt_0_), 
	.A(U_dsdc_n1755));
   OAI211_X1 U_dsdc_U290 (.ZN(U_dsdc_auto_ref_en_nxt), 
	.C2(U_dsdc_n2063), 
	.C1(U_dsdc_n1492), 
	.B(U_dsdc_n1488), 
	.A(FE_PHN771_U_dsdc_n1540));
   INV_X1 U_dsdc_U289 (.ZN(U_dsdc_n1529), 
	.A(U_dsdc_n1525));
   NOR2_X1 U_dsdc_U286 (.ZN(U_dsdc_n1449), 
	.A2(sdram_req_i), 
	.A1(debug_ref_req));
   INV_X4 U_dsdc_U285 (.ZN(U_dsdc_n1382), 
	.A(U_dsdc_n764));
   NAND2_X1 U_dsdc_U283 (.ZN(U_dsdc_n589), 
	.A2(U_dsdc_n575), 
	.A1(U_dsdc_n1791));
   NAND2_X1 U_dsdc_U282 (.ZN(U_dsdc_n584), 
	.A2(U_dsdc_n580), 
	.A1(U_dsdc_n1791));
   INV_X1 U_dsdc_U280 (.ZN(U_dsdc_n1796), 
	.A(U_dsdc_n589));
   AND2_X2 U_dsdc_U279 (.ZN(U_dsdc_n1352), 
	.A2(U_dsdc_n852), 
	.A1(U_dsdc_n921));
   NAND2_X1 U_dsdc_U278 (.ZN(U_dsdc_n1698), 
	.A2(U_dsdc_n1715), 
	.A1(U_dsdc_n1694));
   OAI21_X1 U_dsdc_U276 (.ZN(U_dsdc_n407), 
	.B2(U_dsdc_n1712), 
	.B1(U_dsdc_init_cnt_4_), 
	.A(U_dsdc_n1710));
   NAND2_X1 U_dsdc_U275 (.ZN(U_dsdc_n776), 
	.A2(U_dsdc_bm_row_addr_1__13_), 
	.A1(U_dsdc_n604));
   NAND2_X1 U_dsdc_U273 (.ZN(U_dsdc_n795), 
	.A2(U_dsdc_bm_row_addr_1__7_), 
	.A1(U_dsdc_n604));
   NAND2_X1 U_dsdc_U272 (.ZN(U_dsdc_n786), 
	.A2(U_dsdc_bm_row_addr_1__9_), 
	.A1(U_dsdc_n604));
   INV_X4 U_dsdc_U271 (.ZN(U_dsdc_n159), 
	.A(U_dsdc_n599));
   NAND2_X1 U_dsdc_U270 (.ZN(U_dsdc_n516), 
	.A2(U_dsdc_bm_row_addr_3__12_), 
	.A1(U_dsdc_n978));
   OAI21_X1 U_dsdc_U269 (.ZN(U_dsdc_n832), 
	.B2(U_dsdc_bm_rc_cnt_2__3_), 
	.B1(U_dsdc_bm_rc_cnt_2__2_), 
	.A(U_dsdc_n159));
   NAND2_X1 U_dsdc_U268 (.ZN(U_dsdc_n777), 
	.A2(U_dsdc_bm_row_addr_2__13_), 
	.A1(U_dsdc_n159));
   NAND2_X1 U_dsdc_U267 (.ZN(U_dsdc_n788), 
	.A2(U_dsdc_bm_row_addr_3__9_), 
	.A1(U_dsdc_n978));
   NAND2_X1 U_dsdc_U266 (.ZN(U_dsdc_n796), 
	.A2(U_dsdc_bm_row_addr_2__7_), 
	.A1(U_dsdc_n159));
   OAI21_X1 U_dsdc_U264 (.ZN(U_dsdc_n830), 
	.B2(U_dsdc_bm_rc_cnt_1__3_), 
	.B1(FE_PHN1221_U_dsdc_bm_rc_cnt_1__2_), 
	.A(U_dsdc_n604));
   INV_X2 U_dsdc_U263 (.ZN(U_dsdc_n372), 
	.A(U_dsdc_n1782));
   NAND2_X4 U_dsdc_U261 (.ZN(U_dsdc_n313), 
	.A2(U_dsdc_n978), 
	.A1(U_dsdc_n1166));
   NOR3_X1 U_dsdc_U260 (.ZN(U_dsdc_n1018), 
	.A3(U_dsdc_n338), 
	.A2(U_dsdc_bm_num_open_bank_3_), 
	.A1(U_dsdc_n1020));
   OAI22_X1 U_dsdc_U259 (.ZN(U_dsdc_N4461), 
	.B2(U_cr_n120), 
	.B1(U_dsdc_n313), 
	.A2(FE_PHN3255_U_dsdc_n1241), 
	.A1(U_dsdc_n1243));
   OAI22_X1 U_dsdc_U258 (.ZN(U_dsdc_N4460), 
	.B2(n95), 
	.B1(U_dsdc_n313), 
	.A2(FE_PHN3513_U_dsdc_bm_ras_cnt_3__0_), 
	.A1(U_dsdc_n1243));
   NOR2_X2 U_dsdc_U257 (.ZN(U_dsdc_n981), 
	.A2(U_dsdc_n817), 
	.A1(U_dsdc_n887));
   NOR3_X1 U_dsdc_U256 (.ZN(U_dsdc_n1311), 
	.A3(U_dsdc_n1309), 
	.A2(cr_delayed_precharge), 
	.A1(U_dsdc_n1310));
   OAI21_X1 U_dsdc_U254 (.ZN(U_dsdc_N4355), 
	.B2(FE_PHN1897_U_dsdc_n1002), 
	.B1(U_dsdc_bm_close_bank_0_), 
	.A(n83));
   NOR3_X1 U_dsdc_U253 (.ZN(U_dsdc_n1287), 
	.A3(U_dsdc_n1557), 
	.A2(U_dsdc_n1285), 
	.A1(U_dsdc_n1286));
   OAI21_X1 U_dsdc_U252 (.ZN(U_dsdc_N4402), 
	.B2(U_dsdc_n997), 
	.B1(U_dsdc_bm_close_bank_1_), 
	.A(U_dsdc_n620));
   OAI21_X2 U_dsdc_U251 (.ZN(U_dsdc_n293), 
	.B2(FE_PHN1093_U_dsdc_n340), 
	.B1(U_dsdc_n1006), 
	.A(U_dsdc_n1005));
   NAND2_X4 U_dsdc_U250 (.ZN(U_dsdc_n310), 
	.A2(U_dsdc_n159), 
	.A1(U_dsdc_n1166));
   AOI22_X1 U_dsdc_U249 (.ZN(U_dsdc_n554), 
	.B2(U_dsdc_n158), 
	.B1(U_dsdc_n1093), 
	.A2(s_read_pipe[2]), 
	.A1(FE_PHN893_U_dsdc_n1092));
   INV_X1 U_dsdc_U248 (.ZN(U_dsdc_n158), 
	.A(FE_PHN1596_U_dsdc_n1091));
   XOR2_X1 U_dsdc_U247 (.Z(U_dsdc_cas_latency_1_), 
	.B(FE_PHN1921_U_dsdc_n1084), 
	.A(FE_PHN1020_U_dsdc_n1085));
   NAND2_X1 U_dsdc_U246 (.ZN(U_dsdc_n[2091]), 
	.A2(FE_PHN1445_U_dsdc_n157), 
	.A1(U_dsdc_n1393));
   AOI211_X1 U_dsdc_U245 (.ZN(U_dsdc_n157), 
	.C2(U_dsdc_n154), 
	.C1(U_dsdc_access_cs_1_), 
	.B(U_dsdc_n156), 
	.A(U_dsdc_n1388));
   OAI211_X1 U_dsdc_U244 (.ZN(U_dsdc_n156), 
	.C2(U_dsdc_n155), 
	.C1(cr_delayed_precharge), 
	.B(U_dsdc_n1389), 
	.A(U_dsdc_n1387));
   INV_X1 U_dsdc_U243 (.ZN(U_dsdc_n155), 
	.A(U_dsdc_n1386));
   NAND3_X1 U_dsdc_U242 (.ZN(U_dsdc_n154), 
	.A3(U_dsdc_n153), 
	.A2(U_dsdc_n1385), 
	.A1(U_dsdc_n2069));
   NOR2_X1 U_dsdc_U241 (.ZN(U_dsdc_n153), 
	.A2(U_dsdc_n1383), 
	.A1(U_dsdc_n1384));
   OAI21_X1 U_dsdc_U240 (.ZN(U_dsdc_n366), 
	.B2(U_dsdc_n151), 
	.B1(U_dsdc_n462), 
	.A(U_dsdc_n152));
   AOI21_X1 U_dsdc_U239 (.ZN(U_dsdc_n152), 
	.B2(U_dsdc_n462), 
	.B1(U_dsdc_n1791), 
	.A(U_dsdc_n1797));
   INV_X1 U_dsdc_U238 (.ZN(U_dsdc_n151), 
	.A(U_dsdc_n1800));
   OAI211_X1 U_dsdc_U237 (.ZN(U_dsdc_n417), 
	.C2(U_dsdc_n148), 
	.C1(U_dsdc_init_cnt_14_), 
	.B(U_dsdc_n150), 
	.A(U_dsdc_n149));
   NAND2_X1 U_dsdc_U236 (.ZN(U_dsdc_n150), 
	.A2(cr_t_init[14]), 
	.A1(U_dsdc_n1722));
   NAND3_X1 U_dsdc_U235 (.ZN(U_dsdc_n149), 
	.A3(U_dsdc_n482), 
	.A2(U_dsdc_init_cnt_14_), 
	.A1(U_dsdc_n1676));
   NAND2_X1 U_dsdc_U234 (.ZN(U_dsdc_n148), 
	.A2(U_dsdc_n147), 
	.A1(U_dsdc_n1715));
   INV_X1 U_dsdc_U233 (.ZN(U_dsdc_n147), 
	.A(U_dsdc_n482));
   AOI22_X1 U_dsdc_U232 (.ZN(U_dsdc_N4462), 
	.B2(U_dsdc_n144), 
	.B1(FE_PHN3192_U_cr_n128), 
	.A2(U_dsdc_n145), 
	.A1(U_dsdc_n313));
   AOI22_X1 U_dsdc_U230 (.ZN(U_dsdc_n145), 
	.B2(U_dsdc_n1244), 
	.B1(U_dsdc_bm_ras_cnt_3__3_), 
	.A2(FE_PHN1497_U_dsdc_n1238), 
	.A1(FE_PHN1891_U_dsdc_bm_ras_cnt_3__2_));
   AOI22_X1 U_dsdc_U229 (.ZN(U_dsdc_N4475), 
	.B2(U_dsdc_n144), 
	.B1(n96), 
	.A2(U_dsdc_n143), 
	.A1(U_dsdc_n313));
   INV_X1 U_dsdc_U228 (.ZN(U_dsdc_n144), 
	.A(U_dsdc_n313));
   AOI22_X1 U_dsdc_U227 (.ZN(U_dsdc_n143), 
	.B2(U_dsdc_n1234), 
	.B1(U_dsdc_bm_rc_cnt_3__3_), 
	.A2(U_dsdc_n1228), 
	.A1(FE_PHN1219_U_dsdc_bm_rc_cnt_3__2_));
   OAI211_X1 U_dsdc_U226 (.ZN(U_dsdc_n288), 
	.C2(U_dsdc_n139), 
	.C1(U_dsdc_n1382), 
	.B(U_dsdc_n142), 
	.A(U_dsdc_n140));
   OAI211_X1 U_dsdc_U225 (.ZN(U_dsdc_n142), 
	.C2(U_dsdc_DP_OP_1642_126_2028_n7), 
	.C1(U_dsdc_DP_OP_1642_126_2028_n15), 
	.B(U_dsdc_n141), 
	.A(U_dsdc_n1380));
   NAND2_X1 U_dsdc_U224 (.ZN(U_dsdc_n141), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n7), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n15));
   NAND2_X1 U_dsdc_U223 (.ZN(U_dsdc_n140), 
	.A2(U_dsdc_N1764), 
	.A1(U_dsdc_n1381));
   AOI21_X1 U_dsdc_U222 (.ZN(U_dsdc_n139), 
	.B2(U_dsdc_data_cnt_2_), 
	.B1(FE_PHN773_U_dsdc_n1823), 
	.A(U_dsdc_n1822));
   OAI21_X1 U_dsdc_U221 (.ZN(U_dsdc_n1354), 
	.B2(debug_ref_req), 
	.B1(U_dsdc_n1473), 
	.A(U_dsdc_n1038));
   NOR4_X1 U_dsdc_U219 (.ZN(U_dsdc_n1590), 
	.A4(U_dsdc_n137), 
	.A3(U_dsdc_n1580), 
	.A2(U_dsdc_n1667), 
	.A1(U_dsdc_n1581));
   NAND3_X1 U_dsdc_U218 (.ZN(U_dsdc_n137), 
	.A3(U_dsdc_n92), 
	.A2(U_dsdc_n1578), 
	.A1(U_dsdc_n1579));
   OR3_X1 U_dsdc_U216 (.ZN(U_dsdc_n613), 
	.A3(U_dsdc_N4239), 
	.A2(U_dsdc_N4240), 
	.A1(U_dsdc_N4241));
   OAI21_X1 U_dsdc_U213 (.ZN(U_dsdc_n982), 
	.B2(U_dsdc_n385), 
	.B1(cr_num_open_banks[4]), 
	.A(U_dsdc_n134));
   OAI221_X1 U_dsdc_U212 (.ZN(U_dsdc_n134), 
	.C2(n92), 
	.C1(U_dsdc_n131), 
	.B2(U_dsdc_bm_num_open_bank_3_), 
	.B1(U_dsdc_n131), 
	.A(U_dsdc_n133));
   AOI22_X1 U_dsdc_U211 (.ZN(U_dsdc_n133), 
	.B2(U_dsdc_n179), 
	.B1(cr_num_open_banks[3]), 
	.A2(U_dsdc_n385), 
	.A1(cr_num_open_banks[4]));
   AOI21_X1 U_dsdc_U209 (.ZN(U_dsdc_n131), 
	.B2(cr_num_open_banks[2]), 
	.B1(U_dsdc_n338), 
	.A(U_dsdc_n130));
   NOR2_X1 U_dsdc_U208 (.ZN(U_dsdc_n130), 
	.A2(U_dsdc_n129), 
	.A1(U_dsdc_n128));
   AOI22_X1 U_dsdc_U207 (.ZN(U_dsdc_n129), 
	.B2(cr_num_open_banks[0]), 
	.B1(FE_PHN1093_U_dsdc_n340), 
	.A2(U_dsdc_n180), 
	.A1(cr_num_open_banks[1]));
   OAI22_X1 U_dsdc_U206 (.ZN(U_dsdc_n128), 
	.B2(U_dsdc_n180), 
	.B1(cr_num_open_banks[1]), 
	.A2(U_dsdc_n338), 
	.A1(cr_num_open_banks[2]));
   NAND3_X1 U_dsdc_U204 (.ZN(U_dsdc_n496), 
	.A3(U_dsdc_n126), 
	.A2(U_dsdc_n493), 
	.A1(U_dsdc_n125));
   AOI22_X1 U_dsdc_U203 (.ZN(U_dsdc_n126), 
	.B2(U_dsdc_bm_row_addr_0__3_), 
	.B1(U_dsdc_n801), 
	.A2(U_dsdc_bm_row_addr_0__7_), 
	.A1(U_dsdc_n816));
   AOI21_X1 U_dsdc_U202 (.ZN(U_dsdc_n125), 
	.B2(U_dsdc_n803), 
	.B1(U_dsdc_bm_row_addr_0__9_), 
	.A(U_dsdc_n572));
   OAI211_X1 U_dsdc_U201 (.ZN(U_dsdc_n286), 
	.C2(U_dsdc_n120), 
	.C1(U_dsdc_n1382), 
	.B(U_dsdc_n124), 
	.A(U_dsdc_n121));
   OAI221_X1 U_dsdc_U200 (.ZN(U_dsdc_n124), 
	.C2(U_dsdc_DP_OP_1642_126_2028_n11), 
	.C1(U_dsdc_n123), 
	.B2(U_dsdc_n25), 
	.B1(U_dsdc_DP_OP_1642_126_2028_n28), 
	.A(U_dsdc_n1380));
   INV_X1 U_dsdc_U199 (.ZN(U_dsdc_n123), 
	.A(U_dsdc_DP_OP_1642_126_2028_n28));
   NAND2_X1 U_dsdc_U197 (.ZN(U_dsdc_n121), 
	.A2(U_dsdc_n1381), 
	.A1(U_dsdc_N1762));
   AOI21_X1 U_dsdc_U196 (.ZN(U_dsdc_n120), 
	.B2(U_dsdc_n1444), 
	.B1(U_dsdc_data_cnt_0_), 
	.A(U_dsdc_n1825));
   AOI22_X1 U_dsdc_U185 (.ZN(U_dsdc_N4415), 
	.B2(U_dsdc_n108), 
	.B1(FE_PHN3192_U_cr_n128), 
	.A2(U_dsdc_n109), 
	.A1(U_dsdc_n310));
   AOI22_X1 U_dsdc_U183 (.ZN(U_dsdc_n109), 
	.B2(U_dsdc_n1214), 
	.B1(U_dsdc_bm_ras_cnt_2__3_), 
	.A2(FE_PHN1155_U_dsdc_n1210), 
	.A1(U_dsdc_bm_ras_cnt_2__2_));
   AOI22_X1 U_dsdc_U182 (.ZN(U_dsdc_N4428), 
	.B2(U_dsdc_n108), 
	.B1(n96), 
	.A2(U_dsdc_n107), 
	.A1(U_dsdc_n310));
   INV_X1 U_dsdc_U181 (.ZN(U_dsdc_n108), 
	.A(U_dsdc_n310));
   AOI22_X1 U_dsdc_U180 (.ZN(U_dsdc_n107), 
	.B2(U_dsdc_n1207), 
	.B1(U_dsdc_bm_rc_cnt_2__3_), 
	.A2(U_dsdc_n1203), 
	.A1(FE_PHN1222_U_dsdc_bm_rc_cnt_2__2_));
   OAI21_X1 U_dsdc_U179 (.ZN(U_dsdc_N4141), 
	.B2(U_dsdc_n105), 
	.B1(U_dsdc_n1166), 
	.A(U_dsdc_n106));
   NAND2_X1 U_dsdc_U178 (.ZN(U_dsdc_n106), 
	.A2(U_dsdc_n1166), 
	.A1(cr_t_rcd[2]));
   NAND2_X1 U_dsdc_U177 (.ZN(U_dsdc_n105), 
	.A2(U_dsdc_rcd_cnt_2_), 
	.A1(U_dsdc_n1165));
   OAI21_X1 U_dsdc_U172 (.ZN(U_dsdc_N4129), 
	.B2(U_dsdc_n1393), 
	.B1(FE_PHN788_U_dsdc_n554), 
	.A(U_dsdc_n101));
   NAND3_X1 U_dsdc_U171 (.ZN(U_dsdc_n101), 
	.A3(FE_PHN1153_U_dsdc_cas_latency_cnt_3_), 
	.A2(FE_PHN1585_U_dsdc_n1094), 
	.A1(U_dsdc_n1393));
   AOI22_X1 U_dsdc_U170 (.ZN(U_dsdc_n231), 
	.B2(U_dsdc_n100), 
	.B1(U_dsdc_n98), 
	.A2(U_dsdc_n434), 
	.A1(U_dsdc_n99));
   NOR2_X1 U_dsdc_U169 (.ZN(U_dsdc_n100), 
	.A2(U_dsdc_n1971), 
	.A1(U_dsdc_n434));
   NAND2_X1 U_dsdc_U168 (.ZN(U_dsdc_n99), 
	.A2(U_dsdc_n1973), 
	.A1(U_dsdc_bm_bank_age_0__3_));
   AOI22_X1 U_dsdc_U167 (.ZN(U_dsdc_n98), 
	.B2(U_dsdc_n458), 
	.B1(U_dsdc_n1972), 
	.A2(U_dsdc_n2081), 
	.A1(U_dsdc_bm_bank_age_0__3_));
   NOR3_X1 U_dsdc_U160 (.ZN(U_dsdc_n325), 
	.A3(U_dsdc_n92), 
	.A2(U_dsdc_row_cnt_0_), 
	.A1(U_dsdc_row_cnt_1_));
   INV_X1 U_dsdc_U159 (.ZN(U_dsdc_n92), 
	.A(U_dsdc_n1791));
   XNOR2_X1 U_dsdc_U156 (.ZN(U_dsdc_N1767), 
	.B(hiu_burst_size[5]), 
	.A(U_dsdc_n90));
   AOI22_X1 U_dsdc_U155 (.ZN(U_dsdc_n90), 
	.B2(U_dsdc_DP_OP_1642_126_2028_n34), 
	.B1(U_dsdc_DP_OP_1642_126_2028_n42), 
	.A2(U_dsdc_N1991), 
	.A1(hiu_burst_size[4]));
   AOI21_X1 U_dsdc_U154 (.ZN(U_dsdc_n514), 
	.B2(U_dsdc_n801), 
	.B1(U_dsdc_n798), 
	.A(U_dsdc_n89));
   NOR3_X1 U_dsdc_U153 (.ZN(U_dsdc_n89), 
	.A3(U_dsdc_bm_row_addr_0__13_), 
	.A2(U_dsdc_n785), 
	.A1(U_dsdc_n800));
   AOI21_X2 U_dsdc_U152 (.ZN(U_dsdc_n548), 
	.B2(U_dsdc_n159), 
	.B1(U_dsdc_bm_row_addr_2__14_), 
	.A(U_dsdc_n88));
   NAND2_X2 U_dsdc_U151 (.ZN(U_dsdc_n88), 
	.A2(U_dsdc_n87), 
	.A1(U_dsdc_n547));
   AOI22_X2 U_dsdc_U150 (.ZN(U_dsdc_n87), 
	.B2(U_dsdc_bm_row_addr_1__14_), 
	.B1(U_dsdc_n604), 
	.A2(U_dsdc_bm_row_addr_0__14_), 
	.A1(U_dsdc_n998));
   AND2_X4 U_dsdc_U149 (.ZN(U_dsdc_n813), 
	.A2(U_dsdc_n86), 
	.A1(U_dsdc_n799));
   AOI22_X1 U_dsdc_U148 (.ZN(U_dsdc_n86), 
	.B2(U_dsdc_n604), 
	.B1(U_dsdc_bm_row_addr_1__1_), 
	.A2(U_dsdc_n978), 
	.A1(U_dsdc_bm_row_addr_3__1_));
   AOI221_X1 U_dsdc_U147 (.ZN(U_dsdc_cas_cnt_nxt[1]), 
	.C2(U_dsdc_n1282), 
	.C1(FE_PHN1335_U_dsdc_n1281), 
	.B2(U_dsdc_n1282), 
	.B1(FE_PHN1161_U_dsdc_n1339), 
	.A(U_dsdc_n1340));
   AOI22_X1 U_dsdc_U146 (.ZN(U_dsdc_N4368), 
	.B2(U_dsdc_n621), 
	.B1(FE_PHN3192_U_cr_n128), 
	.A2(U_dsdc_n84), 
	.A1(U_dsdc_n620));
   AOI22_X1 U_dsdc_U144 (.ZN(U_dsdc_n84), 
	.B2(U_dsdc_n1200), 
	.B1(U_dsdc_bm_ras_cnt_1__3_), 
	.A2(FE_PHN1154_U_dsdc_n1196), 
	.A1(FE_PHN1889_U_dsdc_bm_ras_cnt_1__2_));
   AOI22_X1 U_dsdc_U143 (.ZN(U_dsdc_N4381), 
	.B2(U_dsdc_n621), 
	.B1(n96), 
	.A2(U_dsdc_n82), 
	.A1(U_dsdc_n620));
   AOI22_X1 U_dsdc_U141 (.ZN(U_dsdc_n82), 
	.B2(U_dsdc_n1193), 
	.B1(U_dsdc_bm_rc_cnt_1__3_), 
	.A2(U_dsdc_n1189), 
	.A1(FE_PHN1221_U_dsdc_bm_rc_cnt_1__2_));
   OAI21_X1 U_dsdc_U140 (.ZN(U_dsdc_N4284), 
	.B2(U_dsdc_n80), 
	.B1(U_dsdc_n1166), 
	.A(U_dsdc_n81));
   NAND2_X1 U_dsdc_U139 (.ZN(U_dsdc_n81), 
	.A2(U_dsdc_n1166), 
	.A1(cr_t_ras_min[3]));
   NAND2_X1 U_dsdc_U138 (.ZN(U_dsdc_n80), 
	.A2(FE_PHN841_U_dsdc_bm_ras_cnt_max_3_), 
	.A1(FE_PHN1200_U_dsdc_n1161));
   OAI211_X1 U_dsdc_U131 (.ZN(U_dsdc_n290), 
	.C2(U_dsdc_n72), 
	.C1(U_dsdc_n1382), 
	.B(U_dsdc_n75), 
	.A(U_dsdc_n73));
   OAI211_X1 U_dsdc_U130 (.ZN(U_dsdc_n75), 
	.C2(U_dsdc_DP_OP_1642_126_2028_n13), 
	.C1(U_dsdc_DP_OP_1642_126_2028_n3), 
	.B(U_dsdc_n74), 
	.A(U_dsdc_n1380));
   NAND2_X1 U_dsdc_U129 (.ZN(U_dsdc_n74), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n13), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n3));
   NAND2_X1 U_dsdc_U128 (.ZN(U_dsdc_n73), 
	.A2(U_dsdc_N1766), 
	.A1(U_dsdc_n1381));
   AOI21_X1 U_dsdc_U127 (.ZN(U_dsdc_n72), 
	.B2(U_dsdc_n1820), 
	.B1(U_dsdc_data_cnt_4_), 
	.A(U_dsdc_n762));
   NOR2_X1 U_dsdc_U126 (.ZN(U_dsdc_n972), 
	.A2(U_dsdc_n945), 
	.A1(U_dsdc_n71));
   AOI211_X1 U_dsdc_U125 (.ZN(U_dsdc_n71), 
	.C2(U_dsdc_n1428), 
	.C1(U_dsdc_n1041), 
	.B(debug_ref_req), 
	.A(U_dsdc_n2014));
   INV_X1 U_dsdc_U124 (.ZN(U_dsdc_n494), 
	.A(U_dsdc_n70));
   AOI22_X1 U_dsdc_U123 (.ZN(U_dsdc_n70), 
	.B2(U_dsdc_bm_row_addr_0__1_), 
	.B1(U_dsdc_n814), 
	.A2(U_dsdc_bm_row_addr_0__13_), 
	.A1(U_dsdc_n800));
   AOI22_X1 U_dsdc_U122 (.ZN(U_dsdc_n515), 
	.B2(U_dsdc_bm_row_addr_0__12_), 
	.B1(U_dsdc_n998), 
	.A2(U_dsdc_bm_row_addr_1__12_), 
	.A1(U_dsdc_n604));
   OAI211_X1 U_dsdc_U121 (.ZN(U_dsdc_term_cnt_nxt[4]), 
	.C2(U_dsdc_n63), 
	.C1(U_dsdc_n457), 
	.B(U_dsdc_n69), 
	.A(U_dsdc_n66));
   OAI211_X1 U_dsdc_U120 (.ZN(U_dsdc_n69), 
	.C2(U_dsdc_n67), 
	.C1(U_dsdc_N1991), 
	.B(U_dsdc_n68), 
	.A(U_dsdc_n1379));
   NAND2_X1 U_dsdc_U119 (.ZN(U_dsdc_n68), 
	.A2(U_dsdc_n67), 
	.A1(U_dsdc_N1991));
   AND2_X1 U_dsdc_U118 (.ZN(U_dsdc_n67), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n30), 
	.A1(U_dsdc_N1990));
   AOI222_X1 U_dsdc_U117 (.ZN(U_dsdc_n66), 
	.C2(U_dsdc_n1648), 
	.C1(U_dsdc_n1424), 
	.B2(U_dsdc_n1649), 
	.B1(U_dsdc_n65), 
	.A2(U_dsdc_N1991), 
	.A1(n89));
   NOR3_X1 U_dsdc_U116 (.ZN(U_dsdc_n65), 
	.A3(U_dsdc_term_cnt_2_), 
	.A2(U_dsdc_term_cnt_4_), 
	.A1(U_dsdc_term_cnt_3_));
   AOI21_X1 U_dsdc_U114 (.ZN(U_dsdc_n63), 
	.B2(U_dsdc_n62), 
	.B1(U_dsdc_term_cnt_3_), 
	.A(U_dsdc_n1647));
   INV_X1 U_dsdc_U113 (.ZN(U_dsdc_n62), 
	.A(U_dsdc_n1646));
   AOI22_X1 U_dsdc_U112 (.ZN(U_dsdc_N4321), 
	.B2(U_dsdc_n59), 
	.B1(FE_PHN3192_U_cr_n128), 
	.A2(U_dsdc_n60), 
	.A1(n83));
   AOI22_X1 U_dsdc_U110 (.ZN(U_dsdc_n60), 
	.B2(U_dsdc_n1186), 
	.B1(U_dsdc_bm_ras_cnt_0__3_), 
	.A2(FE_PHN1156_U_dsdc_n1182), 
	.A1(U_dsdc_bm_ras_cnt_0__2_));
   AOI22_X1 U_dsdc_U109 (.ZN(U_dsdc_N4334), 
	.B2(U_dsdc_n59), 
	.B1(n96), 
	.A2(U_dsdc_n58), 
	.A1(n83));
   INV_X1 U_dsdc_U108 (.ZN(U_dsdc_n59), 
	.A(n83));
   AOI22_X1 U_dsdc_U107 (.ZN(U_dsdc_n58), 
	.B2(U_dsdc_n1179), 
	.B1(U_dsdc_bm_rc_cnt_0__3_), 
	.A2(FE_PHN945_U_dsdc_n1175), 
	.A1(U_dsdc_bm_rc_cnt_0__2_));
   XOR2_X1 U_dsdc_U100 (.Z(U_dsdc_n1085), 
	.B(FE_PHN955_s_read_pipe_1_), 
	.A(FE_PHN1402_U_dsdc_n1462));
   OR4_X1 U_dsdc_U99 (.ZN(U_dsdc_n1483), 
	.A4(U_dsdc_bm_bank_status_0_), 
	.A3(FE_PHN1593_U_dsdc_bm_bank_status_1_), 
	.A2(U_dsdc_bm_bank_status_2_), 
	.A1(U_dsdc_bm_bank_status_3_));
   AOI222_X1 U_dsdc_U98 (.ZN(U_dsdc_n1281), 
	.C2(U_dsdc_n1270), 
	.C1(hiu_burst_size[1]), 
	.B2(U_dsdc_n1269), 
	.B1(FE_PHN1896_U_dsdc_r_burst_size_1_), 
	.A2(U_dsdc_n1268), 
	.A1(U_dsdc_cas_cnt_1_));
   NOR3_X2 U_dsdc_U97 (.ZN(U_dsdc_n740), 
	.A3(U_dsdc_n53), 
	.A2(U_dsdc_data_cnt_1_), 
	.A1(U_dsdc_data_cnt_0_));
   OR4_X1 U_dsdc_U96 (.ZN(U_dsdc_n53), 
	.A4(U_dsdc_data_cnt_4_), 
	.A3(U_dsdc_data_cnt_2_), 
	.A2(U_dsdc_data_cnt_3_), 
	.A1(U_dsdc_data_cnt_5_));
   INV_X1 U_dsdc_U95 (.ZN(U_dsdc_n477), 
	.A(U_dsdc_n52));
   AOI222_X1 U_dsdc_U94 (.ZN(U_dsdc_n52), 
	.C2(U_dsdc_n476), 
	.C1(U_dsdc_bm_bank_age_3__2_), 
	.B2(U_dsdc_n1839), 
	.B1(U_dsdc_bm_bank_age_1__2_), 
	.A2(U_dsdc_bm_bank_age_2__2_), 
	.A1(U_dsdc_n1840));
   AOI22_X2 U_dsdc_U92 (.ZN(U_dsdc_n51), 
	.B2(U_dsdc_n802), 
	.B1(debug_ad_row_addr[9]), 
	.A2(U_dsdc_n805), 
	.A1(debug_ad_row_addr[15]));
   AOI22_X1 U_dsdc_U91 (.ZN(U_dsdc_n562), 
	.B2(U_dsdc_bm_row_addr_0__2_), 
	.B1(U_dsdc_n998), 
	.A2(U_dsdc_bm_row_addr_1__2_), 
	.A1(U_dsdc_n604));
   OAI21_X1 U_dsdc_U87 (.ZN(U_dsdc_term_cnt_nxt[2]), 
	.B2(U_dsdc_n200), 
	.B1(U_dsdc_n1643), 
	.A(U_dsdc_n48));
   AOI21_X1 U_dsdc_U86 (.ZN(U_dsdc_n48), 
	.B2(n89), 
	.B1(U_dsdc_N1989), 
	.A(U_dsdc_n47));
   OAI21_X1 U_dsdc_U85 (.ZN(U_dsdc_n47), 
	.B2(U_dsdc_term_cnt_2_), 
	.B1(U_dsdc_n1645), 
	.A(U_dsdc_n46));
   AOI22_X1 U_dsdc_U84 (.ZN(U_dsdc_n46), 
	.B2(U_dsdc_n45), 
	.B1(U_dsdc_n1379), 
	.A2(U_dsdc_n770), 
	.A1(U_dsdc_r_cas_latency_2_));
   XOR2_X1 U_dsdc_U83 (.Z(U_dsdc_n45), 
	.B(U_dsdc_DP_OP_1642_126_2028_n31), 
	.A(U_dsdc_N1989));
   INV_X4 U_dsdc_U82 (.ZN(U_dsdc_n291), 
	.A(U_dsdc_n44));
   AOI222_X1 U_dsdc_U81 (.ZN(U_dsdc_n44), 
	.C2(U_dsdc_n43), 
	.C1(U_dsdc_n764), 
	.B2(U_dsdc_n1381), 
	.B1(U_dsdc_N1767), 
	.A2(U_dsdc_n1380), 
	.A1(U_dsdc_C880_DATA5_5));
   XOR2_X1 U_dsdc_U80 (.Z(U_dsdc_n43), 
	.B(U_dsdc_n762), 
	.A(U_dsdc_data_cnt_5_));
   OAI22_X1 U_dsdc_U79 (.ZN(U_dsdc_n281), 
	.B2(U_dsdc_n440), 
	.B1(U_dsdc_n42), 
	.A2(U_dsdc_n41), 
	.A1(U_dsdc_n2073));
   AND3_X1 U_dsdc_U78 (.ZN(U_dsdc_n42), 
	.A3(U_dsdc_n2075), 
	.A2(U_dsdc_n2071), 
	.A1(U_dsdc_n2072));
   AOI221_X1 U_dsdc_U77 (.ZN(U_dsdc_n41), 
	.C2(U_dsdc_n721), 
	.C1(U_dsdc_n39), 
	.B2(U_dsdc_n721), 
	.B1(U_dsdc_n1872), 
	.A(U_dsdc_n40));
   INV_X1 U_dsdc_U76 (.ZN(U_dsdc_n40), 
	.A(U_dsdc_n974));
   NAND2_X1 U_dsdc_U75 (.ZN(U_dsdc_n39), 
	.A2(U_dsdc_n991), 
	.A1(U_dsdc_n2069));
   NAND3_X1 U_dsdc_U71 (.ZN(U_dsdc_n979), 
	.A3(U_dsdc_n35), 
	.A2(U_dsdc_n34), 
	.A1(U_dsdc_n36));
   NAND2_X1 U_dsdc_U70 (.ZN(U_dsdc_n36), 
	.A2(U_dsdc_n998), 
	.A1(U_dsdc_n1181));
   AOI22_X1 U_dsdc_U69 (.ZN(U_dsdc_n35), 
	.B2(U_dsdc_n1237), 
	.B1(U_dsdc_n978), 
	.A2(U_dsdc_n1209), 
	.A1(U_dsdc_n159));
   AOI21_X1 U_dsdc_U68 (.ZN(U_dsdc_n34), 
	.B2(U_dsdc_n604), 
	.B1(U_dsdc_n1195), 
	.A(U_dsdc_n1294));
   INV_X1 U_dsdc_U67 (.ZN(U_dsdc_n495), 
	.A(U_dsdc_n33));
   AOI22_X1 U_dsdc_U66 (.ZN(U_dsdc_n33), 
	.B2(U_dsdc_bm_row_addr_0__11_), 
	.B1(U_addrdec_n231), 
	.A2(U_dsdc_bm_row_addr_0__15_), 
	.A1(U_dsdc_n806));
   NAND3_X1 U_dsdc_U62 (.ZN(U_dsdc_term_cnt_nxt[1]), 
	.A3(U_dsdc_n30), 
	.A2(U_dsdc_n28), 
	.A1(U_dsdc_n1645));
   AOI22_X1 U_dsdc_U61 (.ZN(U_dsdc_n30), 
	.B2(n89), 
	.B1(U_dsdc_N1988), 
	.A2(U_dsdc_n29), 
	.A1(U_dsdc_term_cnt_1_));
   OAI22_X1 U_dsdc_U60 (.ZN(U_dsdc_n29), 
	.B2(U_dsdc_n463), 
	.B1(U_dsdc_n1646), 
	.A2(U_dsdc_n1636), 
	.A1(FE_PHN671_U_dsdc_n1637));
   AOI22_X1 U_dsdc_U59 (.ZN(U_dsdc_n28), 
	.B2(U_dsdc_n27), 
	.B1(U_dsdc_n1379), 
	.A2(U_dsdc_n770), 
	.A1(U_dsdc_r_cas_latency_1_));
   XOR2_X1 U_dsdc_U58 (.Z(U_dsdc_n27), 
	.B(U_dsdc_N1988), 
	.A(U_dsdc_N1987));
   INV_X1 U_dsdc_U57 (.ZN(U_dsdc_n1093), 
	.A(U_dsdc_n26));
   AOI22_X1 U_dsdc_U56 (.ZN(U_dsdc_n26), 
	.B2(FE_PHN1402_U_dsdc_n1462), 
	.B1(FE_PHN955_s_read_pipe_1_), 
	.A2(FE_PHN1020_U_dsdc_n1085), 
	.A1(FE_PHN1921_U_dsdc_n1084));
   AOI222_X1 U_dsdc_U55 (.ZN(U_dsdc_n1276), 
	.C2(U_dsdc_n1270), 
	.C1(hiu_burst_size[3]), 
	.B2(U_dsdc_n1269), 
	.B1(FE_PHN1892_U_dsdc_r_burst_size_3_), 
	.A2(U_dsdc_n1268), 
	.A1(U_dsdc_cas_cnt_3_));
   OAI22_X1 U_dsdc_U54 (.ZN(U_dsdc_n163), 
	.B2(U_dsdc_n601), 
	.B1(U_dsdc_n162), 
	.A2(U_dsdc_n25), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n28));
   INV_X1 U_dsdc_U53 (.ZN(U_dsdc_n25), 
	.A(U_dsdc_DP_OP_1642_126_2028_n11));
   NAND2_X1 U_dsdc_U52 (.ZN(U_dsdc_n716), 
	.A2(U_dsdc_n24), 
	.A1(U_dsdc_n937));
   AOI21_X1 U_dsdc_U51 (.ZN(U_dsdc_n24), 
	.B2(U_dsdc_n759), 
	.B1(U_dsdc_n672), 
	.A(U_dsdc_n683));
   AND2_X1 U_dsdc_U50 (.ZN(U_dsdc_n884), 
	.A2(U_dsdc_n23), 
	.A1(U_dsdc_n22));
   AOI22_X1 U_dsdc_U49 (.ZN(U_dsdc_n23), 
	.B2(U_dsdc_bm_bank_status_3_), 
	.B1(U_dsdc_n978), 
	.A2(U_dsdc_bm_bank_status_0_), 
	.A1(U_dsdc_n998));
   AOI22_X1 U_dsdc_U48 (.ZN(U_dsdc_n22), 
	.B2(U_dsdc_bm_bank_status_2_), 
	.B1(U_dsdc_n159), 
	.A2(FE_PHN1593_U_dsdc_bm_bank_status_1_), 
	.A1(U_dsdc_n604));
   NOR4_X1 U_dsdc_U47 (.ZN(U_dsdc_n1428), 
	.A4(cr_mode_reg_update), 
	.A3(cr_do_self_ref_rp), 
	.A2(cr_exn_mode_reg_update), 
	.A1(cr_do_initialize));
   OAI221_X1 U_dsdc_U42 (.ZN(U_dsdc_n[2090]), 
	.C2(U_dsdc_n1417), 
	.C1(U_dsdc_n355), 
	.B2(U_dsdc_n2069), 
	.B1(U_dsdc_n355), 
	.A(U_dsdc_n18));
   NOR4_X1 U_dsdc_U41 (.ZN(U_dsdc_n18), 
	.A4(U_dsdc_n17), 
	.A3(U_dsdc_n1363), 
	.A2(U_dsdc_n1412), 
	.A1(U_dsdc_n1344));
   OAI211_X1 U_dsdc_U40 (.ZN(U_dsdc_n17), 
	.C2(U_dsdc_n1805), 
	.C1(U_dsdc_n2071), 
	.B(U_dsdc_n16), 
	.A(U_dsdc_n1979));
   OR2_X1 U_dsdc_U39 (.ZN(U_dsdc_n16), 
	.A2(U_dsdc_n1496), 
	.A1(U_dsdc_n1650));
   XNOR2_X1 U_dsdc_U37 (.ZN(U_dsdc_DP_OP_1642_126_2028_n20), 
	.B(U_dsdc_DP_OP_1642_126_2028_n85), 
	.A(U_dsdc_n15));
   NAND2_X1 U_dsdc_U36 (.ZN(U_dsdc_n15), 
	.A2(U_dsdc_n753), 
	.A1(U_dsdc_r_cas_latency_2_));
   OAI211_X1 U_dsdc_U35 (.ZN(U_dsdc_n492), 
	.C2(U_dsdc_n800), 
	.C1(U_dsdc_n785), 
	.B(U_dsdc_n14), 
	.A(U_dsdc_n572));
   NAND2_X1 U_dsdc_U34 (.ZN(U_dsdc_n14), 
	.A2(debug_ad_row_addr[11]), 
	.A1(U_dsdc_n810));
   OAI211_X1 U_dsdc_U32 (.ZN(U_dsdc_term_cnt_nxt[0]), 
	.C2(U_dsdc_n8), 
	.C1(U_dsdc_term_cnt_0_), 
	.B(U_dsdc_n12), 
	.A(U_dsdc_n11));
   NAND2_X1 U_dsdc_U31 (.ZN(U_dsdc_n12), 
	.A2(n89), 
	.A1(U_dsdc_N1987));
   AOI222_X1 U_dsdc_U30 (.ZN(U_dsdc_n11), 
	.C2(U_dsdc_n770), 
	.C1(U_dsdc_r_cas_latency_0_), 
	.B2(U_dsdc_n10), 
	.B1(U_dsdc_term_cnt_0_), 
	.A2(U_dsdc_n1379), 
	.A1(U_dsdc_n9));
   NOR2_X1 U_dsdc_U29 (.ZN(U_dsdc_n10), 
	.A2(FE_PHN671_U_dsdc_n1637), 
	.A1(U_dsdc_n1636));
   INV_X1 U_dsdc_U28 (.ZN(U_dsdc_n9), 
	.A(U_dsdc_N1987));
   AOI21_X1 U_dsdc_U27 (.ZN(U_dsdc_n8), 
	.B2(U_dsdc_n1642), 
	.B1(FE_PHN671_U_dsdc_n1637), 
	.A(U_dsdc_n1639));
   NAND2_X1 U_dsdc_U26 (.ZN(U_dsdc_n1320), 
	.A2(U_dsdc_n7), 
	.A1(U_dsdc_n1043));
   NAND2_X1 U_dsdc_U25 (.ZN(U_dsdc_n7), 
	.A2(U_dsdc_n1286), 
	.A1(U_dsdc_n6));
   NAND3_X1 U_dsdc_U24 (.ZN(U_dsdc_n6), 
	.A3(U_dsdc_n1411), 
	.A2(U_dsdc_n1042), 
	.A1(U_dsdc_n1041));
   NAND3_X2 U_dsdc_U23 (.ZN(U_dsdc_n2007), 
	.A3(U_dsdc_n5), 
	.A2(U_dsdc_n717), 
	.A1(U_dsdc_n3));
   AOI211_X1 U_dsdc_U22 (.ZN(U_dsdc_n5), 
	.C2(U_dsdc_n1412), 
	.C1(U_dsdc_n1061), 
	.B(U_dsdc_n716), 
	.A(U_dsdc_n4));
   AOI21_X1 U_dsdc_U21 (.ZN(U_dsdc_n4), 
	.B2(U_dsdc_n1980), 
	.B1(U_dsdc_n181), 
	.A(U_dsdc_n1064));
   AOI21_X1 U_dsdc_U20 (.ZN(U_dsdc_n3), 
	.B2(U_dsdc_n2), 
	.B1(U_dsdc_n881), 
	.A(U_dsdc_n2012));
   INV_X1 U_dsdc_U19 (.ZN(U_dsdc_n2), 
	.A(U_dsdc_n1299));
   XNOR2_X1 U_dsdc_U18 (.ZN(U_dsdc_DP_OP_1642_126_2028_n21), 
	.B(U_dsdc_DP_OP_1642_126_2028_n85), 
	.A(U_dsdc_n1));
   NAND2_X1 U_dsdc_U17 (.ZN(U_dsdc_n1), 
	.A2(U_dsdc_n753), 
	.A1(U_dsdc_r_cas_latency_1_));
   NOR2_X2 U_dsdc_U15 (.ZN(U_dsdc_n1393), 
	.A2(U_dsdc_n1364), 
	.A1(U_dsdc_n1124));
   AOI222_X1 U_dsdc_U13 (.ZN(U_dsdc_n763), 
	.C2(U_dsdc_N1765), 
	.C1(U_dsdc_n1381), 
	.B2(U_dsdc_n764), 
	.B1(U_dsdc_n1821), 
	.A2(U_dsdc_C880_DATA5_3), 
	.A1(U_dsdc_n1380));
   AOI222_X1 U_dsdc_U12 (.ZN(U_dsdc_n765), 
	.C2(U_dsdc_N1763), 
	.C1(U_dsdc_n1381), 
	.B2(U_dsdc_n764), 
	.B1(U_dsdc_n1824), 
	.A2(U_dsdc_C880_DATA5_1), 
	.A1(U_dsdc_n1380));
   NAND2_X2 U_dsdc_U11 (.ZN(U_dsdc_n1286), 
	.A2(U_dsdc_n983), 
	.A1(U_dsdc_n900));
   INV_X4 U_dsdc_U10 (.ZN(U_dsdc_n620), 
	.A(U_dsdc_n621));
   AOI22_X2 U_dsdc_U9 (.ZN(U_dsdc_DP_OP_1642_126_2028_n8), 
	.B2(U_dsdc_DP_OP_1642_126_2028_n21), 
	.B1(U_dsdc_DP_OP_1642_126_2028_n58), 
	.A2(U_dsdc_n163), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n9));
   NAND2_X2 U_dsdc_U5 (.ZN(U_dsdc_n914), 
	.A2(U_dsdc_n818), 
	.A1(U_dsdc_n887));
   INV_X4 U_dsdc_U4 (.ZN(U_dsdc_n887), 
	.A(U_dsdc_n483));
   DFFR_X2 U_dsdc_term_cnt_reg_0_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n463), 
	.Q(U_dsdc_term_cnt_0_), 
	.D(FE_PHN740_U_dsdc_term_cnt_nxt_0_), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dsdc_r_row_addr_reg_0_ (.RN(FE_OFN50_HRESETn), 
	.QN(U_dsdc_n453), 
	.Q(U_dsdc_r_row_addr_0_), 
	.D(FE_PHN2030_U_dsdc_n255), 
	.CK(HCLK__L5_N33));
   DFFR_X2 U_dsdc_r_row_addr_reg_1_ (.RN(FE_OFN191_HRESETn), 
	.QN(U_dsdc_n452), 
	.Q(U_dsdc_r_row_addr_1_), 
	.D(FE_PHN2033_U_dsdc_n262), 
	.CK(HCLK__L5_N33));
   DFFR_X2 U_dsdc_r_row_addr_reg_2_ (.RN(FE_OFN36_HRESETn), 
	.QN(U_dsdc_n451), 
	.Q(U_dsdc_r_row_addr_2_), 
	.D(FE_PHN2029_U_dsdc_n263), 
	.CK(HCLK__L5_N29));
   DFFR_X2 U_dsdc_r_row_addr_reg_3_ (.RN(FE_OFN191_HRESETn), 
	.QN(U_dsdc_n450), 
	.Q(U_dsdc_r_row_addr_3_), 
	.D(FE_PHN2031_U_dsdc_n264), 
	.CK(HCLK__L5_N33));
   DFFR_X2 U_dsdc_r_row_addr_reg_7_ (.RN(FE_OFN50_HRESETn), 
	.QN(U_dsdc_n449), 
	.Q(U_dsdc_r_row_addr_7_), 
	.D(FE_PHN2027_U_dsdc_n268), 
	.CK(HCLK__L5_N33));
   DFFR_X2 U_dsdc_r_row_addr_reg_9_ (.RN(FE_OFN50_HRESETn), 
	.QN(U_dsdc_n448), 
	.Q(U_dsdc_r_row_addr_9_), 
	.D(FE_PHN2032_U_dsdc_n270), 
	.CK(HCLK__L5_N33));
   DFFR_X2 U_dsdc_r_row_addr_reg_11_ (.RN(FE_OFN50_HRESETn), 
	.QN(U_dsdc_n447), 
	.Q(U_dsdc_r_row_addr_11_), 
	.D(FE_PHN1269_U_dsdc_n257), 
	.CK(HCLK__L5_N29));
   DFFR_X2 U_dsdc_r_row_addr_reg_13_ (.RN(FE_OFN50_HRESETn), 
	.QN(U_dsdc_n454), 
	.Q(U_dsdc_r_row_addr_13_), 
	.D(FE_PHN1480_U_dsdc_n259), 
	.CK(HCLK__L5_N33));
   DFFR_X2 U_dsdc_r_row_addr_reg_14_ (.RN(FE_OFN50_HRESETn), 
	.QN(U_dsdc_n455), 
	.Q(U_dsdc_r_row_addr_14_), 
	.D(FE_PHN1479_U_dsdc_n260), 
	.CK(HCLK__L5_N33));
   DFFR_X2 U_dsdc_r_row_addr_reg_15_ (.RN(FE_OFN50_HRESETn), 
	.QN(U_dsdc_n456), 
	.Q(U_dsdc_r_row_addr_15_), 
	.D(FE_PHN1478_U_dsdc_n261), 
	.CK(HCLK__L5_N34));
   DFFR_X2 U_dsdc_r_burst_size_reg_3_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n299), 
	.Q(U_dsdc_r_burst_size_3_), 
	.D(FE_PHN3299_U_dsdc_n274), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_r_burst_size_reg_4_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n301), 
	.Q(U_dsdc_r_burst_size_4_), 
	.D(FE_PHN3289_U_dsdc_n275), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_r_burst_size_reg_5_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n172), 
	.Q(U_dsdc_r_burst_size_5_), 
	.D(FE_PHN3293_U_dsdc_n276), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_r_burst_size_reg_0_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n182), 
	.Q(U_dsdc_r_burst_size_0_), 
	.D(FE_PHN2040_U_dsdc_n271), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_access_cs_reg_2_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dsdc_n355), 
	.Q(U_dsdc_access_cs_2_), 
	.D(FE_PHN3105_U_dsdc_n_2090_), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dsdc_r_wrapped_burst_reg (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n328), 
	.Q(U_dsdc_r_wrapped_burst), 
	.D(FE_PHN2038_U_dsdc_n277), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_i_col_addr_reg_1_ (.RN(FE_OFN36_HRESETn), 
	.QN(U_dsdc_n354), 
	.Q(U_dsdc_i_col_addr_1_), 
	.D(FE_PHN1484_U_dsdc_n319), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_dsdc_delta_delay_reg_0_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n461), 
	.Q(U_dsdc_delta_delay_0_), 
	.D(FE_PHN951_U_dsdc_n216), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_early_term_flag_reg (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n306), 
	.Q(U_dsdc_early_term_flag), 
	.D(FE_PHN1493_U_dsdc_n282), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dsdc_data_flag_reg (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n440), 
	.Q(U_dsdc_data_flag), 
	.D(FE_PHN1016_U_dsdc_n281), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dsdc_rcar_cnt2_reg_3_ (.RN(FE_OFN142_HRESETn), 
	.QN(U_dsdc_n430), 
	.Q(U_dsdc_rcar_cnt2_3_), 
	.D(FE_PHN960_U_dsdc_rcar_cnt2_nxt_3_), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dsdc_mrd_cnt_reg_0_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_dsdc_n199), 
	.Q(U_dsdc_mrd_cnt_0_), 
	.D(FE_PHN796_U_dsdc_N4174), 
	.CK(HCLK__L5_N11));
   DFFR_X2 U_dsdc_mrd_cnt_reg_1_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_dsdc_n429), 
	.Q(U_dsdc_mrd_cnt_1_), 
	.D(FE_PHN1521_U_dsdc_n423), 
	.CK(HCLK__L5_N11));
   DFFR_X2 U_dsdc_num_init_ref_cnt_reg_2_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_dsdc_n473), 
	.Q(U_dsdc_num_init_ref_cnt_2_), 
	.D(FE_PHN1143_U_dsdc_num_init_ref_cnt_nxt_2_), 
	.CK(hclk));
   DFFR_X2 U_dsdc_rp_cnt1_reg_0_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_dsdc_n169), 
	.Q(U_dsdc_rp_cnt1_0_), 
	.D(FE_PHN1198_U_dsdc_rp_cnt1_nxt_0_), 
	.CK(HCLK__L5_N11));
   DFFR_X2 U_dsdc_rp_cnt1_reg_2_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_dsdc_n427), 
	.Q(U_dsdc_rp_cnt1_2_), 
	.D(FE_PHN1199_U_dsdc_rp_cnt1_nxt_2_), 
	.CK(HCLK__L5_N11));
   DFFR_X2 U_dsdc_rp_cnt1_reg_1_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_dsdc_n198), 
	.Q(U_dsdc_rp_cnt1_1_), 
	.D(FE_PHN1087_U_dsdc_rp_cnt1_nxt_1_), 
	.CK(HCLK__L5_N11));
   DFFR_X2 U_dsdc_r_cas_latency_reg_0_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n342), 
	.Q(U_dsdc_r_cas_latency_0_), 
	.D(FE_PHN1249_U_dsdc_add_x_2600_1_n8), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_bm_num_open_bank_reg_3_ (.RN(FE_OFN186_HRESETn), 
	.QN(U_dsdc_n179), 
	.Q(U_dsdc_bm_num_open_bank_3_), 
	.D(FE_PHN865_U_dsdc_n296), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_dsdc_operation_cs_reg_3_ (.RN(FE_OFN142_HRESETn), 
	.QN(U_dsdc_n196), 
	.Q(U_dsdc_operation_cs_3_), 
	.D(FE_PHN931_U_dsdc_n2094), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dsdc_row_cnt_reg_12_ (.RN(FE_OFN186_HRESETn), 
	.QN(U_dsdc_n203), 
	.Q(U_dsdc_row_cnt_12_), 
	.D(FE_PHN1120_U_dsdc_n369), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_dsdc_bm_bank_age_reg_0__0_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n201), 
	.Q(U_dsdc_bm_bank_age_0__0_), 
	.D(FE_PHN895_U_dsdc_n283), 
	.CK(HCLK__L5_N30));
   DFFR_X2 U_dsdc_bm_bank_age_reg_2__2_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n336), 
	.Q(U_dsdc_bm_bank_age_2__2_), 
	.D(FE_PHN863_U_dsdc_n211), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_data_cnt_reg_1_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n436), 
	.Q(U_dsdc_data_cnt_1_), 
	.D(FE_PHN836_U_dsdc_n287), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_bm_bank_age_reg_2__0_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n353), 
	.Q(U_dsdc_bm_bank_age_2__0_), 
	.D(FE_PHN992_U_dsdc_n209), 
	.CK(HCLK__L5_N30));
   DFFR_X2 U_dsdc_bm_bank_age_reg_1__0_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n352), 
	.Q(U_dsdc_bm_bank_age_1__0_), 
	.D(FE_PHN917_U_dsdc_n223), 
	.CK(HCLK__L5_N30));
   DFFR_X2 U_dsdc_wrapped_pop_flag_reg (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_wrapped_pop_flag), 
	.D(FE_PHN1144_U_dsdc_wrapped_pop_flag_nxt), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_num_init_ref_cnt_reg_0_ (.RN(FE_OFN63_HRESETn), 
	.Q(U_dsdc_num_init_ref_cnt_0_), 
	.D(FE_PHN996_U_dsdc_num_init_ref_cnt_nxt_0_), 
	.CK(hclk));
   DFFR_X2 U_dsdc_num_init_ref_cnt_reg_1_ (.RN(FE_OFN63_HRESETn), 
	.Q(U_dsdc_num_init_ref_cnt_1_), 
	.D(FE_PHN797_U_dsdc_num_init_ref_cnt_nxt_1_), 
	.CK(hclk));
   DFFR_X2 U_dsdc_rp_cnt2_reg_0_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_dsdc_n171), 
	.D(FE_PHN1054_U_dsdc_rp_cnt2_nxt_0_), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_dsdc_write_start_reg (.RN(FE_OFN39_HRESETn), 
	.QN(U_dsdc_n433), 
	.D(FE_PHN1470_U_dsdc_write_start_nxt), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_dsdc_rcd_cnt_reg_1_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_dsdc_n326), 
	.D(FE_PHN1491_U_dsdc_N4140), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_dsdc_wtr_cnt_reg_1_ (.RN(FE_OFN142_HRESETn), 
	.QN(U_dsdc_n194), 
	.D(FE_PHN1242_U_dsdc_wtr_cnt_nxt_1_), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dsdc_cas_cnt_reg_0_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n327), 
	.D(U_dsdc_cas_cnt_nxt[0]), 
	.CK(HCLK__L5_N31));
   DFFR_X2 U_dsdc_xsr_cnt_reg_6_ (.RN(FE_OFN142_HRESETn), 
	.QN(U_dsdc_n359), 
	.D(FE_PHN1095_U_dsdc_n392), 
	.CK(hclk));
   DFFR_X2 U_dsdc_terminate_reg (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n181), 
	.Q(U_dsdc_n165), 
	.D(hiu_terminate), 
	.CK(HCLK__L5_N28));
   XOR2_X1 U_dsdc_DP_OP_1642_126_2028_U42 (.Z(U_dsdc_N2002), 
	.B(U_dsdc_N1990), 
	.A(U_dsdc_DP_OP_1642_126_2028_n30));
   AND2_X2 U_dsdc_DP_OP_1642_126_2028_U45 (.ZN(U_dsdc_DP_OP_1642_126_2028_n30), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n31), 
	.A1(U_dsdc_N1989));
   AND2_X2 U_dsdc_DP_OP_1642_126_2028_U47 (.ZN(U_dsdc_DP_OP_1642_126_2028_n31), 
	.A2(U_dsdc_N1987), 
	.A1(U_dsdc_N1988));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U1 (.Z(U_dsdc_C880_DATA5_5), 
	.B(U_dsdc_DP_OP_1642_126_2028_n12), 
	.A(U_dsdc_DP_OP_1642_126_2028_n1));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U2 (.Z(U_dsdc_DP_OP_1642_126_2028_n1), 
	.B(U_dsdc_DP_OP_1642_126_2028_n62), 
	.A(U_dsdc_DP_OP_1642_126_2028_n85));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U6 (.Z(U_dsdc_DP_OP_1642_126_2028_n3), 
	.B(U_dsdc_DP_OP_1642_126_2028_n61), 
	.A(U_dsdc_DP_OP_1642_126_2028_n85));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U7 (.Z(U_dsdc_C880_DATA5_3), 
	.B(U_dsdc_DP_OP_1642_126_2028_n5), 
	.A(U_dsdc_DP_OP_1642_126_2028_n14));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U10 (.Z(U_dsdc_DP_OP_1642_126_2028_n5), 
	.B(U_dsdc_DP_OP_1642_126_2028_n60), 
	.A(U_dsdc_DP_OP_1642_126_2028_n19));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U14 (.Z(U_dsdc_DP_OP_1642_126_2028_n7), 
	.B(U_dsdc_DP_OP_1642_126_2028_n59), 
	.A(U_dsdc_DP_OP_1642_126_2028_n20));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U15 (.Z(U_dsdc_C880_DATA5_1), 
	.B(U_dsdc_DP_OP_1642_126_2028_n9), 
	.A(U_dsdc_n163));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U18 (.Z(U_dsdc_DP_OP_1642_126_2028_n9), 
	.B(U_dsdc_DP_OP_1642_126_2028_n58), 
	.A(U_dsdc_DP_OP_1642_126_2028_n21));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U51 (.Z(U_dsdc_N1766), 
	.B(U_dsdc_DP_OP_1642_126_2028_n42), 
	.A(U_dsdc_DP_OP_1642_126_2028_n34));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U54 (.Z(U_dsdc_DP_OP_1642_126_2028_n34), 
	.B(U_dsdc_N1991), 
	.A(hiu_burst_size[4]));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U55 (.Z(U_dsdc_N1765), 
	.B(U_dsdc_DP_OP_1642_126_2028_n43), 
	.A(U_dsdc_DP_OP_1642_126_2028_n36));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U58 (.Z(U_dsdc_DP_OP_1642_126_2028_n36), 
	.B(U_dsdc_N1990), 
	.A(hiu_burst_size[3]));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U59 (.Z(U_dsdc_N1764), 
	.B(U_dsdc_DP_OP_1642_126_2028_n38), 
	.A(U_dsdc_DP_OP_1642_126_2028_n44));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U62 (.Z(U_dsdc_DP_OP_1642_126_2028_n38), 
	.B(U_dsdc_N1989), 
	.A(hiu_burst_size[2]));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U63 (.Z(U_dsdc_N1763), 
	.B(U_dsdc_DP_OP_1642_126_2028_n40), 
	.A(U_dsdc_DP_OP_1642_126_2028_n45));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U66 (.Z(U_dsdc_DP_OP_1642_126_2028_n40), 
	.B(U_dsdc_N1988), 
	.A(hiu_burst_size[1]));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U67 (.Z(U_dsdc_N1762), 
	.B(U_dsdc_N1987), 
	.A(hiu_burst_size[0]));
   AND2_X4 U_dsdc_DP_OP_1642_126_2028_U68 (.ZN(U_dsdc_DP_OP_1642_126_2028_n45), 
	.A2(hiu_burst_size[0]), 
	.A1(U_dsdc_N1987));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U69 (.Z(U_dsdc_N1990), 
	.B(U_dsdc_DP_OP_1642_126_2028_n50), 
	.A(U_dsdc_r_cas_latency_3_));
   AND2_X4 U_dsdc_DP_OP_1642_126_2028_U70 (.ZN(U_dsdc_N1991), 
	.A2(U_dsdc_r_cas_latency_3_), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n50));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U71 (.Z(U_dsdc_N1989), 
	.B(U_dsdc_DP_OP_1642_126_2028_n51), 
	.A(U_dsdc_DP_OP_1642_126_2028_n47));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U74 (.Z(U_dsdc_DP_OP_1642_126_2028_n47), 
	.B(U_dsdc_r_cas_latency_2_), 
	.A(U_dsdc_delta_delay_2_));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U75 (.Z(U_dsdc_N1988), 
	.B(U_dsdc_DP_OP_1642_126_2028_n49), 
	.A(U_dsdc_DP_OP_1642_126_2028_n52));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U78 (.Z(U_dsdc_DP_OP_1642_126_2028_n49), 
	.B(U_dsdc_r_cas_latency_1_), 
	.A(U_dsdc_delta_delay_1_));
   XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U79 (.Z(U_dsdc_N1987), 
	.B(U_dsdc_r_cas_latency_0_), 
	.A(U_dsdc_delta_delay_0_));
   AND2_X4 U_dsdc_DP_OP_1642_126_2028_U80 (.ZN(U_dsdc_DP_OP_1642_126_2028_n52), 
	.A2(U_dsdc_delta_delay_0_), 
	.A1(U_dsdc_r_cas_latency_0_));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U77 (.ZN(U_dsdc_DP_OP_1642_126_2028_n48), 
	.B2(U_dsdc_delta_delay_1_), 
	.B1(U_dsdc_r_cas_latency_1_), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n52), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n49));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U76 (.ZN(U_dsdc_DP_OP_1642_126_2028_n51), 
	.A(U_dsdc_DP_OP_1642_126_2028_n48));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U65 (.ZN(U_dsdc_DP_OP_1642_126_2028_n39), 
	.B2(hiu_burst_size[1]), 
	.B1(U_dsdc_N1988), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n45), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n40));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U64 (.ZN(U_dsdc_DP_OP_1642_126_2028_n44), 
	.A(U_dsdc_DP_OP_1642_126_2028_n39));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U61 (.ZN(U_dsdc_DP_OP_1642_126_2028_n37), 
	.B2(hiu_burst_size[2]), 
	.B1(U_dsdc_N1989), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n44), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n38));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U60 (.ZN(U_dsdc_DP_OP_1642_126_2028_n43), 
	.A(U_dsdc_DP_OP_1642_126_2028_n37));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U73 (.ZN(U_dsdc_DP_OP_1642_126_2028_n46), 
	.B2(U_dsdc_delta_delay_2_), 
	.B1(U_dsdc_r_cas_latency_2_), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n47), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n51));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U72 (.ZN(U_dsdc_DP_OP_1642_126_2028_n50), 
	.A(U_dsdc_DP_OP_1642_126_2028_n46));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U57 (.ZN(U_dsdc_DP_OP_1642_126_2028_n35), 
	.B2(hiu_burst_size[3]), 
	.B1(U_dsdc_N1990), 
	.A2(U_dsdc_DP_OP_1642_126_2028_n36), 
	.A1(U_dsdc_DP_OP_1642_126_2028_n43));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U56 (.ZN(U_dsdc_DP_OP_1642_126_2028_n42), 
	.A(U_dsdc_DP_OP_1642_126_2028_n35));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U29 (.ZN(U_dsdc_DP_OP_1642_126_2028_n23), 
	.B2(U_dsdc_DP_OP_1642_126_2028_I5_5_), 
	.B1(U_dsdc_DP_OP_1642_126_2028_I6), 
	.A2(U_dsdc_DP_OP_1642_126_2028_I4), 
	.A1(U_dsdc_N1767));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U30 (.ZN(U_dsdc_DP_OP_1642_126_2028_n62), 
	.A(U_dsdc_DP_OP_1642_126_2028_n23));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U34 (.ZN(U_dsdc_DP_OP_1642_126_2028_n25), 
	.B2(U_dsdc_DP_OP_1642_126_2028_I5_3_), 
	.B1(U_dsdc_DP_OP_1642_126_2028_I6), 
	.A2(U_dsdc_DP_OP_1642_126_2028_I4), 
	.A1(U_dsdc_N1765));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U33 (.ZN(U_dsdc_DP_OP_1642_126_2028_n60), 
	.A(U_dsdc_DP_OP_1642_126_2028_n25));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U36 (.ZN(U_dsdc_DP_OP_1642_126_2028_n26), 
	.B2(U_dsdc_DP_OP_1642_126_2028_I5_2_), 
	.B1(U_dsdc_DP_OP_1642_126_2028_I6), 
	.A2(U_dsdc_DP_OP_1642_126_2028_I4), 
	.A1(U_dsdc_N1764));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U35 (.ZN(U_dsdc_DP_OP_1642_126_2028_n59), 
	.A(U_dsdc_DP_OP_1642_126_2028_n26));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U38 (.ZN(U_dsdc_DP_OP_1642_126_2028_n27), 
	.B2(U_dsdc_DP_OP_1642_126_2028_I5_1_), 
	.B1(U_dsdc_DP_OP_1642_126_2028_I6), 
	.A2(U_dsdc_DP_OP_1642_126_2028_I4), 
	.A1(U_dsdc_N1763));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U37 (.ZN(U_dsdc_DP_OP_1642_126_2028_n58), 
	.A(U_dsdc_DP_OP_1642_126_2028_n27));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U40 (.ZN(U_dsdc_DP_OP_1642_126_2028_n28), 
	.B2(U_dsdc_DP_OP_1642_126_2028_I5_0_), 
	.B1(U_dsdc_DP_OP_1642_126_2028_I6), 
	.A2(U_dsdc_DP_OP_1642_126_2028_I4), 
	.A1(U_dsdc_N1762));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U16 (.ZN(U_dsdc_DP_OP_1642_126_2028_n15), 
	.A(U_dsdc_DP_OP_1642_126_2028_n8));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U12 (.ZN(U_dsdc_DP_OP_1642_126_2028_n14), 
	.A(U_dsdc_DP_OP_1642_126_2028_n6));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U8 (.ZN(U_dsdc_DP_OP_1642_126_2028_n13), 
	.A(U_dsdc_DP_OP_1642_126_2028_n4));
   AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U32 (.ZN(U_dsdc_DP_OP_1642_126_2028_n24), 
	.B2(U_dsdc_DP_OP_1642_126_2028_I5_4_), 
	.B1(U_dsdc_DP_OP_1642_126_2028_I6), 
	.A2(U_dsdc_DP_OP_1642_126_2028_I4), 
	.A1(U_dsdc_N1766));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U31 (.ZN(U_dsdc_DP_OP_1642_126_2028_n61), 
	.A(U_dsdc_DP_OP_1642_126_2028_n24));
   INV_X4 U_dsdc_DP_OP_1642_126_2028_U4 (.ZN(U_dsdc_DP_OP_1642_126_2028_n12), 
	.A(U_dsdc_DP_OP_1642_126_2028_n2));
   DFFR_X2 U_dsdc_miu_push_n_reg (.RN(FE_OFN51_HRESETn), 
	.QN(ctl_push_n), 
	.Q(n82), 
	.D(FE_PHN981_U_dsdc_n329), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_dsdc_bm_bank_age_reg_2__1_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n178), 
	.Q(U_dsdc_bm_bank_age_2__1_), 
	.D(FE_PHN764_U_dsdc_n210), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_age_reg_2__3_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n459), 
	.Q(U_dsdc_bm_bank_age_2__3_), 
	.D(FE_PHN994_U_dsdc_n212), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_bank_age_reg_2__4_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n350), 
	.Q(U_dsdc_bm_bank_age_2__4_), 
	.D(FE_PHN898_U_dsdc_n213), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_ref_ack_reg (.RN(FE_OFN39_HRESETn), 
	.Q(ctl_ref_ack), 
	.D(U_dsdc_N430), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_dsdc_data_cnt_reg_5_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_data_cnt_5_), 
	.D(FE_PHN786_U_dsdc_n291), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_data_cnt_reg_4_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_data_cnt_4_), 
	.D(FE_PHN706_U_dsdc_n290), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_data_cnt_reg_3_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n437), 
	.Q(U_dsdc_data_cnt_3_), 
	.D(FE_PHN790_U_dsdc_n289), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_data_cnt_reg_2_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_data_cnt_2_), 
	.D(FE_PHN697_U_dsdc_n288), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_term_cnt_reg_1_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_term_cnt_1_), 
	.D(FE_PHN767_U_dsdc_term_cnt_nxt_1_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_term_cnt_reg_2_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n200), 
	.Q(U_dsdc_term_cnt_2_), 
	.D(FE_PHN833_U_dsdc_term_cnt_nxt_2_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_term_cnt_reg_3_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_term_cnt_3_), 
	.D(FE_PHN834_U_dsdc_term_cnt_nxt_3_), 
	.CK(HCLK__L5_N12));
   DFFS_X2 U_dsdc_miu_pop_n_reg (.SN(FE_OFN63_HRESETn), 
	.Q(ctl_pop_n), 
	.D(FE_PHN1447_U_dsdc_N429), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_dsdc_delta_delay_reg_2_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n467), 
	.Q(U_dsdc_delta_delay_2_), 
	.D(FE_PHN989_U_dsdc_n214), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_delta_delay_reg_1_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n464), 
	.Q(U_dsdc_delta_delay_1_), 
	.D(FE_PHN1529_U_dsdc_n215), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_bank_age_reg_3__0_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n304), 
	.Q(U_dsdc_bm_bank_age_3__0_), 
	.D(FE_PHN1050_U_dsdc_n218), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_age_reg_3__1_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n302), 
	.Q(U_dsdc_bm_bank_age_3__1_), 
	.D(FE_PHN792_U_dsdc_n219), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_age_reg_3__2_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n303), 
	.Q(U_dsdc_bm_bank_age_3__2_), 
	.D(FE_PHN842_U_dsdc_n220), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_age_reg_3__3_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n284), 
	.Q(U_dsdc_bm_bank_age_3__3_), 
	.D(FE_PHN998_U_dsdc_n221), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_age_reg_3__4_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n351), 
	.Q(U_dsdc_bm_bank_age_3__4_), 
	.D(FE_PHN864_U_dsdc_n222), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_status_reg_3_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n396), 
	.Q(U_dsdc_bm_bank_status_3_), 
	.D(U_dsdc_N4496), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_age_reg_1__1_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n335), 
	.Q(U_dsdc_bm_bank_age_1__1_), 
	.D(FE_PHN781_U_dsdc_n224), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_bank_age_reg_1__2_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n337), 
	.Q(U_dsdc_bm_bank_age_1__2_), 
	.D(FE_PHN799_U_dsdc_n225), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_bank_age_reg_1__3_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n460), 
	.Q(U_dsdc_bm_bank_age_1__3_), 
	.D(FE_PHN959_U_dsdc_n226), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_bank_age_reg_1__4_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n349), 
	.Q(U_dsdc_bm_bank_age_1__4_), 
	.D(FE_PHN899_U_dsdc_n227), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_bank_status_reg_1_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n383), 
	.Q(U_dsdc_bm_bank_status_1_), 
	.D(U_dsdc_N4402), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_bank_age_reg_0__1_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n435), 
	.Q(U_dsdc_bm_bank_age_0__1_), 
	.D(FE_PHN814_U_dsdc_n228), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_age_reg_0__2_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n334), 
	.Q(U_dsdc_bm_bank_age_0__2_), 
	.D(FE_PHN745_U_dsdc_n229), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_age_reg_0__3_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n458), 
	.Q(U_dsdc_bm_bank_age_0__3_), 
	.D(FE_PHN862_U_dsdc_n230), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_age_reg_0__4_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n434), 
	.Q(U_dsdc_bm_bank_age_0__4_), 
	.D(FE_PHN3053_U_dsdc_n231), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_bank_status_reg_0_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n384), 
	.Q(U_dsdc_bm_bank_status_0_), 
	.D(U_dsdc_N4355), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_num_open_bank_reg_0_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n340), 
	.Q(U_dsdc_bm_num_open_bank_0_), 
	.D(FE_PHN4293_U_dsdc_n293), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_num_open_bank_reg_1_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_dsdc_n180), 
	.Q(U_dsdc_bm_num_open_bank_1_), 
	.D(FE_PHN940_U_dsdc_n294), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_num_open_bank_reg_2_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n338), 
	.Q(U_dsdc_bm_num_open_bank_2_), 
	.D(FE_PHN901_U_dsdc_n295), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_num_open_bank_reg_4_ (.RN(FE_OFN186_HRESETn), 
	.QN(U_dsdc_n385), 
	.Q(U_dsdc_bm_num_open_bank_4_), 
	.D(FE_PHN937_U_dsdc_n297), 
	.CK(HCLK__L5_N28));
   DFFS_X2 U_dsdc_r_bm_close_all_reg (.SN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_r_bm_close_all), 
	.D(FE_PHN683_U_dsdc_n1394), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_cas_latency_cnt_reg_2_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n331), 
	.Q(U_dsdc_cas_latency_cnt_2_), 
	.D(FE_PHN1092_U_dsdc_N4128), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_cas_latency_cnt_reg_1_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_cas_latency_cnt_1_), 
	.D(FE_PHN1028_U_dsdc_N4127), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_cas_latency_cnt_reg_0_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_cas_latency_cnt_0_), 
	.D(FE_PHN4522_U_dsdc_n300), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_cas_latency_cnt_reg_3_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_cas_latency_cnt_3_), 
	.D(U_dsdc_N4129), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__12_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__12_), 
	.D(FE_PHN2381_U_dsdc_N4348), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__12_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__12_), 
	.D(FE_PHN2395_U_dsdc_N4395), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__12_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__12_), 
	.D(FE_PHN1485_U_dsdc_N4442), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__12_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__12_), 
	.D(FE_PHN1481_U_dsdc_N4489), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__11_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__11_), 
	.D(FE_PHN2424_U_dsdc_N4347), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__11_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__11_), 
	.D(FE_PHN1202_U_dsdc_N4394), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__11_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__11_), 
	.D(FE_PHN1205_U_dsdc_N4441), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__11_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__11_), 
	.D(FE_PHN2400_U_dsdc_N4488), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__10_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__10_), 
	.D(FE_PHN1570_U_dsdc_N4346), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__10_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__10_), 
	.D(FE_PHN2384_U_dsdc_N4393), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__10_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__10_), 
	.D(FE_PHN2418_U_dsdc_N4440), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__10_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__10_), 
	.D(FE_PHN1573_U_dsdc_N4487), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__9_ (.RN(FE_OFN50_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__9_), 
	.D(FE_PHN2423_U_dsdc_N4345), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__9_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__9_), 
	.D(FE_PHN2392_U_dsdc_N4392), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__9_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__9_), 
	.D(FE_PHN1300_U_dsdc_N4439), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__9_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__9_), 
	.D(FE_PHN2387_U_dsdc_N4486), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__8_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__8_), 
	.D(FE_PHN2382_U_dsdc_N4344), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__8_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__8_), 
	.D(FE_PHN2398_U_dsdc_N4391), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__8_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__8_), 
	.D(FE_PHN2405_U_dsdc_N4438), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__8_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__8_), 
	.D(FE_PHN1572_U_dsdc_N4485), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__7_ (.RN(FE_OFN50_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__7_), 
	.D(FE_PHN2419_U_dsdc_N4343), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__7_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__7_), 
	.D(FE_PHN2394_U_dsdc_N4390), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__7_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__7_), 
	.D(FE_PHN2390_U_dsdc_N4437), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__7_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__7_), 
	.D(FE_PHN1279_U_dsdc_N4484), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_r_col_addr_reg_1_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_r_col_addr_1_), 
	.D(FE_PHN3442_U_dsdc_n240), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_ras_cnt_max_reg_2_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n428), 
	.Q(U_dsdc_bm_ras_cnt_max_2_), 
	.D(FE_PHN995_U_dsdc_N4283), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_ras_cnt_max_reg_1_ (.RN(FE_OFN141_HRESETn), 
	.Q(U_dsdc_bm_ras_cnt_max_1_), 
	.D(U_dsdc_N4282), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_max_reg_0_ (.RN(FE_OFN141_HRESETn), 
	.Q(U_dsdc_bm_ras_cnt_max_0_), 
	.D(FE_PHN1413_U_dsdc_N4281), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_max_reg_3_ (.RN(FE_OFN141_HRESETn), 
	.Q(U_dsdc_bm_ras_cnt_max_3_), 
	.D(U_dsdc_N4284), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_rcd_cnt_reg_0_ (.RN(FE_OFN148_HRESETn), 
	.QN(U_dsdc_n174), 
	.Q(U_dsdc_rcd_cnt_0_), 
	.D(FE_PHN1262_U_dsdc_N4139), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_rcd_cnt_reg_2_ (.RN(FE_OFN59_HRESETn), 
	.Q(U_dsdc_rcd_cnt_2_), 
	.D(FE_PHN2978_U_dsdc_N4141), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__15_ (.RN(FE_OFN191_HRESETn), 
	.QN(U_dsdc_n425), 
	.Q(U_dsdc_bm_row_addr_0__15_), 
	.D(FE_PHN2408_U_dsdc_N4351), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__14_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__14_), 
	.D(FE_PHN1299_U_dsdc_N4350), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__13_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__13_), 
	.D(FE_PHN1209_U_dsdc_N4349), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__6_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__6_), 
	.D(FE_PHN2401_U_dsdc_N4342), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__5_ (.RN(FE_OFN50_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__5_), 
	.D(FE_PHN2425_U_dsdc_N4341), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__4_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__4_), 
	.D(FE_PHN1582_U_dsdc_N4340), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__3_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__3_), 
	.D(FE_PHN1329_U_dsdc_N4339), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__2_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__2_), 
	.D(FE_PHN2388_U_dsdc_N4338), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__1_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__1_), 
	.D(FE_PHN1322_U_dsdc_N4337), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_0__0_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_0__0_), 
	.D(FE_PHN2410_U_dsdc_N4336), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_0__2_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_rc_cnt_0__2_), 
	.D(FE_PHN3189_U_dsdc_N4334), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_0__1_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n402), 
	.Q(U_dsdc_bm_rc_cnt_0__1_), 
	.D(FE_PHN1294_U_dsdc_N4333), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_0__0_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n192), 
	.Q(U_dsdc_bm_rc_cnt_0__0_), 
	.D(FE_PHN1268_U_dsdc_N4332), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_0__3_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n441), 
	.Q(U_dsdc_bm_rc_cnt_0__3_), 
	.D(U_dsdc_N4335), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_0__2_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_ras_cnt_0__2_), 
	.D(FE_PHN3108_U_dsdc_N4321), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_0__1_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n424), 
	.Q(U_dsdc_bm_ras_cnt_0__1_), 
	.D(FE_PHN997_U_dsdc_N4320), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_0__0_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n189), 
	.Q(U_dsdc_bm_ras_cnt_0__0_), 
	.D(FE_PHN1288_U_dsdc_N4319), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_0__3_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n363), 
	.Q(U_dsdc_bm_ras_cnt_0__3_), 
	.D(FE_PHN1590_U_dsdc_N4322), 
	.CK(HCLK__L5_N28));
   DFFS_X2 U_dsdc_r_bm_open_bank_reg_0_ (.SN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_r_bm_open_bank[0]), 
	.Q(U_dsdc_n168), 
	.D(n83), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__15_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__15_), 
	.D(FE_PHN1206_U_dsdc_N4398), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__14_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__14_), 
	.D(FE_PHN2413_U_dsdc_N4397), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__13_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__13_), 
	.D(FE_PHN2386_U_dsdc_N4396), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__6_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__6_), 
	.D(FE_PHN2414_U_dsdc_N4389), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__5_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__5_), 
	.D(FE_PHN2404_U_dsdc_N4388), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__4_ (.RN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_n339), 
	.Q(U_dsdc_bm_row_addr_1__4_), 
	.D(FE_PHN2373_U_dsdc_N4387), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__3_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__3_), 
	.D(FE_PHN2396_U_dsdc_N4386), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__2_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__2_), 
	.D(FE_PHN2391_U_dsdc_N4385), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__1_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__1_), 
	.D(FE_PHN2399_U_dsdc_N4384), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_1__0_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_1__0_), 
	.D(FE_PHN1303_U_dsdc_N4383), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_1__2_ (.RN(FE_OFN173_HRESETn), 
	.Q(U_dsdc_bm_rc_cnt_1__2_), 
	.D(FE_PHN3034_U_dsdc_N4381), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_1__1_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n419), 
	.Q(U_dsdc_bm_rc_cnt_1__1_), 
	.D(FE_PHN1306_U_dsdc_N4380), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_1__0_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n193), 
	.Q(U_dsdc_bm_rc_cnt_1__0_), 
	.D(FE_PHN1271_U_dsdc_N4379), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_1__3_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n438), 
	.Q(U_dsdc_bm_rc_cnt_1__3_), 
	.D(U_dsdc_N4382), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_1__2_ (.RN(FE_OFN173_HRESETn), 
	.Q(U_dsdc_bm_ras_cnt_1__2_), 
	.D(FE_PHN3182_U_dsdc_N4368), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_1__1_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n420), 
	.Q(U_dsdc_bm_ras_cnt_1__1_), 
	.D(FE_PHN1026_U_dsdc_N4367), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_1__0_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n186), 
	.Q(U_dsdc_bm_ras_cnt_1__0_), 
	.D(FE_PHN2377_U_dsdc_N4366), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_1__3_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n364), 
	.Q(U_dsdc_bm_ras_cnt_1__3_), 
	.D(FE_PHN1496_U_dsdc_N4369), 
	.CK(HCLK__L5_N29));
   DFFS_X2 U_dsdc_r_bm_open_bank_reg_1_ (.SN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_r_bm_open_bank[1]), 
	.Q(U_dsdc_n356), 
	.D(U_dsdc_n307), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__15_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__15_), 
	.D(FE_PHN1204_U_dsdc_N4445), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__14_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__14_), 
	.D(FE_PHN2406_U_dsdc_N4444), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__13_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__13_), 
	.D(FE_PHN2383_U_dsdc_N4443), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__6_ (.RN(FE_OFN50_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__6_), 
	.D(FE_PHN1580_U_dsdc_N4436), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__5_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__5_), 
	.D(FE_PHN1575_U_dsdc_N4435), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__4_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__4_), 
	.D(FE_PHN1578_U_dsdc_N4434), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__3_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__3_), 
	.D(FE_PHN2407_U_dsdc_N4433), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__2_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__2_), 
	.D(FE_PHN2389_U_dsdc_N4432), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__1_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__1_), 
	.D(FE_PHN1291_U_dsdc_N4431), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_2__0_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_2__0_), 
	.D(FE_PHN2411_U_dsdc_N4430), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_2__2_ (.RN(FE_OFN173_HRESETn), 
	.Q(U_dsdc_bm_rc_cnt_2__2_), 
	.D(FE_PHN3033_U_dsdc_N4428), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_2__1_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n401), 
	.Q(U_dsdc_bm_rc_cnt_2__1_), 
	.D(FE_PHN1311_U_dsdc_N4427), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_2__0_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n191), 
	.Q(U_dsdc_bm_rc_cnt_2__0_), 
	.D(FE_PHN1275_U_dsdc_N4426), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_2__3_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n439), 
	.Q(U_dsdc_bm_rc_cnt_2__3_), 
	.D(FE_PHN1489_U_dsdc_N4429), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_2__2_ (.RN(FE_OFN173_HRESETn), 
	.Q(U_dsdc_bm_ras_cnt_2__2_), 
	.D(FE_PHN3109_U_dsdc_N4415), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_2__1_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n422), 
	.Q(U_dsdc_bm_ras_cnt_2__1_), 
	.D(FE_PHN1315_U_dsdc_N4414), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_2__0_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n188), 
	.Q(U_dsdc_bm_ras_cnt_2__0_), 
	.D(FE_PHN1410_U_dsdc_N4413), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_2__3_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n365), 
	.Q(U_dsdc_bm_ras_cnt_2__3_), 
	.D(FE_PHN1495_U_dsdc_N4416), 
	.CK(HCLK__L5_N31));
   DFFS_X2 U_dsdc_r_bm_open_bank_reg_2_ (.SN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_n164), 
	.D(U_dsdc_n310), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__15_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__15_), 
	.D(FE_PHN2416_U_dsdc_N4492), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__14_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__14_), 
	.D(FE_PHN2409_U_dsdc_N4491), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__13_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__13_), 
	.D(FE_PHN2380_U_dsdc_N4490), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__6_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__6_), 
	.D(FE_PHN2402_U_dsdc_N4483), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__5_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__5_), 
	.D(FE_PHN1581_U_dsdc_N4482), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__4_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__4_), 
	.D(FE_PHN1576_U_dsdc_N4481), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__3_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__3_), 
	.D(FE_PHN2397_U_dsdc_N4480), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__2_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__2_), 
	.D(FE_PHN1292_U_dsdc_N4479), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__1_ (.RN(FE_OFN191_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__1_), 
	.D(FE_PHN2393_U_dsdc_N4478), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_bm_row_addr_reg_3__0_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_bm_row_addr_3__0_), 
	.D(FE_PHN2417_U_dsdc_N4477), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_3__2_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_bm_rc_cnt_3__2_), 
	.D(FE_PHN3013_U_dsdc_N4475), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_3__1_ (.RN(FE_OFN36_HRESETn), 
	.QN(U_dsdc_n400), 
	.Q(U_dsdc_bm_rc_cnt_3__1_), 
	.D(FE_PHN1310_U_dsdc_N4474), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_3__0_ (.RN(FE_OFN36_HRESETn), 
	.QN(U_dsdc_n190), 
	.Q(U_dsdc_bm_rc_cnt_3__0_), 
	.D(FE_PHN1287_U_dsdc_N4473), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_rc_cnt_reg_3__3_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n442), 
	.Q(U_dsdc_bm_rc_cnt_3__3_), 
	.D(FE_PHN1486_U_dsdc_N4476), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_3__2_ (.RN(FE_OFN141_HRESETn), 
	.Q(U_dsdc_bm_ras_cnt_3__2_), 
	.D(FE_PHN3245_U_dsdc_N4462), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_3__1_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n421), 
	.Q(U_dsdc_bm_ras_cnt_3__1_), 
	.D(FE_PHN921_U_dsdc_N4461), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_3__0_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n187), 
	.Q(U_dsdc_bm_ras_cnt_3__0_), 
	.D(FE_PHN1090_U_dsdc_N4460), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_bm_ras_cnt_reg_3__3_ (.RN(FE_OFN141_HRESETn), 
	.QN(U_dsdc_n382), 
	.Q(U_dsdc_bm_ras_cnt_3__3_), 
	.D(U_dsdc_N4463), 
	.CK(HCLK__L5_N31));
   DFFS_X2 U_dsdc_r_bm_open_bank_reg_3_ (.SN(FE_OFN45_HRESETn), 
	.QN(U_dsdc_r_bm_open_bank[3]), 
	.Q(U_dsdc_n185), 
	.D(U_dsdc_n313), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_rcar_cnt2_reg_2_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_rcar_cnt2_2_), 
	.D(FE_PHN751_U_dsdc_rcar_cnt2_nxt_2_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_rcar_cnt2_reg_1_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_rcar_cnt2_1_), 
	.D(FE_PHN900_U_dsdc_rcar_cnt2_nxt_1_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_rcar_cnt2_reg_0_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_rcar_cnt2_0_), 
	.D(FE_PHN1213_U_dsdc_rcar_cnt2_nxt_0_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_wtr_cnt_reg_2_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_wtr_cnt_2_), 
	.D(FE_PHN742_U_dsdc_wtr_cnt_nxt_2_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_wtr_cnt_reg_0_ (.RN(FE_OFN142_HRESETn), 
	.QN(U_dsdc_n398), 
	.Q(U_dsdc_wtr_cnt_0_), 
	.D(FE_PHN933_U_dsdc_wtr_cnt_nxt_0_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_r_row_addr_reg_10_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_r_row_addr_10_), 
	.D(FE_PHN3431_U_dsdc_n256), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_r_row_addr_reg_12_ (.RN(FE_OFN50_HRESETn), 
	.Q(U_dsdc_r_row_addr_12_), 
	.D(FE_PHN1326_U_dsdc_n258), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_dsdc_r_row_addr_reg_4_ (.RN(FE_OFN50_HRESETn), 
	.Q(U_dsdc_r_row_addr_4_), 
	.D(FE_PHN3440_U_dsdc_n265), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_dsdc_r_row_addr_reg_5_ (.RN(FE_OFN50_HRESETn), 
	.Q(U_dsdc_r_row_addr_5_), 
	.D(FE_PHN3415_U_dsdc_n266), 
	.CK(HCLK__L5_N33));
   DFFR_X1 U_dsdc_r_row_addr_reg_6_ (.RN(FE_OFN50_HRESETn), 
	.Q(U_dsdc_r_row_addr_6_), 
	.D(FE_PHN3407_U_dsdc_n267), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_r_row_addr_reg_8_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_r_row_addr_8_), 
	.D(FE_PHN3446_U_dsdc_n269), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_cas_cnt_reg_5_ (.RN(FE_OFN141_HRESETn), 
	.Q(U_dsdc_cas_cnt_5_), 
	.D(FE_PHN1338_U_dsdc_cas_cnt_nxt_5_), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_cas_cnt_reg_4_ (.RN(FE_OFN141_HRESETn), 
	.Q(U_dsdc_cas_cnt_4_), 
	.D(U_dsdc_cas_cnt_nxt[4]), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_cas_cnt_reg_3_ (.RN(FE_OFN141_HRESETn), 
	.Q(U_dsdc_cas_cnt_3_), 
	.D(FE_PHN3194_U_dsdc_cas_cnt_nxt_3_), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_cas_cnt_reg_2_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_cas_cnt_2_), 
	.D(FE_PHN3087_U_dsdc_cas_cnt_nxt_2_), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_cas_cnt_reg_1_ (.RN(FE_OFN141_HRESETn), 
	.Q(U_dsdc_cas_cnt_1_), 
	.D(FE_PHN1218_U_dsdc_cas_cnt_nxt_1_), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_r_burst_size_reg_1_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_r_burst_size_1_), 
	.D(U_dsdc_n272), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_r_burst_size_reg_2_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_r_burst_size_2_), 
	.D(FE_PHN2044_U_dsdc_n273), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_r_close_bank_addr_reg_0_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n292), 
	.Q(U_dsdc_r_close_bank_addr_0_), 
	.D(U_dsdc_close_bank_addr_0_), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_r_bm_close_bank_reg_1_ (.RN(FE_OFN173_HRESETn), 
	.Q(U_dsdc_r_bm_close_bank_1_), 
	.D(U_dsdc_bm_close_bank_1_), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_r_bm_close_bank_reg_0_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_r_bm_close_bank_0_), 
	.D(U_dsdc_bm_close_bank_0_), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_r_bm_close_bank_reg_3_ (.RN(FE_OFN45_HRESETn), 
	.Q(U_dsdc_r_bm_close_bank_3_), 
	.D(U_dsdc_bm_close_bank_3_), 
	.CK(HCLK__L5_N30));
   DFFR_X1 U_dsdc_r_close_bank_addr_reg_1_ (.RN(FE_OFN173_HRESETn), 
	.Q(U_dsdc_r_close_bank_addr_1_), 
	.D(U_dsdc_close_bank_addr_1_), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_auto_ref_en_reg (.RN(FE_OFN39_HRESETn), 
	.QN(n94), 
	.Q(ctl_auto_ref_en), 
	.D(FE_PHN757_U_dsdc_auto_ref_en_nxt), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_dsdc_init_cnt_reg_15_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_dsdc_init_cnt_15_), 
	.D(FE_PHN1295_U_dsdc_n418), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_dsdc_init_cnt_reg_14_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_dsdc_init_cnt_14_), 
	.D(FE_PHN1328_U_dsdc_n417), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_dsdc_init_cnt_reg_13_ (.RN(FE_OFN172_HRESETn), 
	.Q(U_dsdc_init_cnt_13_), 
	.D(FE_PHN3081_U_dsdc_n416), 
	.CK(hclk));
   DFFR_X1 U_dsdc_init_cnt_reg_12_ (.RN(FE_OFN172_HRESETn), 
	.Q(U_dsdc_init_cnt_12_), 
	.D(FE_PHN3112_U_dsdc_n415), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_init_cnt_reg_11_ (.RN(FE_OFN172_HRESETn), 
	.Q(U_dsdc_init_cnt_11_), 
	.D(FE_PHN3127_U_dsdc_n414), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_init_cnt_reg_10_ (.RN(FE_OFN172_HRESETn), 
	.Q(U_dsdc_init_cnt_10_), 
	.D(FE_PHN1216_U_dsdc_n413), 
	.CK(hclk));
   DFFR_X1 U_dsdc_init_cnt_reg_9_ (.RN(FE_OFN172_HRESETn), 
	.Q(U_dsdc_init_cnt_9_), 
	.D(FE_PHN922_U_dsdc_n412), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_init_cnt_reg_8_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_dsdc_init_cnt_8_), 
	.D(FE_PHN3119_U_dsdc_n411), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_dsdc_init_cnt_reg_7_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_dsdc_init_cnt_7_), 
	.D(FE_PHN925_U_dsdc_n410), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_dsdc_init_cnt_reg_6_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_dsdc_init_cnt_6_), 
	.D(FE_PHN1215_U_dsdc_n409), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_init_cnt_reg_5_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_dsdc_init_cnt_5_), 
	.D(FE_PHN942_U_dsdc_n408), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_init_cnt_reg_4_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_dsdc_init_cnt_4_), 
	.D(FE_PHN3123_U_dsdc_n407), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_init_cnt_reg_3_ (.RN(FE_OFN172_HRESETn), 
	.Q(U_dsdc_init_cnt_3_), 
	.D(FE_PHN938_U_dsdc_n406), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_init_cnt_reg_2_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_dsdc_n468), 
	.Q(U_dsdc_init_cnt_2_), 
	.D(FE_PHN1047_U_dsdc_n405), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_init_cnt_reg_1_ (.RN(FE_OFN31_HRESETn), 
	.Q(U_dsdc_init_cnt_1_), 
	.D(FE_PHN1099_U_dsdc_n404), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_init_cnt_reg_0_ (.RN(FE_OFN172_HRESETn), 
	.Q(U_dsdc_init_cnt_0_), 
	.D(FE_PHN1658_U_dsdc_n403), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_dsdc_row_cnt_reg_0_ (.RN(FE_OFN186_HRESETn), 
	.QN(U_dsdc_n462), 
	.Q(U_dsdc_row_cnt_0_), 
	.D(FE_PHN1623_U_dsdc_n366), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_10_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n208), 
	.Q(U_dsdc_row_cnt_10_), 
	.D(FE_PHN1121_U_dsdc_n367), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_11_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_row_cnt_11_), 
	.D(FE_PHN986_U_dsdc_n368), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_13_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n197), 
	.Q(U_dsdc_row_cnt_13_), 
	.D(FE_PHN987_U_dsdc_n370), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_14_ (.RN(FE_OFN186_HRESETn), 
	.QN(U_dsdc_n202), 
	.Q(U_dsdc_row_cnt_14_), 
	.D(FE_PHN1122_U_dsdc_n371), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_15_ (.RN(FE_OFN186_HRESETn), 
	.QN(U_dsdc_n426), 
	.Q(U_dsdc_row_cnt_15_), 
	.D(FE_PHN1123_U_dsdc_n372), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_1_ (.RN(FE_OFN186_HRESETn), 
	.QN(U_dsdc_n465), 
	.Q(U_dsdc_row_cnt_1_), 
	.D(FE_PHN1247_U_dsdc_n373), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_2_ (.RN(FE_OFN36_HRESETn), 
	.QN(U_dsdc_n204), 
	.Q(U_dsdc_row_cnt_2_), 
	.D(FE_PHN905_U_dsdc_n374), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_3_ (.RN(FE_OFN186_HRESETn), 
	.Q(U_dsdc_row_cnt_3_), 
	.D(FE_PHN953_U_dsdc_n375), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_4_ (.RN(FE_OFN36_HRESETn), 
	.QN(U_dsdc_n207), 
	.Q(U_dsdc_row_cnt_4_), 
	.D(FE_PHN1045_U_dsdc_n376), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_row_cnt_reg_5_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_row_cnt_5_), 
	.D(FE_PHN985_U_dsdc_n377), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_row_cnt_reg_6_ (.RN(FE_OFN36_HRESETn), 
	.QN(U_dsdc_n206), 
	.Q(U_dsdc_row_cnt_6_), 
	.D(FE_PHN983_U_dsdc_n378), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_row_cnt_reg_7_ (.RN(FE_OFN36_HRESETn), 
	.Q(U_dsdc_row_cnt_7_), 
	.D(FE_PHN906_U_dsdc_n379), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_row_cnt_reg_8_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n205), 
	.Q(U_dsdc_row_cnt_8_), 
	.D(FE_PHN1046_U_dsdc_n380), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_row_cnt_reg_9_ (.RN(FE_OFN44_HRESETn), 
	.Q(U_dsdc_row_cnt_9_), 
	.D(FE_PHN984_U_dsdc_n381), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_rcar_cnt1_reg_3_ (.RN(FE_OFN63_HRESETn), 
	.Q(U_dsdc_rcar_cnt1_3_), 
	.D(FE_PHN1053_U_dsdc_rcar_cnt1_nxt_3_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_rcar_cnt1_reg_2_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_rcar_cnt1_2_), 
	.D(FE_PHN1051_U_dsdc_rcar_cnt1_nxt_2_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_rcar_cnt1_reg_1_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_rcar_cnt1_1_), 
	.D(FE_PHN1208_U_dsdc_rcar_cnt1_nxt_1_), 
	.CK(hclk));
   DFFR_X1 U_dsdc_rcar_cnt1_reg_0_ (.RN(FE_OFN63_HRESETn), 
	.Q(U_dsdc_rcar_cnt1_0_), 
	.D(FE_PHN2037_U_dsdc_rcar_cnt1_nxt_0_), 
	.CK(hclk));
   DFFR_X1 U_dsdc_xsr_cnt_reg_0_ (.RN(FE_OFN63_HRESETn), 
	.Q(U_dsdc_xsr_cnt_0_), 
	.D(FE_PHN1659_U_dsdc_n386), 
	.CK(hclk));
   DFFR_X1 U_dsdc_xsr_cnt_reg_1_ (.RN(FE_OFN63_HRESETn), 
	.Q(U_dsdc_xsr_cnt_1_), 
	.D(FE_PHN1023_U_dsdc_n387), 
	.CK(hclk));
   DFFR_X1 U_dsdc_xsr_cnt_reg_2_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_xsr_cnt_2_), 
	.D(FE_PHN1210_U_dsdc_n388), 
	.CK(hclk));
   DFFR_X1 U_dsdc_xsr_cnt_reg_3_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_xsr_cnt_3_), 
	.D(FE_PHN896_U_dsdc_n389), 
	.CK(hclk));
   DFFR_X1 U_dsdc_xsr_cnt_reg_4_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_xsr_cnt_4_), 
	.D(FE_PHN1321_U_dsdc_n390), 
	.CK(hclk));
   DFFR_X1 U_dsdc_xsr_cnt_reg_5_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_xsr_cnt_5_), 
	.D(FE_PHN1001_U_dsdc_n391), 
	.CK(hclk));
   DFFR_X1 U_dsdc_xsr_cnt_reg_7_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_xsr_cnt_7_), 
	.D(FE_PHN1323_U_dsdc_n393), 
	.CK(hclk));
   DFFR_X1 U_dsdc_xsr_cnt_reg_8_ (.RN(FE_OFN142_HRESETn), 
	.Q(U_dsdc_xsr_cnt_8_), 
	.D(FE_PHN1094_U_dsdc_n394), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_operation_cs_reg_2_ (.RN(FE_OFN142_HRESETn), 
	.QN(U_dsdc_n341), 
	.Q(U_dsdc_operation_cs_2_), 
	.D(FE_PHN3473_U_dsdc_n2095), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_operation_cs_reg_4_ (.RN(FE_OFN142_HRESETn), 
	.QN(U_dsdc_n432), 
	.D(FE_PHN854_U_dsdc_n2093), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_num_init_ref_cnt_reg_3_ (.RN(FE_OFN63_HRESETn), 
	.Q(U_dsdc_num_init_ref_cnt_3_), 
	.D(FE_PHN964_U_dsdc_n431), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_dsdc_operation_cs_reg_0_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_dsdc_n344), 
	.Q(U_dsdc_operation_cs_0_), 
	.D(FE_PHN882_U_dsdc_n2097), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_operation_cs_reg_1_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_dsdc_n343), 
	.Q(U_dsdc_operation_cs_1_), 
	.D(FE_PHN758_U_dsdc_n2096), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_t_xp_cnt_reg_1_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dsdc_n474), 
	.Q(U_dsdc_t_xp_cnt_1_), 
	.D(FE_PHN1683_U_dsdc_N4229), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_t_xp_cnt_reg_0_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dsdc_n239), 
	.Q(U_dsdc_t_xp_cnt_0_), 
	.D(FE_PHN1430_U_dsdc_N4228), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_access_cs_reg_4_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dsdc_n167), 
	.Q(U_dsdc_access_cs_4_), 
	.D(FE_PHN1012_U_dsdc_n_2088_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_wr_cnt_reg_2_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_dsdc_wr_cnt_2_), 
	.D(FE_PHN891_U_dsdc_wr_cnt_nxt_2_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_wr_cnt_reg_1_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_dsdc_n195), 
	.D(FE_PHN1381_U_dsdc_wr_cnt_nxt_1_), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_wr_cnt_reg_0_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_dsdc_n397), 
	.Q(U_dsdc_wr_cnt_0_), 
	.D(FE_PHN1173_U_dsdc_wr_cnt_nxt_0_), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_access_cs_reg_3_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dsdc_n173), 
	.Q(U_dsdc_access_cs_3_), 
	.D(FE_PHN990_U_dsdc_n_2089_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_rp_cnt2_reg_2_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_dsdc_rp_cnt2_2_), 
	.D(FE_PHN924_U_dsdc_rp_cnt2_nxt_2_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_rp_cnt2_reg_1_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_dsdc_n309), 
	.D(FE_PHN838_U_dsdc_rp_cnt2_nxt_1_), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_dsdc_r_rw_reg (.SN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n166), 
	.Q(U_dsdc_r_rw), 
	.D(FE_PHN4397_U_dsdc_n279), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_r_chip_slct_reg_0_ (.RN(FE_OFN44_HRESETn), 
	.QN(U_dsdc_n361), 
	.Q(U_dsdc_r_chip_slct_0_), 
	.D(FE_PHN1483_U_dsdc_n280), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_dsdc_access_cs_reg_0_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dsdc_n170), 
	.Q(U_dsdc_access_cs_0_), 
	.D(U_dsdc_n[2092]), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_term_cnt_reg_4_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n457), 
	.Q(U_dsdc_term_cnt_4_), 
	.D(FE_PHN835_U_dsdc_term_cnt_nxt_4_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_data_cnt_reg_0_ (.RN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_n347), 
	.Q(U_dsdc_data_cnt_0_), 
	.D(FE_PHN696_U_dsdc_n286), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_access_cs_reg_1_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dsdc_n298), 
	.Q(U_dsdc_access_cs_1_), 
	.D(U_dsdc_n[2091]), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dsdc_bm_bank_status_reg_2_ (.RN(FE_OFN173_HRESETn), 
	.QN(U_dsdc_n395), 
	.Q(U_dsdc_bm_bank_status_2_), 
	.D(U_dsdc_N4449), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_r_bm_close_bank_reg_2_ (.RN(FE_OFN173_HRESETn), 
	.Q(U_dsdc_r_bm_close_bank_2_), 
	.D(U_dsdc_bm_close_bank_2_), 
	.CK(HCLK__L5_N29));
   DFFR_X1 U_dsdc_r_cas_latency_reg_1_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_r_cas_latency_1_), 
	.D(FE_PHN907_U_dsdc_cas_latency_1_), 
	.CK(HCLK__L5_N31));
   DFFR_X1 U_dsdc_r_cas_latency_reg_2_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dsdc_r_cas_latency_2_), 
	.D(U_dsdc_cas_latency_2_), 
	.CK(HCLK__L5_N31));
   DFFS_X2 U_dsdc_r_cas_latency_reg_3_ (.SN(FE_OFN64_HRESETn), 
	.QN(U_dsdc_r_cas_latency_3_), 
	.D(FE_PHN788_U_dsdc_n554), 
	.CK(HCLK__L5_N31));
   OAI22_X1 U_cr_U595 (.ZN(U_cr_n507), 
	.B2(U_cr_n17), 
	.B1(U_cr_n519), 
	.A2(U_cr_n531), 
	.A1(FE_PHN2432_n27));
   NAND2_X1 U_cr_U594 (.ZN(U_cr_n504), 
	.A2(hiu_rw), 
	.A1(U_cr_n17));
   AOI22_X1 U_cr_U593 (.ZN(U_cr_n387), 
	.B2(cr_row_addr_width[1]), 
	.B1(U_cr_n407), 
	.A2(s_read_pipe[0]), 
	.A1(U_cr_n422));
   INV_X4 U_cr_U591 (.ZN(U_cr_n204), 
	.A(U_cr_n487));
   INV_X4 U_cr_U590 (.ZN(U_cr_n203), 
	.A(U_cr_n492));
   NAND3_X2 U_cr_U589 (.ZN(U_cr_n182), 
	.A3(U_cr_n179), 
	.A2(U_cr_n185), 
	.A1(U_cr_n180));
   NOR2_X2 U_cr_U588 (.ZN(U_cr_n424), 
	.A2(U_cr_n308), 
	.A1(hiu_haddr[2]));
   NAND3_X2 U_cr_U587 (.ZN(U_cr_n416), 
	.A3(U_cr_n283), 
	.A2(U_cr_n320), 
	.A1(U_cr_n227));
   OR2_X4 U_cr_U586 (.ZN(U_cr_n25), 
	.A2(U_cr_n263), 
	.A1(hiu_haddr[2]));
   NAND3_X2 U_cr_U585 (.ZN(U_cr_n391), 
	.A3(U_cr_n227), 
	.A2(hiu_haddr[2]), 
	.A1(U_cr_n283));
   INV_X4 U_cr_U584 (.ZN(U_cr_n430), 
	.A(U_cr_n391));
   AOI221_X2 U_cr_U583 (.ZN(U_cr_n239), 
	.C2(U_addrdec_n40), 
	.C1(ad_cr_data_mask[3]), 
	.B2(big_endian), 
	.B1(ad_cr_data_mask[0]), 
	.A(U_cr_n237));
   NOR2_X2 U_cr_U582 (.ZN(U_cr_n258), 
	.A2(U_cr_n241), 
	.A1(big_endian));
   NOR2_X2 U_cr_U581 (.ZN(U_cr_n259), 
	.A2(U_cr_n241), 
	.A1(U_cr_n242));
   NOR2_X2 U_cr_U580 (.ZN(U_cr_n215), 
	.A2(U_cr_n416), 
	.A1(U_cr_n526));
   INV_X4 U_cr_U579 (.ZN(U_cr_n229), 
	.A(U_cr_n230));
   INV_X4 U_cr_U578 (.ZN(U_cr_n312), 
	.A(U_cr_n313));
   INV_X4 U_cr_U577 (.ZN(U_cr_n538), 
	.A(U_cr_n536));
   INV_X4 U_cr_U576 (.ZN(U_cr_n304), 
	.A(U_cr_n305));
   INV_X4 U_cr_U575 (.ZN(U_cr_n288), 
	.A(U_cr_n289));
   NAND3_X1 U_cr_U574 (.ZN(U_cr_n174), 
	.A3(U_cr_n23), 
	.A2(U_cr_n17), 
	.A1(U_cr_n194));
   NOR2_X2 U_cr_U573 (.ZN(U_cr_n499), 
	.A2(U_addrdec_n40), 
	.A1(U_cr_n182));
   INV_X4 U_cr_U572 (.ZN(U_cr_n267), 
	.A(U_cr_n268));
   AND2_X4 U_cr_U571 (.ZN(U_cr_n511), 
	.A2(U_cr_n223), 
	.A1(FE_PHN4616_n27));
   NOR2_X2 U_cr_U570 (.ZN(U_cr_n221), 
	.A2(U_cr_n416), 
	.A1(U_cr_n544));
   NOR2_X2 U_cr_U569 (.ZN(U_cr_n307), 
	.A2(U_cr_n358), 
	.A1(U_cr_n544));
   NOR2_X2 U_cr_U568 (.ZN(U_cr_n542), 
	.A2(U_cr_n334), 
	.A1(U_cr_n544));
   INV_X4 U_cr_U567 (.ZN(U_cr_n292), 
	.A(U_cr_n294));
   INV_X4 U_cr_U566 (.ZN(U_cr_n269), 
	.A(U_cr_n270));
   NAND3_X1 U_cr_U565 (.ZN(U_cr_n195), 
	.A3(FE_PHN2432_n27), 
	.A2(U_cr_n194), 
	.A1(hiu_reg_req));
   XNOR2_X2 U_cr_U564 (.ZN(U_cr_N574), 
	.B(U_cr_n210), 
	.A(U_cr_sctlr_16_));
   XNOR2_X2 U_cr_U563 (.ZN(U_cr_N577), 
	.B(U_cr_n282), 
	.A(U_cr_stmg0r_26));
   INV_X4 U_cr_U562 (.ZN(U_cr_n205), 
	.A(U_cr_n236));
   INV_X4 U_cr_U561 (.ZN(U_cr_n396), 
	.A(U_cr_n422));
   AOI222_X2 U_cr_U560 (.ZN(U_cr_n531), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[11]), 
	.B2(hiu_wr_data[27]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[3]), 
	.A1(U_addrdec_n40));
   INV_X4 U_cr_U559 (.ZN(U_cr_n334), 
	.A(U_cr_n424));
   NAND3_X2 U_cr_U558 (.ZN(U_cr_n315), 
	.A3(U_cr_n283), 
	.A2(hiu_addr[4]), 
	.A1(U_cr_n284));
   INV_X4 U_cr_U557 (.ZN(U_cr_n358), 
	.A(U_cr_n423));
   NAND2_X2 U_cr_U556 (.ZN(U_cr_n487), 
	.A2(big_endian), 
	.A1(U_cr_n182));
   NAND2_X2 U_cr_U555 (.ZN(U_cr_n492), 
	.A2(U_addrdec_n40), 
	.A1(U_cr_n182));
   AOI221_X2 U_cr_U554 (.ZN(U_cr_n223), 
	.C2(ad_cr_data_mask[1]), 
	.C1(big_endian), 
	.B2(ad_cr_data_mask[2]), 
	.B1(U_addrdec_n40), 
	.A(U_cr_n205));
   INV_X4 U_cr_U553 (.ZN(U_cr_n231), 
	.A(U_cr_n232));
   AOI21_X2 U_cr_U552 (.ZN(U_cr_n187), 
	.B2(FE_PHN1401_U_cr_cr_cs_1_), 
	.B1(hiu_rw), 
	.A(FE_PHN837_U_cr_cr_cs_0_));
   INV_X4 U_cr_U551 (.ZN(U_cr_n199), 
	.A(U_cr_n190));
   OAI211_X2 U_cr_U550 (.ZN(cr_pop_n), 
	.C2(U_cr_n24), 
	.C1(U_cr_n187), 
	.B(U_cr_n199), 
	.A(U_cr_n186));
   AOI222_X2 U_cr_U548 (.ZN(U_cr_n548), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[0]), 
	.B2(hiu_wr_data[16]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[8]), 
	.A1(FE_OFN357_U_addrdec_n40));
   NOR3_X2 U_cr_U547 (.ZN(U_cr_n212), 
	.A3(FE_OFN220_hiu_burst_size_0_), 
	.A2(hiu_burst_size[5]), 
	.A1(hiu_burst_size[3]));
   NAND3_X2 U_cr_U546 (.ZN(U_cr_n550), 
	.A3(U_cr_n211), 
	.A2(U_cr_n212), 
	.A1(hiu_burst_size[1]));
   NAND2_X2 U_cr_U545 (.ZN(U_cr_n318), 
	.A2(U_cr_n550), 
	.A1(hiu_haddr[1]));
   NOR4_X2 U_cr_U544 (.ZN(U_cr_n227), 
	.A4(hiu_addr[4]), 
	.A3(hiu_addr[6]), 
	.A2(hiu_addr[7]), 
	.A1(hiu_addr[5]));
   NAND2_X2 U_cr_U543 (.ZN(U_cr_n236), 
	.A2(U_cr_n200), 
	.A1(U_cr_n202));
   NAND2_X2 U_cr_U542 (.ZN(U_cr_n262), 
	.A2(U_cr_n239), 
	.A1(U_cr_n238));
   NAND2_X2 U_cr_U541 (.ZN(U_cr_n241), 
	.A2(FE_PHN4616_n27), 
	.A1(U_cr_n239));
   NAND2_X2 U_cr_U540 (.ZN(U_cr_n257), 
	.A2(U_cr_n239), 
	.A1(U_cr_n240));
   AOI22_X2 U_cr_U539 (.ZN(U_cr_n244), 
	.B2(U_cr_n257), 
	.B1(cr_t_rc[2]), 
	.A2(U_cr_n258), 
	.A1(hiu_wr_data[24]));
   AOI222_X2 U_cr_U538 (.ZN(U_cr_n546), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[1]), 
	.B2(hiu_wr_data[17]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[9]), 
	.A1(FE_OFN357_U_addrdec_n40));
   AOI22_X2 U_cr_U537 (.ZN(U_cr_n246), 
	.B2(U_cr_n257), 
	.B1(cr_t_rc[3]), 
	.A2(U_cr_n258), 
	.A1(FE_OFN227_hiu_data_25_));
   OAI211_X2 U_cr_U536 (.ZN(U_cr_N414), 
	.C2(U_cr_n262), 
	.C1(U_cr_n546), 
	.B(U_cr_n245), 
	.A(U_cr_n246));
   AOI222_X2 U_cr_U535 (.ZN(U_cr_n545), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[2]), 
	.B2(hiu_wr_data[18]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[10]), 
	.A1(FE_OFN357_U_addrdec_n40));
   AOI22_X2 U_cr_U534 (.ZN(U_cr_n248), 
	.B2(U_cr_n257), 
	.B1(U_cr_stmg0r_26), 
	.A2(U_cr_n258), 
	.A1(hiu_wr_data[26]));
   OAI211_X2 U_cr_U533 (.ZN(U_cr_N415), 
	.C2(U_cr_n262), 
	.C1(U_cr_n545), 
	.B(U_cr_n247), 
	.A(U_cr_n248));
   AOI22_X2 U_cr_U532 (.ZN(U_cr_n252), 
	.B2(U_cr_n257), 
	.B1(cr_t_xsr[5]), 
	.A2(U_cr_n258), 
	.A1(hiu_wr_data[28]));
   AOI22_X2 U_cr_U531 (.ZN(U_cr_n250), 
	.B2(U_cr_n257), 
	.B1(cr_t_xsr[4]), 
	.A2(U_cr_n258), 
	.A1(hiu_wr_data[27]));
   AOI22_X2 U_cr_U530 (.ZN(U_cr_n254), 
	.B2(U_cr_n257), 
	.B1(cr_t_xsr[6]), 
	.A2(U_cr_n258), 
	.A1(FE_OFN224_hiu_data_29_));
   AOI22_X2 U_cr_U529 (.ZN(U_cr_n261), 
	.B2(U_cr_n257), 
	.B1(cr_t_xsr[8]), 
	.A2(U_cr_n258), 
	.A1(hiu_wr_data[31]));
   AOI22_X2 U_cr_U528 (.ZN(U_cr_n256), 
	.B2(U_cr_n257), 
	.B1(cr_t_xsr[7]), 
	.A2(U_cr_n258), 
	.A1(FE_OFN223_hiu_data_30_));
   INV_X4 U_cr_U527 (.ZN(U_cr_n317), 
	.A(U_cr_n318));
   AOI221_X2 U_cr_U526 (.ZN(U_cr_n213), 
	.C2(ad_cr_data_mask[0]), 
	.C1(U_addrdec_n40), 
	.B2(ad_cr_data_mask[3]), 
	.B1(big_endian), 
	.A(U_cr_n205));
   AOI222_X2 U_cr_U525 (.ZN(U_cr_n529), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[13]), 
	.B2(hiu_wr_data[29]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[5]), 
	.A1(FE_OFN357_U_addrdec_n40));
   INV_X4 U_cr_U524 (.ZN(U_cr_n214), 
	.A(U_cr_n215));
   AOI22_X2 U_cr_U523 (.ZN(U_cr_N300), 
	.B2(U_cr_n214), 
	.B1(U_cr_n21), 
	.A2(U_cr_n529), 
	.A1(U_cr_n215));
   AOI222_X2 U_cr_U522 (.ZN(U_cr_n530), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[12]), 
	.B2(hiu_wr_data[28]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[4]), 
	.A1(U_addrdec_n40));
   AOI22_X2 U_cr_U521 (.ZN(U_cr_N299), 
	.B2(U_cr_n214), 
	.B1(U_cr_n66), 
	.A2(U_cr_n530), 
	.A1(U_cr_n215));
   AOI222_X2 U_cr_U520 (.ZN(U_cr_n528), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[14]), 
	.B2(hiu_wr_data[30]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[6]), 
	.A1(FE_OFN357_U_addrdec_n40));
   AOI22_X2 U_cr_U519 (.ZN(U_cr_N301), 
	.B2(U_cr_n214), 
	.B1(U_cr_n42), 
	.A2(FE_OFN333_U_cr_n528), 
	.A1(U_cr_n215));
   NAND2_X2 U_cr_U518 (.ZN(U_cr_n263), 
	.A2(U_cr_n227), 
	.A1(hiu_haddr[3]));
   INV_X4 U_cr_U517 (.ZN(U_cr_n272), 
	.A(U_cr_n273));
   AOI22_X2 U_cr_U516 (.ZN(U_cr_N554), 
	.B2(U_cr_n272), 
	.B1(U_cr_n139), 
	.A2(U_cr_n530), 
	.A1(U_cr_n273));
   AOI22_X2 U_cr_U515 (.ZN(U_cr_N555), 
	.B2(U_cr_n272), 
	.B1(U_cr_n132), 
	.A2(U_cr_n529), 
	.A1(U_cr_n273));
   AOI22_X2 U_cr_U514 (.ZN(U_cr_N556), 
	.B2(U_cr_n272), 
	.B1(U_cr_n40), 
	.A2(U_cr_n528), 
	.A1(U_cr_n273));
   AOI221_X2 U_cr_U513 (.ZN(U_cr_N551), 
	.C2(U_cr_n272), 
	.C1(U_cr_n39), 
	.B2(U_cr_n273), 
	.B1(U_cr_n516), 
	.A(clear_sr_dp));
   AOI22_X2 U_cr_U512 (.ZN(U_cr_N390), 
	.B2(U_cr_n229), 
	.B1(FE_PHN3106_U_cr_n43), 
	.A2(U_cr_n516), 
	.A1(U_cr_n230));
   AOI222_X2 U_cr_U511 (.ZN(U_cr_n527), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[15]), 
	.B2(hiu_wr_data[31]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[7]), 
	.A1(FE_OFN357_U_addrdec_n40));
   AOI22_X2 U_cr_U510 (.ZN(U_cr_N396), 
	.B2(U_cr_n229), 
	.B1(U_cr_n133), 
	.A2(U_cr_n527), 
	.A1(U_cr_n230));
   AOI22_X2 U_cr_U509 (.ZN(U_cr_N392), 
	.B2(U_cr_n229), 
	.B1(U_cr_n120), 
	.A2(U_cr_n531), 
	.A1(U_cr_n230));
   AOI22_X2 U_cr_U508 (.ZN(U_cr_N394), 
	.B2(U_cr_n229), 
	.B1(U_cr_n54), 
	.A2(U_cr_n529), 
	.A1(U_cr_n230));
   AOI22_X2 U_cr_U507 (.ZN(U_cr_N736), 
	.B2(U_cr_n312), 
	.B1(U_cr_n156), 
	.A2(U_cr_n531), 
	.A1(U_cr_n313));
   NOR3_X2 U_cr_U506 (.ZN(U_cr_n525), 
	.A3(U_cr_n315), 
	.A2(U_cr_n316), 
	.A1(U_cr_n320));
   INV_X4 U_cr_U505 (.ZN(U_cr_n543), 
	.A(U_cr_n525));
   AOI22_X2 U_cr_U504 (.ZN(U_cr_n83), 
	.B2(U_cr_n538), 
	.B1(U_cr_n152), 
	.A2(U_cr_n530), 
	.A1(U_cr_n536));
   AOI22_X2 U_cr_U503 (.ZN(U_cr_N740), 
	.B2(U_cr_n312), 
	.B1(U_cr_n159), 
	.A2(FE_OFN336_U_cr_n527), 
	.A1(U_cr_n313));
   AOI22_X2 U_cr_U502 (.ZN(U_cr_N693), 
	.B2(U_cr_n304), 
	.B1(U_cr_n124), 
	.A2(U_cr_n529), 
	.A1(U_cr_n305));
   AOI22_X2 U_cr_U501 (.ZN(U_cr_n81), 
	.B2(U_cr_n538), 
	.B1(FE_PHN1642_U_cr_n119), 
	.A2(U_cr_n528), 
	.A1(U_cr_n536));
   AOI22_X2 U_cr_U500 (.ZN(U_cr_n82), 
	.B2(U_cr_n538), 
	.B1(U_cr_n110), 
	.A2(FE_OFN332_U_cr_n529), 
	.A1(U_cr_n536));
   AOI22_X2 U_cr_U499 (.ZN(U_cr_N691), 
	.B2(U_cr_n304), 
	.B1(U_cr_n97), 
	.A2(U_cr_n531), 
	.A1(U_cr_n305));
   NOR3_X2 U_cr_U498 (.ZN(U_cr_n429), 
	.A3(U_cr_n315), 
	.A2(hiu_addr[6]), 
	.A1(hiu_haddr[2]));
   INV_X4 U_cr_U497 (.ZN(U_cr_n170), 
	.A(U_cr_n429));
   AOI22_X2 U_cr_U496 (.ZN(U_cr_N639), 
	.B2(U_cr_n288), 
	.B1(U_cr_n113), 
	.A2(FE_OFN336_U_cr_n527), 
	.A1(U_cr_n289));
   AOI22_X2 U_cr_U495 (.ZN(U_cr_n80), 
	.B2(U_cr_n538), 
	.B1(FE_PHN1634_U_cr_n167), 
	.A2(FE_OFN336_U_cr_n527), 
	.A1(U_cr_n536));
   AOI22_X2 U_cr_U494 (.ZN(U_cr_N637), 
	.B2(U_cr_n288), 
	.B1(U_cr_n112), 
	.A2(FE_OFN332_U_cr_n529), 
	.A1(U_cr_n289));
   AOI22_X2 U_cr_U493 (.ZN(U_cr_N694), 
	.B2(U_cr_n304), 
	.B1(U_cr_n125), 
	.A2(FE_OFN333_U_cr_n528), 
	.A1(U_cr_n305));
   AOI22_X2 U_cr_U492 (.ZN(U_cr_N692), 
	.B2(U_cr_n304), 
	.B1(U_cr_n26), 
	.A2(U_cr_n530), 
	.A1(U_cr_n305));
   AOI22_X2 U_cr_U491 (.ZN(U_cr_N737), 
	.B2(U_cr_n312), 
	.B1(U_cr_n164), 
	.A2(U_cr_n530), 
	.A1(U_cr_n313));
   AOI22_X2 U_cr_U490 (.ZN(U_cr_N695), 
	.B2(U_cr_n304), 
	.B1(U_cr_n100), 
	.A2(U_cr_n527), 
	.A1(U_cr_n305));
   AOI22_X2 U_cr_U489 (.ZN(U_cr_N738), 
	.B2(U_cr_n312), 
	.B1(U_cr_n157), 
	.A2(U_cr_n529), 
	.A1(U_cr_n313));
   AOI22_X2 U_cr_U488 (.ZN(U_cr_N638), 
	.B2(U_cr_n288), 
	.B1(U_cr_n121), 
	.A2(U_cr_n528), 
	.A1(U_cr_n289));
   AOI22_X2 U_cr_U487 (.ZN(U_cr_N635), 
	.B2(U_cr_n288), 
	.B1(U_cr_n69), 
	.A2(FE_OFN326_U_cr_n531), 
	.A1(U_cr_n289));
   AOI22_X2 U_cr_U486 (.ZN(U_cr_N739), 
	.B2(U_cr_n312), 
	.B1(U_cr_n158), 
	.A2(FE_OFN333_U_cr_n528), 
	.A1(U_cr_n313));
   AOI22_X2 U_cr_U485 (.ZN(U_cr_N298), 
	.B2(U_cr_n214), 
	.B1(U_cr_n36), 
	.A2(U_cr_n531), 
	.A1(U_cr_n215));
   AOI22_X2 U_cr_U484 (.ZN(U_cr_N302), 
	.B2(U_cr_n214), 
	.B1(FE_PHN1254_U_cr_n55), 
	.A2(U_cr_n527), 
	.A1(U_cr_n215));
   AOI22_X2 U_cr_U483 (.ZN(U_cr_N553), 
	.B2(U_cr_n272), 
	.B1(U_cr_n58), 
	.A2(U_cr_n531), 
	.A1(U_cr_n273));
   AOI22_X2 U_cr_U482 (.ZN(U_cr_N557), 
	.B2(U_cr_n272), 
	.B1(FE_PHN3600_U_cr_n59), 
	.A2(U_cr_n527), 
	.A1(U_cr_n273));
   AOI221_X2 U_cr_U481 (.ZN(U_cr_N550), 
	.C2(U_cr_n272), 
	.C1(U_cr_n56), 
	.B2(U_cr_n273), 
	.B1(U_cr_n514), 
	.A(ctl_init_done));
   INV_X4 U_cr_U480 (.ZN(U_cr_n532), 
	.A(U_cr_n518));
   INV_X4 U_cr_U479 (.ZN(U_cr_n537), 
	.A(U_cr_n514));
   AOI22_X2 U_cr_U478 (.ZN(U_cr_N389), 
	.B2(U_cr_n229), 
	.B1(FE_PHN2455_U_cr_n20), 
	.A2(U_cr_n514), 
	.A1(U_cr_n230));
   AOI22_X2 U_cr_U477 (.ZN(U_cr_N393), 
	.B2(U_cr_n229), 
	.B1(FE_PHN3192_U_cr_n128), 
	.A2(U_cr_n530), 
	.A1(U_cr_n230));
   AOI22_X2 U_cr_U476 (.ZN(U_cr_N395), 
	.B2(U_cr_n229), 
	.B1(FE_PHN3588_U_cr_n149), 
	.A2(U_cr_n528), 
	.A1(U_cr_n230));
   INV_X4 U_cr_U475 (.ZN(U_cr_n171), 
	.A(U_cr_n25));
   INV_X4 U_cr_U474 (.ZN(U_cr_n407), 
	.A(U_cr_n416));
   NOR2_X2 U_cr_U473 (.ZN(U_cr_n321), 
	.A2(U_cr_n359), 
	.A1(U_cr_n316));
   NAND2_X2 U_cr_U472 (.ZN(U_cr_n412), 
	.A2(U_cr_n321), 
	.A1(hiu_haddr[3]));
   AOI21_X2 U_cr_U471 (.ZN(U_cr_n467), 
	.B2(cr_t_wtr[0]), 
	.B1(U_cr_n171), 
	.A(U_cr_n356));
   NAND2_X2 U_cr_U470 (.ZN(U_cr_n176), 
	.A2(big_endian), 
	.A1(U_cr_n318));
   NOR2_X2 U_cr_U469 (.ZN(U_cr_n177), 
	.A2(U_cr_n174), 
	.A1(U_cr_n188));
   NAND3_X2 U_cr_U468 (.ZN(U_cr_n180), 
	.A3(U_cr_n175), 
	.A2(U_cr_n177), 
	.A1(U_cr_n176));
   NOR2_X2 U_cr_U467 (.ZN(U_cr_n497), 
	.A2(big_endian), 
	.A1(U_cr_n182));
   NOR2_X2 U_cr_U466 (.ZN(U_cr_n421), 
	.A2(hiu_haddr[2]), 
	.A1(U_cr_n412));
   INV_X4 U_cr_U465 (.ZN(U_cr_n431), 
	.A(U_cr_n421));
   NAND2_X2 U_cr_U464 (.ZN(U_cr_n465), 
	.A2(U_cr_n431), 
	.A1(U_cr_n357));
   OAI22_X2 U_cr_U463 (.ZN(U_cr_n365), 
	.B2(U_cr_n26), 
	.B1(U_cr_n358), 
	.A2(U_cr_n359), 
	.A1(U_cr_n360));
   AOI22_X2 U_cr_U462 (.ZN(U_cr_n362), 
	.B2(cr_t_ref[4]), 
	.B1(U_cr_n169), 
	.A2(cr_bank_addr_width[1]), 
	.A1(U_cr_n407));
   NAND3_X2 U_cr_U461 (.ZN(U_cr_n364), 
	.A3(U_cr_n361), 
	.A2(U_cr_n362), 
	.A1(U_cr_n363));
   AOI211_X2 U_cr_U460 (.ZN(U_cr_n463), 
	.C2(U_cr_n554), 
	.C1(U_cr_n525), 
	.B(U_cr_n364), 
	.A(U_cr_n365));
   INV_X4 U_cr_U459 (.ZN(U_cr_n469), 
	.A(U_cr_n499));
   AOI22_X2 U_cr_U458 (.ZN(U_cr_n368), 
	.B2(cr_t_wr[0]), 
	.B1(U_cr_n430), 
	.A2(n[23]), 
	.A1(U_cr_n407));
   AOI22_X2 U_cr_U457 (.ZN(U_cr_n367), 
	.B2(cr_t_ref[12]), 
	.B1(U_cr_n169), 
	.A2(U_cr_sctlr_12_), 
	.A1(U_cr_n422));
   NAND3_X2 U_cr_U456 (.ZN(U_cr_n369), 
	.A3(U_cr_n366), 
	.A2(U_cr_n367), 
	.A1(U_cr_n368));
   AOI211_X2 U_cr_U455 (.ZN(U_cr_n462), 
	.C2(cr_t_init[12]), 
	.C1(U_cr_n171), 
	.B(U_cr_n369), 
	.A(U_cr_n421));
   OAI22_X2 U_cr_U454 (.ZN(U_cr_n370), 
	.B2(U_cr_n492), 
	.B1(U_cr_n462), 
	.A2(U_cr_n469), 
	.A1(U_cr_n463));
   AOI21_X2 U_cr_U453 (.ZN(U_cr_n371), 
	.B2(U_cr_n465), 
	.B1(U_cr_n497), 
	.A(U_cr_n370));
   OAI21_X2 U_cr_U452 (.ZN(cr_reg_data_out[12]), 
	.B2(U_cr_n487), 
	.B1(U_cr_n467), 
	.A(U_cr_n371));
   INV_X4 U_cr_U451 (.ZN(U_cr_n485), 
	.A(U_cr_n497));
   OAI22_X2 U_cr_U450 (.ZN(U_cr_n464), 
	.B2(U_cr_n469), 
	.B1(U_cr_n462), 
	.A2(U_cr_n492), 
	.A1(U_cr_n463));
   AOI21_X2 U_cr_U449 (.ZN(U_cr_n466), 
	.B2(U_cr_n465), 
	.B1(U_cr_n204), 
	.A(U_cr_n464));
   OAI21_X2 U_cr_U448 (.ZN(cr_reg_data_out[4]), 
	.B2(U_cr_n485), 
	.B1(U_cr_n467), 
	.A(U_cr_n466));
   AOI22_X2 U_cr_U447 (.ZN(U_cr_N636), 
	.B2(U_cr_n288), 
	.B1(U_cr_n130), 
	.A2(U_cr_n530), 
	.A1(U_cr_n289));
   AOI22_X2 U_cr_U446 (.ZN(U_cr_n84), 
	.B2(U_cr_n538), 
	.B1(FE_PHN3549_U_cr_n165), 
	.A2(FE_OFN326_U_cr_n531), 
	.A1(U_cr_n536));
   AOI22_X2 U_cr_U445 (.ZN(U_cr_n331), 
	.B2(cr_num_init_ref[2]), 
	.B1(U_cr_n171), 
	.A2(gpo[2]), 
	.A1(U_cr_n169));
   AOI21_X2 U_cr_U444 (.ZN(U_cr_n450), 
	.B2(cr_exn_mode_reg_update), 
	.B1(U_cr_n422), 
	.A(U_cr_n333));
   AOI22_X2 U_cr_U443 (.ZN(U_cr_n339), 
	.B2(cr_t_init[10]), 
	.B1(U_cr_n171), 
	.A2(cr_t_ref[10]), 
	.A1(U_cr_n169));
   AOI22_X2 U_cr_U442 (.ZN(U_cr_n338), 
	.B2(cr_t_rp[1]), 
	.B1(U_cr_n430), 
	.A2(n[25]), 
	.A1(U_cr_n407));
   NAND2_X2 U_cr_U441 (.ZN(U_cr_n378), 
	.A2(U_cr_n320), 
	.A1(U_cr_n321));
   AOI211_X2 U_cr_U440 (.ZN(U_cr_n336), 
	.C2(U_cr_n551), 
	.C1(U_cr_n525), 
	.B(U_cr_n335), 
	.A(U_cr_n393));
   NAND4_X2 U_cr_U439 (.ZN(U_cr_n448), 
	.A4(U_cr_n336), 
	.A3(U_cr_n337), 
	.A2(U_cr_n338), 
	.A1(U_cr_n339));
   AOI22_X2 U_cr_U438 (.ZN(U_cr_n342), 
	.B2(cr_t_init[2]), 
	.B1(U_cr_n171), 
	.A2(cr_t_ref[2]), 
	.A1(U_cr_n169));
   NAND3_X2 U_cr_U437 (.ZN(U_cr_n343), 
	.A3(U_cr_n340), 
	.A2(U_cr_n341), 
	.A1(U_cr_n342));
   AOI211_X2 U_cr_U436 (.ZN(U_cr_n446), 
	.C2(U_cr_n556), 
	.C1(U_cr_n525), 
	.B(U_cr_n343), 
	.A(U_cr_n393));
   NOR2_X2 U_cr_U435 (.ZN(U_cr_n392), 
	.A2(U_cr_n412), 
	.A1(U_cr_n320));
   AOI211_X2 U_cr_U434 (.ZN(U_cr_n445), 
	.C2(U_cr_srefr[26]), 
	.C1(U_cr_n169), 
	.B(U_cr_n392), 
	.A(U_cr_n344));
   OAI22_X2 U_cr_U433 (.ZN(U_cr_n345), 
	.B2(U_cr_n485), 
	.B1(U_cr_n445), 
	.A2(U_cr_n469), 
	.A1(U_cr_n446));
   AOI21_X2 U_cr_U432 (.ZN(U_cr_n346), 
	.B2(U_cr_n448), 
	.B1(U_cr_n203), 
	.A(U_cr_n345));
   OAI22_X2 U_cr_U431 (.ZN(U_cr_n447), 
	.B2(U_cr_n487), 
	.B1(U_cr_n445), 
	.A2(U_cr_n492), 
	.A1(U_cr_n446));
   AOI21_X2 U_cr_U430 (.ZN(U_cr_n449), 
	.B2(U_cr_n448), 
	.B1(U_cr_n499), 
	.A(U_cr_n447));
   OAI21_X2 U_cr_U429 (.ZN(cr_reg_data_out[2]), 
	.B2(U_cr_n485), 
	.B1(U_cr_n450), 
	.A(U_cr_n449));
   INV_X4 U_cr_U428 (.ZN(U_cr_n534), 
	.A(U_cr_n516));
   OAI22_X2 U_cr_U427 (.ZN(U_cr_n372), 
	.B2(U_cr_n19), 
	.B1(U_cr_n170), 
	.A2(U_cr_n34), 
	.A1(U_cr_n391));
   AOI211_X2 U_cr_U426 (.ZN(U_cr_n474), 
	.C2(cr_t_wtr[1]), 
	.C1(U_cr_n171), 
	.B(U_cr_n372), 
	.A(U_cr_n421));
   NAND2_X2 U_cr_U425 (.ZN(U_cr_n472), 
	.A2(U_cr_n431), 
	.A1(U_cr_n373));
   NAND2_X2 U_cr_U424 (.ZN(U_cr_n376), 
	.A2(U_cr_n374), 
	.A1(U_cr_n375));
   AOI211_X2 U_cr_U423 (.ZN(U_cr_n470), 
	.C2(cr_t_ref[13]), 
	.C1(U_cr_n169), 
	.B(U_cr_n376), 
	.A(U_cr_n377));
   AOI22_X2 U_cr_U422 (.ZN(U_cr_n379), 
	.B2(cr_exn_mode_value[5]), 
	.B1(U_cr_n423), 
	.A2(cr_t_ras_min[3]), 
	.A1(U_cr_n430));
   NAND4_X2 U_cr_U421 (.ZN(U_cr_n382), 
	.A4(U_cr_n378), 
	.A3(U_cr_n379), 
	.A2(U_cr_n380), 
	.A1(U_cr_n381));
   AOI211_X2 U_cr_U420 (.ZN(U_cr_n468), 
	.C2(cr_ref_all_after_sr), 
	.C1(U_cr_n422), 
	.B(U_cr_n382), 
	.A(U_cr_n383));
   OAI22_X2 U_cr_U419 (.ZN(U_cr_n384), 
	.B2(U_cr_n469), 
	.B1(U_cr_n468), 
	.A2(U_cr_n492), 
	.A1(U_cr_n470));
   AOI21_X2 U_cr_U418 (.ZN(U_cr_n385), 
	.B2(U_cr_n472), 
	.B1(U_cr_n497), 
	.A(U_cr_n384));
   OAI22_X2 U_cr_U417 (.ZN(U_cr_n471), 
	.B2(U_cr_n492), 
	.B1(U_cr_n468), 
	.A2(U_cr_n469), 
	.A1(U_cr_n470));
   AOI21_X2 U_cr_U416 (.ZN(U_cr_n473), 
	.B2(U_cr_n472), 
	.B1(U_cr_n204), 
	.A(U_cr_n471));
   OAI21_X2 U_cr_U415 (.ZN(cr_reg_data_out[5]), 
	.B2(U_cr_n485), 
	.B1(U_cr_n474), 
	.A(U_cr_n473));
   AOI22_X2 U_cr_U414 (.ZN(U_cr_n347), 
	.B2(cr_exn_mode_value[3]), 
	.B1(U_cr_n423), 
	.A2(cr_t_ras_min[1]), 
	.A1(U_cr_n430));
   NAND4_X2 U_cr_U413 (.ZN(U_cr_n350), 
	.A4(U_cr_n378), 
	.A3(U_cr_n347), 
	.A2(U_cr_n348), 
	.A1(U_cr_n349));
   AOI211_X2 U_cr_U412 (.ZN(U_cr_n461), 
	.C2(cr_delayed_precharge), 
	.C1(U_cr_n422), 
	.B(U_cr_n350), 
	.A(U_cr_n351));
   AOI22_X2 U_cr_U411 (.ZN(U_cr_n457), 
	.B2(U_cr_srefr[27]), 
	.B1(U_cr_n169), 
	.A2(cr_t_xsr[4]), 
	.A1(U_cr_n430));
   AOI22_X2 U_cr_U410 (.ZN(U_cr_n442), 
	.B2(U_addrdec_n40), 
	.B1(U_cr_n457), 
	.A2(U_cr_n461), 
	.A1(big_endian));
   AOI22_X2 U_cr_U409 (.ZN(U_cr_n352), 
	.B2(cr_num_init_ref[3]), 
	.B1(U_cr_n171), 
	.A2(U_cr_n572), 
	.A1(U_cr_n422));
   OAI211_X2 U_cr_U408 (.ZN(U_cr_n459), 
	.C2(U_cr_n32), 
	.C1(U_cr_n391), 
	.B(U_cr_n352), 
	.A(U_cr_n353));
   AOI22_X2 U_cr_U407 (.ZN(U_cr_n354), 
	.B2(U_cr_n459), 
	.B1(U_cr_n204), 
	.A2(U_cr_n181), 
	.A1(FE_PHN948_U_cr_n442));
   AOI22_X2 U_cr_U406 (.ZN(U_cr_N470), 
	.B2(U_cr_n267), 
	.B1(U_cr_n135), 
	.A2(U_cr_n528), 
	.A1(U_cr_n268));
   AOI22_X2 U_cr_U405 (.ZN(U_cr_N468), 
	.B2(U_cr_n267), 
	.B1(U_cr_n134), 
	.A2(U_cr_n530), 
	.A1(U_cr_n268));
   AOI22_X2 U_cr_U404 (.ZN(U_cr_N471), 
	.B2(U_cr_n267), 
	.B1(U_cr_n142), 
	.A2(U_cr_n527), 
	.A1(U_cr_n268));
   AOI22_X2 U_cr_U403 (.ZN(U_cr_N469), 
	.B2(U_cr_n267), 
	.B1(U_cr_n141), 
	.A2(U_cr_n529), 
	.A1(U_cr_n268));
   AOI22_X2 U_cr_U402 (.ZN(U_cr_N467), 
	.B2(U_cr_n267), 
	.B1(U_cr_n150), 
	.A2(U_cr_n531), 
	.A1(U_cr_n268));
   OAI22_X2 U_cr_U401 (.ZN(U_cr_n458), 
	.B2(U_cr_n469), 
	.B1(U_cr_n456), 
	.A2(U_cr_n487), 
	.A1(U_cr_n457));
   AOI21_X2 U_cr_U400 (.ZN(U_cr_n460), 
	.B2(U_cr_n459), 
	.B1(U_cr_n497), 
	.A(U_cr_n458));
   AOI221_X2 U_cr_U399 (.ZN(U_cr_n216), 
	.C2(ad_cr_data_mask[1]), 
	.C1(U_addrdec_n40), 
	.B2(ad_cr_data_mask[2]), 
	.B1(big_endian), 
	.A(U_cr_n205));
   NOR2_X2 U_cr_U398 (.ZN(U_cr_n275), 
	.A2(U_cr_n544), 
	.A1(U_cr_n396));
   INV_X4 U_cr_U397 (.ZN(U_cr_n274), 
	.A(U_cr_n275));
   AOI22_X2 U_cr_U396 (.ZN(U_cr_N563), 
	.B2(U_cr_n274), 
	.B1(U_cr_n35), 
	.A2(U_cr_n291), 
	.A1(U_cr_n275));
   AOI22_X2 U_cr_U395 (.ZN(U_cr_N564), 
	.B2(U_cr_n274), 
	.B1(FE_PHN3107_U_cr_n44), 
	.A2(U_cr_n293), 
	.A1(U_cr_n275));
   AOI22_X2 U_cr_U394 (.ZN(U_cr_N558), 
	.B2(U_cr_n274), 
	.B1(U_cr_n41), 
	.A2(U_cr_n548), 
	.A1(U_cr_n275));
   AOI22_X2 U_cr_U393 (.ZN(U_cr_N560), 
	.B2(U_cr_n274), 
	.B1(U_cr_n155), 
	.A2(U_cr_n545), 
	.A1(U_cr_n275));
   AOI221_X2 U_cr_U392 (.ZN(U_cr_N559), 
	.C2(U_cr_n274), 
	.C1(U_cr_n61), 
	.B2(U_cr_n275), 
	.B1(U_cr_n546), 
	.A(ctl_mode_reg_done));
   AOI22_X2 U_cr_U391 (.ZN(U_cr_n517), 
	.B2(FE_OFN357_U_addrdec_n40), 
	.B1(hiu_wr_data[18]), 
	.A2(hiu_wr_data[10]), 
	.A1(U_cr_n168));
   NAND2_X2 U_cr_U390 (.ZN(U_cr_n512), 
	.A2(U_cr_n240), 
	.A1(U_cr_n223));
   NOR2_X2 U_cr_U389 (.ZN(U_cr_n506), 
	.A2(U_cr_n512), 
	.A1(U_cr_n396));
   INV_X4 U_cr_U388 (.ZN(U_cr_n508), 
	.A(U_cr_n506));
   NAND2_X2 U_cr_U387 (.ZN(U_cr_n276), 
	.A2(U_cr_n223), 
	.A1(U_cr_n238));
   NOR2_X2 U_cr_U386 (.ZN(U_cr_n279), 
	.A2(U_cr_n396), 
	.A1(U_cr_n276));
   AOI22_X2 U_cr_U385 (.ZN(U_cr_n281), 
	.B2(U_cr_n532), 
	.B1(U_cr_n279), 
	.A2(U_cr_n508), 
	.A1(cr_exn_mode_reg_update));
   NAND2_X2 U_cr_U384 (.ZN(U_cr_n280), 
	.A2(U_cr_n511), 
	.A1(U_cr_n422));
   AOI221_X2 U_cr_U383 (.ZN(U_cr_N567), 
	.C2(U_cr_n281), 
	.C1(U_cr_n280), 
	.B2(U_cr_n281), 
	.B1(U_cr_n517), 
	.A(ctl_ext_mode_reg_done));
   NAND4_X2 U_cr_U382 (.ZN(U_cr_n495), 
	.A4(U_cr_n408), 
	.A3(U_cr_n409), 
	.A2(U_cr_n410), 
	.A1(U_cr_n411));
   NAND2_X2 U_cr_U381 (.ZN(U_cr_n453), 
	.A2(big_endian), 
	.A1(U_cr_n13));
   AOI21_X2 U_cr_U380 (.ZN(U_cr_n415), 
	.B2(cr_s_ready_valid), 
	.B1(U_cr_n422), 
	.A(U_cr_n414));
   OAI21_X2 U_cr_U379 (.ZN(U_cr_n494), 
	.B2(U_cr_n31), 
	.B1(U_cr_n416), 
	.A(U_cr_n415));
   NAND2_X2 U_cr_U378 (.ZN(U_cr_n451), 
	.A2(U_addrdec_n40), 
	.A1(U_cr_n13));
   OAI22_X2 U_cr_U377 (.ZN(cr_reg_data_out[17]), 
	.B2(U_cr_n451), 
	.B1(U_cr_n417), 
	.A2(U_cr_n453), 
	.A1(U_cr_n418));
   AOI22_X2 U_cr_U376 (.ZN(U_cr_n484), 
	.B2(U_cr_srefr[31]), 
	.B1(U_cr_n429), 
	.A2(cr_t_xsr[8]), 
	.A1(U_cr_n430));
   NAND4_X2 U_cr_U375 (.ZN(U_cr_n481), 
	.A4(U_cr_n399), 
	.A3(U_cr_n400), 
	.A2(U_cr_n401), 
	.A1(U_cr_n402));
   AOI22_X2 U_cr_U374 (.ZN(U_cr_n405), 
	.B2(cr_t_ref[15]), 
	.B1(U_cr_n169), 
	.A2(s_sa[0]), 
	.A1(U_cr_n407));
   NAND2_X2 U_cr_U373 (.ZN(U_cr_n406), 
	.A2(U_cr_n404), 
	.A1(U_cr_n405));
   AOI21_X2 U_cr_U372 (.ZN(U_cr_n438), 
	.B2(U_cr_n422), 
	.B1(U_cr_sctlr_15_), 
	.A(U_cr_n406));
   AOI22_X2 U_cr_U371 (.ZN(U_cr_n437), 
	.B2(gpo[7]), 
	.B1(U_cr_n169), 
	.A2(cr_t_rc[1]), 
	.A1(U_cr_n430));
   AOI22_X2 U_cr_U370 (.ZN(U_cr_n482), 
	.B2(U_addrdec_n40), 
	.B1(U_cr_n437), 
	.A2(U_cr_n438), 
	.A1(big_endian));
   AOI22_X2 U_cr_U369 (.ZN(U_cr_n483), 
	.B2(FE_PHN1163_U_cr_n482), 
	.B1(U_cr_n181), 
	.A2(U_cr_n203), 
	.A1(U_cr_n481));
   AOI22_X2 U_cr_U368 (.ZN(U_cr_n513), 
	.B2(FE_OFN357_U_addrdec_n40), 
	.B1(hiu_wr_data[16]), 
	.A2(U_cr_n168), 
	.A1(hiu_wr_data[8]));
   AOI22_X2 U_cr_U367 (.ZN(U_cr_n277), 
	.B2(U_cr_n508), 
	.B1(U_cr_sctlr_16_), 
	.A2(U_cr_n537), 
	.A1(U_cr_n279));
   OAI21_X2 U_cr_U366 (.ZN(U_cr_N565), 
	.B2(U_cr_n280), 
	.B1(U_cr_n513), 
	.A(U_cr_n277));
   AOI22_X2 U_cr_U365 (.ZN(U_cr_n515), 
	.B2(FE_OFN357_U_addrdec_n40), 
	.B1(hiu_wr_data[17]), 
	.A2(U_cr_n168), 
	.A1(hiu_wr_data[9]));
   AOI22_X2 U_cr_U364 (.ZN(U_cr_n278), 
	.B2(U_cr_n508), 
	.B1(cr_s_ready_valid), 
	.A2(U_cr_n534), 
	.A1(U_cr_n279));
   OAI21_X2 U_cr_U363 (.ZN(U_cr_N566), 
	.B2(U_cr_n280), 
	.B1(U_cr_n515), 
	.A(U_cr_n278));
   AOI22_X2 U_cr_U362 (.ZN(U_cr_n519), 
	.B2(U_addrdec_n40), 
	.B1(hiu_wr_data[19]), 
	.A2(U_cr_n168), 
	.A1(hiu_wr_data[11]));
   OAI22_X2 U_cr_U361 (.ZN(U_cr_n509), 
	.B2(U_cr_n506), 
	.B1(U_cr_n572), 
	.A2(U_cr_n507), 
	.A1(U_cr_n508));
   INV_X4 U_cr_U360 (.ZN(U_cr_n73), 
	.A(U_cr_n509));
   AOI22_X2 U_cr_U359 (.ZN(U_cr_n455), 
	.B2(U_addrdec_n40), 
	.B1(U_cr_n403), 
	.A2(U_cr_n481), 
	.A1(big_endian));
   AOI22_X2 U_cr_U358 (.ZN(U_cr_N561), 
	.B2(U_cr_n274), 
	.B1(FE_PHN2051_U_cr_n18), 
	.A2(FE_OFN0_U_cr_n314), 
	.A1(U_cr_n275));
   AOI22_X2 U_cr_U357 (.ZN(U_cr_N562), 
	.B2(U_cr_n274), 
	.B1(FE_PHN1473_U_cr_n27), 
	.A2(U_cr_n290), 
	.A1(U_cr_n275));
   AOI21_X2 U_cr_U356 (.ZN(U_cr_n323), 
	.B2(U_cr_n422), 
	.B1(cr_do_initialize), 
	.A(U_cr_n393));
   NAND4_X2 U_cr_U355 (.ZN(U_cr_n490), 
	.A4(U_cr_n322), 
	.A3(U_cr_n323), 
	.A2(U_cr_n324), 
	.A1(U_cr_n325));
   AOI22_X2 U_cr_U354 (.ZN(U_cr_n326), 
	.B2(cr_num_init_ref[0]), 
	.B1(U_cr_n171), 
	.A2(gpo[0]), 
	.A1(U_cr_n169));
   AOI21_X2 U_cr_U353 (.ZN(U_cr_n488), 
	.B2(U_cr_sctlr_16_), 
	.B1(U_cr_n422), 
	.A(U_cr_n328));
   OAI22_X2 U_cr_U352 (.ZN(U_cr_n489), 
	.B2(U_cr_n485), 
	.B1(U_cr_n486), 
	.A2(U_cr_n487), 
	.A1(U_cr_n488));
   AOI21_X2 U_cr_U351 (.ZN(U_cr_n491), 
	.B2(U_cr_n490), 
	.B1(U_cr_n499), 
	.A(U_cr_n489));
   OAI22_X2 U_cr_U350 (.ZN(U_cr_n329), 
	.B2(U_cr_n487), 
	.B1(U_cr_n486), 
	.A2(U_cr_n485), 
	.A1(U_cr_n488));
   AOI21_X2 U_cr_U349 (.ZN(U_cr_n330), 
	.B2(U_cr_n490), 
	.B1(U_cr_n203), 
	.A(U_cr_n329));
   OAI21_X2 U_cr_U348 (.ZN(cr_reg_data_out[0]), 
	.B2(U_cr_n469), 
	.B1(U_cr_n493), 
	.A(U_cr_n330));
   INV_X4 U_cr_U347 (.ZN(U_cr_n220), 
	.A(U_cr_n221));
   AOI22_X2 U_cr_U346 (.ZN(U_cr_N306), 
	.B2(U_cr_n220), 
	.B1(U_cr_n38), 
	.A2(FE_OFN1_U_cr_n541), 
	.A1(U_cr_n221));
   AOI22_X2 U_cr_U345 (.ZN(U_cr_N310), 
	.B2(U_cr_n220), 
	.B1(U_cr_n52), 
	.A2(U_cr_n293), 
	.A1(U_cr_n221));
   INV_X4 U_cr_U344 (.ZN(U_cr_n510), 
	.A(U_cr_n276));
   NAND2_X2 U_cr_U343 (.ZN(U_cr_n233), 
	.A2(U_cr_n430), 
	.A1(U_cr_n510));
   NAND2_X2 U_cr_U342 (.ZN(U_cr_n235), 
	.A2(U_cr_n430), 
	.A1(U_cr_n511));
   NOR2_X2 U_cr_U341 (.ZN(U_cr_n234), 
	.A2(U_cr_n391), 
	.A1(U_cr_n512));
   OAI222_X2 U_cr_U340 (.ZN(U_cr_N408), 
	.C2(U_cr_n234), 
	.C1(U_cr_n32), 
	.B2(U_cr_n519), 
	.B1(U_cr_n235), 
	.A2(U_cr_n531), 
	.A1(U_cr_n233));
   AOI22_X2 U_cr_U339 (.ZN(U_cr_n295), 
	.B2(FE_OFN357_U_addrdec_n40), 
	.B1(hiu_wr_data[22]), 
	.A2(U_cr_n168), 
	.A1(hiu_wr_data[14]));
   OAI222_X2 U_cr_U338 (.ZN(U_cr_N411), 
	.C2(U_cr_n528), 
	.C1(U_cr_n233), 
	.B2(U_cr_n234), 
	.B1(FE_OFN23_U_cr_n64), 
	.A2(FE_PHN1015_U_cr_n295), 
	.A1(U_cr_n235));
   OAI222_X2 U_cr_U337 (.ZN(U_cr_N405), 
	.C2(U_cr_n234), 
	.C1(FE_PHN1407_U_cr_n104), 
	.B2(U_cr_n513), 
	.B1(U_cr_n235), 
	.A2(U_cr_n514), 
	.A1(U_cr_n233));
   AOI22_X2 U_cr_U336 (.ZN(U_cr_N305), 
	.B2(U_cr_n220), 
	.B1(U_cr_n22), 
	.A2(U_cr_n545), 
	.A1(U_cr_n221));
   AOI22_X2 U_cr_U335 (.ZN(U_cr_N304), 
	.B2(U_cr_n220), 
	.B1(FE_PHN3113_U_cr_n63), 
	.A2(U_cr_n546), 
	.A1(U_cr_n221));
   AOI22_X2 U_cr_U334 (.ZN(U_cr_N303), 
	.B2(U_cr_n220), 
	.B1(U_cr_n70), 
	.A2(U_cr_n548), 
	.A1(U_cr_n221));
   AOI22_X2 U_cr_U333 (.ZN(U_cr_N307), 
	.B2(U_cr_n220), 
	.B1(FE_PHN1645_U_cr_n65), 
	.A2(FE_OFN0_U_cr_n314), 
	.A1(U_cr_n221));
   NAND2_X2 U_cr_U332 (.ZN(U_cr_n299), 
	.A2(U_cr_n169), 
	.A1(U_cr_n510));
   NAND2_X2 U_cr_U331 (.ZN(U_cr_n298), 
	.A2(U_cr_n169), 
	.A1(U_cr_n511));
   NOR2_X2 U_cr_U330 (.ZN(U_cr_n296), 
	.A2(U_cr_n170), 
	.A1(U_cr_n512));
   OAI222_X2 U_cr_U329 (.ZN(U_cr_N651), 
	.C2(U_cr_n296), 
	.C1(FE_PHN4855_U_cr_n49), 
	.B2(U_cr_n519), 
	.B1(U_cr_n298), 
	.A2(U_cr_n531), 
	.A1(U_cr_n299));
   AOI22_X2 U_cr_U328 (.ZN(U_cr_n520), 
	.B2(FE_OFN357_U_addrdec_n40), 
	.B1(hiu_wr_data[20]), 
	.A2(U_cr_n168), 
	.A1(hiu_wr_data[12]));
   OAI222_X2 U_cr_U327 (.ZN(U_cr_N652), 
	.C2(U_cr_n296), 
	.C1(FE_PHN4798_U_cr_n50), 
	.B2(U_cr_n520), 
	.B1(U_cr_n298), 
	.A2(U_cr_n530), 
	.A1(U_cr_n299));
   AOI22_X2 U_cr_U326 (.ZN(U_cr_n522), 
	.B2(FE_OFN357_U_addrdec_n40), 
	.B1(hiu_wr_data[21]), 
	.A2(U_cr_n168), 
	.A1(hiu_wr_data[13]));
   OAI222_X2 U_cr_U325 (.ZN(U_cr_N410), 
	.C2(U_cr_n529), 
	.C1(U_cr_n233), 
	.B2(U_cr_n234), 
	.B1(U_cr_n34), 
	.A2(U_cr_n522), 
	.A1(U_cr_n235));
   AOI22_X2 U_cr_U324 (.ZN(U_cr_n297), 
	.B2(FE_OFN357_U_addrdec_n40), 
	.B1(hiu_wr_data[23]), 
	.A2(U_cr_n168), 
	.A1(hiu_wr_data[15]));
   OAI222_X2 U_cr_U323 (.ZN(U_cr_N412), 
	.C2(U_cr_n527), 
	.C1(U_cr_n233), 
	.B2(U_cr_n234), 
	.B1(U_cr_n106), 
	.A2(FE_PHN1171_U_cr_n297), 
	.A1(U_cr_n235));
   OAI222_X2 U_cr_U322 (.ZN(U_cr_N653), 
	.C2(U_cr_n296), 
	.C1(FE_PHN4464_U_cr_n19), 
	.B2(U_cr_n522), 
	.B1(U_cr_n298), 
	.A2(U_cr_n529), 
	.A1(U_cr_n299));
   OAI222_X2 U_cr_U321 (.ZN(U_cr_N409), 
	.C2(U_cr_n234), 
	.C1(U_cr_n33), 
	.B2(U_cr_n520), 
	.B1(U_cr_n235), 
	.A2(U_cr_n530), 
	.A1(U_cr_n233));
   OAI222_X2 U_cr_U320 (.ZN(U_cr_N655), 
	.C2(U_cr_n296), 
	.C1(FE_PHN4915_U_cr_n51), 
	.B2(FE_PHN1171_U_cr_n297), 
	.B1(U_cr_n298), 
	.A2(U_cr_n527), 
	.A1(U_cr_n299));
   OAI222_X2 U_cr_U319 (.ZN(U_cr_N654), 
	.C2(U_cr_n296), 
	.C1(FE_PHN4871_U_cr_n46), 
	.B2(FE_PHN1015_U_cr_n295), 
	.B1(U_cr_n298), 
	.A2(U_cr_n528), 
	.A1(U_cr_n299));
   OAI222_X2 U_cr_U318 (.ZN(U_cr_N649), 
	.C2(U_cr_n296), 
	.C1(FE_PHN4265_U_cr_n29), 
	.B2(U_cr_n515), 
	.B1(U_cr_n298), 
	.A2(U_cr_n516), 
	.A1(U_cr_n299));
   OAI222_X2 U_cr_U317 (.ZN(U_cr_N648), 
	.C2(U_cr_n296), 
	.C1(FE_PHN4845_U_cr_n47), 
	.B2(U_cr_n513), 
	.B1(U_cr_n298), 
	.A2(U_cr_n514), 
	.A1(U_cr_n299));
   INV_X4 U_cr_U316 (.ZN(U_cr_n306), 
	.A(U_cr_n307));
   AOI22_X2 U_cr_U315 (.ZN(U_cr_N697), 
	.B2(U_cr_n306), 
	.B1(U_cr_n101), 
	.A2(U_cr_n546), 
	.A1(U_cr_n307));
   INV_X4 U_cr_U314 (.ZN(U_cr_n540), 
	.A(U_cr_n542));
   AOI22_X2 U_cr_U313 (.ZN(U_cr_n91), 
	.B2(U_cr_n540), 
	.B1(U_cr_n163), 
	.A2(FE_OFN1_U_cr_n541), 
	.A1(U_cr_n542));
   AOI22_X2 U_cr_U312 (.ZN(U_cr_N698), 
	.B2(U_cr_n306), 
	.B1(U_cr_n71), 
	.A2(U_cr_n545), 
	.A1(U_cr_n307));
   AOI22_X2 U_cr_U311 (.ZN(U_cr_N699), 
	.B2(U_cr_n306), 
	.B1(U_cr_n102), 
	.A2(FE_OFN1_U_cr_n541), 
	.A1(U_cr_n307));
   AOI22_X2 U_cr_U310 (.ZN(U_cr_N696), 
	.B2(U_cr_n306), 
	.B1(U_cr_n126), 
	.A2(U_cr_n548), 
	.A1(U_cr_n307));
   AOI22_X2 U_cr_U309 (.ZN(U_cr_n89), 
	.B2(U_cr_n540), 
	.B1(U_cr_n162), 
	.A2(U_cr_n546), 
	.A1(U_cr_n542));
   AOI22_X2 U_cr_U308 (.ZN(U_cr_n90), 
	.B2(U_cr_n540), 
	.B1(U_cr_n37), 
	.A2(U_cr_n545), 
	.A1(U_cr_n542));
   AOI22_X2 U_cr_U307 (.ZN(U_cr_N700), 
	.B2(U_cr_n306), 
	.B1(U_cr_n103), 
	.A2(FE_OFN0_U_cr_n314), 
	.A1(U_cr_n307));
   AOI22_X2 U_cr_U306 (.ZN(U_cr_n88), 
	.B2(U_cr_n540), 
	.B1(U_cr_n161), 
	.A2(U_cr_n548), 
	.A1(U_cr_n542));
   AOI22_X2 U_cr_U305 (.ZN(U_cr_N745), 
	.B2(U_cr_n540), 
	.B1(U_cr_n160), 
	.A2(FE_OFN0_U_cr_n314), 
	.A1(U_cr_n542));
   OAI222_X2 U_cr_U304 (.ZN(U_cr_N406), 
	.C2(U_cr_n234), 
	.C1(U_cr_n72), 
	.B2(U_cr_n515), 
	.B1(U_cr_n235), 
	.A2(U_cr_n516), 
	.A1(U_cr_n233));
   OAI222_X2 U_cr_U303 (.ZN(U_cr_N650), 
	.C2(U_cr_n296), 
	.C1(FE_PHN4894_U_cr_n48), 
	.B2(U_cr_n517), 
	.B1(U_cr_n298), 
	.A2(U_cr_n518), 
	.A1(U_cr_n299));
   NAND2_X2 U_cr_U302 (.ZN(U_cr_n226), 
	.A2(U_cr_n407), 
	.A1(U_cr_n511));
   NOR2_X2 U_cr_U301 (.ZN(U_cr_n225), 
	.A2(U_cr_n416), 
	.A1(U_cr_n512));
   NAND2_X2 U_cr_U300 (.ZN(U_cr_n224), 
	.A2(U_cr_n407), 
	.A1(U_cr_n510));
   AOI22_X2 U_cr_U298 (.ZN(U_cr_n434), 
	.B2(U_cr_n494), 
	.B1(U_cr_n497), 
	.A2(U_cr_n495), 
	.A1(U_cr_n499));
   NAND4_X2 U_cr_U297 (.ZN(U_cr_n498), 
	.A4(U_cr_n425), 
	.A3(U_cr_n426), 
	.A2(U_cr_n427), 
	.A1(U_cr_n428));
   NAND2_X2 U_cr_U296 (.ZN(U_cr_n496), 
	.A2(U_cr_n431), 
	.A1(U_cr_n432));
   AOI22_X2 U_cr_U295 (.ZN(U_cr_n433), 
	.B2(U_cr_n496), 
	.B1(U_cr_n204), 
	.A2(U_cr_n498), 
	.A1(U_cr_n203));
   NAND2_X2 U_cr_U294 (.ZN(cr_reg_data_out[1]), 
	.A2(U_cr_n433), 
	.A1(U_cr_n434));
   AOI22_X2 U_cr_U293 (.ZN(U_cr_n501), 
	.B2(U_cr_n494), 
	.B1(U_cr_n204), 
	.A2(U_cr_n495), 
	.A1(U_cr_n203));
   AOI22_X2 U_cr_U292 (.ZN(U_cr_n500), 
	.B2(U_cr_n496), 
	.B1(U_cr_n497), 
	.A2(U_cr_n498), 
	.A1(U_cr_n499));
   NAND2_X2 U_cr_U291 (.ZN(cr_reg_data_out[9]), 
	.A2(U_cr_n500), 
	.A1(U_cr_n501));
   OAI222_X2 U_cr_U290 (.ZN(U_cr_N315), 
	.C2(U_cr_n530), 
	.C1(U_cr_n224), 
	.B2(U_cr_n225), 
	.B1(U_cr_n57), 
	.A2(U_cr_n520), 
	.A1(U_cr_n226));
   OAI222_X2 U_cr_U289 (.ZN(U_cr_N407), 
	.C2(U_cr_n234), 
	.C1(FE_PHN4952_U_cr_n108), 
	.B2(U_cr_n517), 
	.B1(U_cr_n235), 
	.A2(U_cr_n518), 
	.A1(U_cr_n233));
   NAND2_X2 U_cr_U288 (.ZN(U_cr_n524), 
	.A2(U_cr_n171), 
	.A1(U_cr_n510));
   NAND2_X2 U_cr_U287 (.ZN(U_cr_n523), 
	.A2(U_cr_n171), 
	.A1(U_cr_n511));
   NOR2_X2 U_cr_U286 (.ZN(U_cr_n521), 
	.A2(U_cr_n25), 
	.A1(U_cr_n512));
   OAI222_X2 U_cr_U285 (.ZN(U_cr_n75), 
	.C2(U_cr_n521), 
	.C1(U_cr_n117), 
	.B2(U_cr_n515), 
	.B1(U_cr_n523), 
	.A2(U_cr_n516), 
	.A1(U_cr_n524));
   OAI222_X2 U_cr_U284 (.ZN(U_cr_n74), 
	.C2(U_cr_n521), 
	.C1(U_cr_n115), 
	.B2(U_cr_n513), 
	.B1(U_cr_n523), 
	.A2(U_cr_n514), 
	.A1(U_cr_n524));
   AOI22_X2 U_cr_U283 (.ZN(U_cr_N644), 
	.B2(U_cr_n292), 
	.B1(U_cr_n122), 
	.A2(FE_OFN0_U_cr_n314), 
	.A1(U_cr_n294));
   AOI22_X2 U_cr_U282 (.ZN(U_cr_N476), 
	.B2(U_cr_n269), 
	.B1(U_cr_n131), 
	.A2(FE_OFN0_U_cr_n314), 
	.A1(U_cr_n270));
   AOI22_X2 U_cr_U281 (.ZN(U_cr_N646), 
	.B2(U_cr_n292), 
	.B1(U_cr_n123), 
	.A2(U_cr_n291), 
	.A1(U_cr_n294));
   AOI22_X2 U_cr_U280 (.ZN(U_cr_N647), 
	.B2(U_cr_n292), 
	.B1(U_cr_n114), 
	.A2(U_cr_n293), 
	.A1(U_cr_n294));
   AOI22_X2 U_cr_U279 (.ZN(U_cr_N474), 
	.B2(U_cr_n269), 
	.B1(U_cr_n137), 
	.A2(U_cr_n545), 
	.A1(U_cr_n270));
   AOI22_X2 U_cr_U278 (.ZN(U_cr_N643), 
	.B2(U_cr_n292), 
	.B1(U_cr_n111), 
	.A2(FE_OFN1_U_cr_n541), 
	.A1(U_cr_n294));
   AOI22_X2 U_cr_U277 (.ZN(U_cr_N477), 
	.B2(U_cr_n269), 
	.B1(U_cr_n145), 
	.A2(FE_OFN347_U_cr_n290), 
	.A1(U_cr_n270));
   AOI22_X2 U_cr_U276 (.ZN(U_cr_N402), 
	.B2(U_cr_n231), 
	.B1(U_cr_n67), 
	.A2(U_cr_n290), 
	.A1(U_cr_n232));
   AOI22_X2 U_cr_U275 (.ZN(U_cr_N473), 
	.B2(U_cr_n269), 
	.B1(U_cr_n143), 
	.A2(U_cr_n546), 
	.A1(U_cr_n270));
   AOI22_X2 U_cr_U274 (.ZN(U_cr_N641), 
	.B2(U_cr_n292), 
	.B1(U_cr_n105), 
	.A2(U_cr_n546), 
	.A1(U_cr_n294));
   AOI22_X2 U_cr_U273 (.ZN(U_cr_N398), 
	.B2(U_cr_n231), 
	.B1(FE_PHN3505_U_cr_n45), 
	.A2(U_cr_n546), 
	.A1(U_cr_n232));
   AOI22_X2 U_cr_U272 (.ZN(U_cr_N475), 
	.B2(U_cr_n269), 
	.B1(U_cr_n144), 
	.A2(FE_OFN1_U_cr_n541), 
	.A1(U_cr_n270));
   AOI22_X2 U_cr_U271 (.ZN(U_cr_N397), 
	.B2(U_cr_n231), 
	.B1(U_cr_n140), 
	.A2(U_cr_n548), 
	.A1(U_cr_n232));
   AOI22_X2 U_cr_U270 (.ZN(U_cr_N640), 
	.B2(U_cr_n292), 
	.B1(U_cr_n118), 
	.A2(U_cr_n548), 
	.A1(U_cr_n294));
   AOI22_X2 U_cr_U269 (.ZN(U_cr_N472), 
	.B2(U_cr_n269), 
	.B1(U_cr_n136), 
	.A2(U_cr_n548), 
	.A1(U_cr_n270));
   AOI22_X2 U_cr_U268 (.ZN(U_cr_N478), 
	.B2(U_cr_n269), 
	.B1(U_cr_n138), 
	.A2(FE_OFN345_U_cr_n291), 
	.A1(U_cr_n270));
   AOI22_X2 U_cr_U267 (.ZN(U_cr_N400), 
	.B2(U_cr_n231), 
	.B1(FE_PHN3514_U_cr_n148), 
	.A2(FE_OFN1_U_cr_n541), 
	.A1(U_cr_n232));
   AOI22_X2 U_cr_U266 (.ZN(U_cr_N479), 
	.B2(U_cr_n269), 
	.B1(U_cr_n146), 
	.A2(U_cr_n293), 
	.A1(U_cr_n270));
   AOI22_X2 U_cr_U265 (.ZN(U_cr_N645), 
	.B2(U_cr_n292), 
	.B1(U_cr_n68), 
	.A2(U_cr_n290), 
	.A1(U_cr_n294));
   OAI222_X2 U_cr_U264 (.ZN(U_cr_n76), 
	.C2(U_cr_n521), 
	.C1(U_cr_n116), 
	.B2(U_cr_n517), 
	.B1(U_cr_n523), 
	.A2(U_cr_n518), 
	.A1(U_cr_n524));
   OAI222_X2 U_cr_U263 (.ZN(U_cr_n77), 
	.C2(U_cr_n521), 
	.C1(U_cr_n109), 
	.B2(U_cr_n519), 
	.B1(U_cr_n523), 
	.A2(U_cr_n531), 
	.A1(U_cr_n524));
   OAI222_X2 U_cr_U262 (.ZN(U_cr_n78), 
	.C2(U_cr_n521), 
	.C1(FE_PHN4110_U_cr_n53), 
	.B2(U_cr_n520), 
	.B1(U_cr_n523), 
	.A2(U_cr_n530), 
	.A1(U_cr_n524));
   OAI222_X2 U_cr_U261 (.ZN(U_cr_n79), 
	.C2(U_cr_n521), 
	.C1(FE_PHN3988_U_cr_n60), 
	.B2(U_cr_n522), 
	.B1(U_cr_n523), 
	.A2(U_cr_n529), 
	.A1(U_cr_n524));
   OAI22_X2 U_cr_U260 (.ZN(cr_reg_data_out[16]), 
	.B2(U_cr_n453), 
	.B1(U_cr_n493), 
	.A2(U_cr_n451), 
	.A1(U_cr_n488));
   OAI222_X2 U_cr_U259 (.ZN(U_cr_N313), 
	.C2(U_cr_n225), 
	.C1(U_cr_n30), 
	.B2(U_cr_n517), 
	.B1(U_cr_n226), 
	.A2(U_cr_n518), 
	.A1(U_cr_n224));
   NOR2_X2 U_cr_U258 (.ZN(U_cr_n549), 
	.A2(U_cr_n543), 
	.A1(U_cr_n544));
   INV_X4 U_cr_U257 (.ZN(U_cr_n547), 
	.A(U_cr_n549));
   AOI22_X2 U_cr_U256 (.ZN(U_cr_n94), 
	.B2(U_cr_n547), 
	.B1(U_cr_n154), 
	.A2(FE_OFN319_U_cr_n548), 
	.A1(U_cr_n549));
   AOI22_X2 U_cr_U255 (.ZN(U_cr_n92), 
	.B2(U_cr_n547), 
	.B1(U_cr_n153), 
	.A2(U_cr_n545), 
	.A1(U_cr_n549));
   AOI22_X2 U_cr_U254 (.ZN(U_cr_N404), 
	.B2(U_cr_n231), 
	.B1(FE_PHN1482_U_cr_n151), 
	.A2(U_cr_n293), 
	.A1(U_cr_n232));
   AOI22_X2 U_cr_U253 (.ZN(U_cr_N403), 
	.B2(U_cr_n231), 
	.B1(FE_PHN1052_U_cr_n127), 
	.A2(U_cr_n291), 
	.A1(U_cr_n232));
   AOI22_X2 U_cr_U252 (.ZN(U_cr_N401), 
	.B2(U_cr_n231), 
	.B1(U_cr_n107), 
	.A2(FE_OFN0_U_cr_n314), 
	.A1(U_cr_n232));
   AOI22_X2 U_cr_U251 (.ZN(U_cr_N642), 
	.B2(U_cr_n292), 
	.B1(U_cr_n129), 
	.A2(U_cr_n545), 
	.A1(U_cr_n294));
   AOI22_X2 U_cr_U250 (.ZN(U_cr_N399), 
	.B2(U_cr_n231), 
	.B1(FE_PHN3012_U_cr_n147), 
	.A2(U_cr_n545), 
	.A1(U_cr_n232));
   OAI222_X2 U_cr_U249 (.ZN(U_cr_N311), 
	.C2(U_cr_n225), 
	.C1(U_cr_n28), 
	.B2(U_cr_n513), 
	.B1(U_cr_n226), 
	.A2(U_cr_n514), 
	.A1(U_cr_n224));
   OAI22_X2 U_cr_U248 (.ZN(cr_reg_data_out[26]), 
	.B2(U_cr_n453), 
	.B1(U_cr_n446), 
	.A2(U_cr_n451), 
	.A1(U_cr_n445));
   OAI22_X2 U_cr_U247 (.ZN(cr_reg_data_out[18]), 
	.B2(U_cr_n451), 
	.B1(U_cr_n450), 
	.A2(U_cr_n453), 
	.A1(U_cr_n419));
   OAI222_X2 U_cr_U246 (.ZN(U_cr_N312), 
	.C2(U_cr_n225), 
	.C1(U_cr_n31), 
	.B2(U_cr_n516), 
	.B1(U_cr_n224), 
	.A2(U_cr_n515), 
	.A1(U_cr_n226));
   AOI21_X2 U_cr_U245 (.ZN(U_cr_n395), 
	.B2(cr_t_ref[14]), 
	.B1(U_cr_n169), 
	.A(U_cr_n393));
   OAI211_X2 U_cr_U244 (.ZN(U_cr_n478), 
	.C2(U_cr_n35), 
	.C1(U_cr_n396), 
	.B(U_cr_n394), 
	.A(U_cr_n395));
   OAI22_X2 U_cr_U243 (.ZN(cr_reg_data_out[22]), 
	.B2(U_cr_n453), 
	.B1(U_cr_n435), 
	.A2(U_cr_n451), 
	.A1(U_cr_n436));
   AOI22_X2 U_cr_U242 (.ZN(U_cr_n93), 
	.B2(U_cr_n547), 
	.B1(U_cr_n166), 
	.A2(U_cr_n546), 
	.A1(U_cr_n549));
   OAI22_X2 U_cr_U241 (.ZN(cr_reg_data_out[20]), 
	.B2(U_cr_n451), 
	.B1(U_cr_n467), 
	.A2(U_cr_n453), 
	.A1(U_cr_n462));
   OAI22_X2 U_cr_U240 (.ZN(cr_reg_data_out[25]), 
	.B2(U_cr_n453), 
	.B1(U_cr_n440), 
	.A2(U_cr_n451), 
	.A1(U_cr_n441));
   OAI22_X2 U_cr_U239 (.ZN(cr_reg_data_out[24]), 
	.B2(U_cr_n453), 
	.B1(U_cr_n439), 
	.A2(U_cr_n451), 
	.A1(U_cr_n486));
   OAI22_X2 U_cr_U238 (.ZN(cr_reg_data_out[28]), 
	.B2(U_cr_n453), 
	.B1(U_cr_n463), 
	.A2(U_cr_n451), 
	.A1(U_cr_n443));
   OAI22_X2 U_cr_U237 (.ZN(cr_reg_data_out[29]), 
	.B2(U_cr_n451), 
	.B1(U_cr_n444), 
	.A2(U_cr_n453), 
	.A1(U_cr_n468));
   OAI22_X2 U_cr_U236 (.ZN(cr_reg_data_out[19]), 
	.B2(U_cr_n451), 
	.B1(U_cr_n420), 
	.A2(U_cr_n453), 
	.A1(U_cr_n456));
   NAND4_X2 U_cr_U235 (.ZN(U_cr_n475), 
	.A4(U_cr_n386), 
	.A3(U_cr_n387), 
	.A2(U_cr_n388), 
	.A1(U_cr_n389));
   AOI22_X2 U_cr_U234 (.ZN(U_cr_n398), 
	.B2(U_cr_n476), 
	.B1(U_cr_n204), 
	.A2(U_cr_n475), 
	.A1(U_cr_n499));
   AOI22_X2 U_cr_U233 (.ZN(U_cr_n397), 
	.B2(U_cr_n478), 
	.B1(U_cr_n203), 
	.A2(U_cr_n477), 
	.A1(U_cr_n497));
   NAND2_X2 U_cr_U232 (.ZN(cr_reg_data_out[14]), 
	.A2(U_cr_n397), 
	.A1(U_cr_n398));
   OAI22_X2 U_cr_U231 (.ZN(cr_reg_data_out[21]), 
	.B2(U_cr_n451), 
	.B1(U_cr_n474), 
	.A2(U_cr_n453), 
	.A1(U_cr_n470));
   AOI22_X2 U_cr_U230 (.ZN(U_cr_n480), 
	.B2(U_cr_n475), 
	.B1(U_cr_n203), 
	.A2(U_cr_n476), 
	.A1(U_cr_n497));
   AOI22_X2 U_cr_U229 (.ZN(U_cr_n479), 
	.B2(U_cr_n477), 
	.B1(U_cr_n204), 
	.A2(U_cr_n478), 
	.A1(U_cr_n499));
   NAND2_X2 U_cr_U228 (.ZN(cr_reg_data_out[6]), 
	.A2(U_cr_n479), 
	.A1(U_cr_n480));
   OAI22_X2 U_cr_U227 (.ZN(cr_reg_data_out[30]), 
	.B2(U_cr_n451), 
	.B1(U_cr_n452), 
	.A2(U_cr_n453), 
	.A1(U_cr_n454));
   NOR2_X2 U_cr_U226 (.ZN(U_cr_n206), 
	.A2(FE_PHN1473_U_cr_n27), 
	.A1(FE_PHN2051_U_cr_n18));
   NAND2_X2 U_cr_U225 (.ZN(U_cr_n208), 
	.A2(U_cr_n206), 
	.A1(FE_PHN1150_U_cr_sctlr_14_));
   NAND2_X2 U_cr_U224 (.ZN(U_cr_n210), 
	.A2(U_cr_n209), 
	.A1(U_cr_sctlr_15_));
   AOI22_X2 U_cr_U223 (.ZN(U_cr_N573), 
	.B2(FE_PHN3107_U_cr_n44), 
	.B1(U_cr_n208), 
	.A2(U_cr_n209), 
	.A1(U_cr_sctlr_15_));
   NAND2_X2 U_cr_U222 (.ZN(U_cr_n282), 
	.A2(U_cr_stmg0r_1_), 
	.A1(FE_PHN1477_U_cr_stmg0r_0_));
   AOI21_X2 U_cr_U221 (.ZN(U_cr_N571), 
	.B2(FE_PHN1473_U_cr_n27), 
	.B1(FE_PHN2051_U_cr_n18), 
	.A(U_cr_n206));
   INV_X4 U_cr_U219 (.ZN(U_cr_n186), 
	.A(U_cr_n193));
   NOR2_X2 U_cr_U218 (.ZN(U_cr_n423), 
	.A2(U_cr_n308), 
	.A1(U_cr_n320));
   AOI22_X2 U_cr_U217 (.ZN(U_cr_n337), 
	.B2(cr_exn_mode_value[10]), 
	.B1(U_cr_n423), 
	.A2(U_cr_n559), 
	.A1(U_cr_n422));
   NOR2_X2 U_cr_U216 (.ZN(U_cr_n393), 
	.A2(U_cr_n378), 
	.A1(hiu_haddr[3]));
   AOI22_X2 U_cr_U215 (.ZN(U_cr_n374), 
	.B2(U_cr_n407), 
	.B1(FE_PHN1475_cr_s_data_width_early_0_), 
	.A2(U_cr_sctlr_13_), 
	.A1(U_cr_n422));
   AOI22_X2 U_cr_U214 (.ZN(U_cr_n402), 
	.B2(cr_t_ref[7]), 
	.B1(U_cr_n169), 
	.A2(FE_PHN955_s_read_pipe_1_), 
	.A1(U_cr_n422));
   NOR2_X2 U_cr_U213 (.ZN(U_cr_n319), 
	.A2(U_addrdec_n40), 
	.A1(FE_PHN4616_n27));
   NAND2_X1 U_cr_U212 (.ZN(U_cr_n202), 
	.A2(FE_PHN916_U_cr_cr_cs_2_), 
	.A1(U_cr_n187));
   NOR2_X2 U_cr_U211 (.ZN(U_cr_n273), 
	.A2(U_cr_n526), 
	.A1(U_cr_n396));
   INV_X4 U_cr_U210 (.ZN(U_cr_n169), 
	.A(U_cr_n170));
   AOI22_X2 U_cr_U209 (.ZN(U_cr_n361), 
	.B2(U_cr_n566), 
	.B1(U_cr_n424), 
	.A2(cr_ref_all_before_sr), 
	.A1(U_cr_n422));
   AOI22_X2 U_cr_U208 (.ZN(U_cr_n366), 
	.B2(cr_exn_mode_value[12]), 
	.B1(U_cr_n423), 
	.A2(U_cr_n571), 
	.A1(U_cr_n424));
   AOI22_X2 U_cr_U207 (.ZN(U_cr_n341), 
	.B2(cr_t_ras_min[0]), 
	.B1(U_cr_n430), 
	.A2(cr_do_power_down), 
	.A1(U_cr_n422));
   AOI22_X2 U_cr_U206 (.ZN(U_cr_n340), 
	.B2(cr_exn_mode_value[2]), 
	.B1(U_cr_n423), 
	.A2(U_cr_n568), 
	.A1(U_cr_n424));
   AOI22_X2 U_cr_U205 (.ZN(U_cr_n408), 
	.B2(cr_exn_mode_value[9]), 
	.B1(U_cr_n423), 
	.A2(U_cr_n561), 
	.A1(U_cr_n424));
   AOI22_X2 U_cr_U204 (.ZN(U_cr_n399), 
	.B2(cr_exn_mode_value[7]), 
	.B1(U_cr_n423), 
	.A2(U_cr_n563), 
	.A1(U_cr_n424));
   OAI222_X2 U_cr_U203 (.ZN(cr_reg_data_out[15]), 
	.C2(FE_PHN1103_U_cr_n455), 
	.C1(U_cr_n182), 
	.B2(U_cr_n438), 
	.B1(U_cr_n492), 
	.A2(U_cr_n437), 
	.A1(U_cr_n487));
   AOI22_X2 U_cr_U202 (.ZN(U_cr_n322), 
	.B2(cr_exn_mode_value[0]), 
	.B1(U_cr_n423), 
	.A2(U_cr_n570), 
	.A1(U_cr_n424));
   AOI22_X2 U_cr_U201 (.ZN(U_cr_n486), 
	.B2(U_cr_srefr[24]), 
	.B1(U_cr_n429), 
	.A2(cr_t_rc[2]), 
	.A1(U_cr_n430));
   AOI22_X2 U_cr_U200 (.ZN(U_cr_n425), 
	.B2(cr_exn_mode_value[1]), 
	.B1(U_cr_n423), 
	.A2(U_cr_n569), 
	.A1(U_cr_n424));
   NOR2_X2 U_cr_U199 (.ZN(U_cr_n232), 
	.A2(U_cr_n391), 
	.A1(U_cr_n544));
   AOI22_X2 U_cr_U198 (.ZN(U_cr_n386), 
	.B2(cr_exn_mode_value[6]), 
	.B1(U_cr_n423), 
	.A2(U_cr_n564), 
	.A1(U_cr_n424));
   NOR2_X1 U_cr_U197 (.ZN(U_cr_n201), 
	.A2(U_cr_n24), 
	.A1(U_cr_n192));
   NAND3_X1 U_cr_U196 (.ZN(U_cr_n197), 
	.A3(FE_PHN916_U_cr_cr_cs_2_), 
	.A2(FE_PHN837_U_cr_cr_cs_0_), 
	.A1(U_cr_n23));
   INV_X4 U_cr_U194 (.ZN(U_cr_n168), 
	.A(U_cr_n242));
   NOR2_X2 U_cr_U193 (.ZN(U_cr_n230), 
	.A2(U_cr_n391), 
	.A1(U_cr_n526));
   NOR2_X2 U_cr_U192 (.ZN(U_cr_n313), 
	.A2(U_cr_n334), 
	.A1(U_cr_n526));
   NOR2_X2 U_cr_U191 (.ZN(U_cr_n536), 
	.A2(U_cr_n543), 
	.A1(U_cr_n526));
   NOR2_X2 U_cr_U190 (.ZN(U_cr_n305), 
	.A2(U_cr_n358), 
	.A1(U_cr_n526));
   NOR2_X2 U_cr_U189 (.ZN(U_cr_n289), 
	.A2(U_cr_n170), 
	.A1(U_cr_n526));
   NOR2_X2 U_cr_U188 (.ZN(U_cr_n268), 
	.A2(U_cr_n25), 
	.A1(U_cr_n526));
   NAND2_X2 U_cr_U187 (.ZN(U_cr_n544), 
	.A2(U_cr_n216), 
	.A1(U_cr_n217));
   AOI22_X2 U_cr_U186 (.ZN(U_cr_n409), 
	.B2(n[26]), 
	.B1(U_cr_n407), 
	.A2(cr_mode_reg_update), 
	.A1(U_cr_n422));
   NOR2_X2 U_cr_U185 (.ZN(U_cr_n294), 
	.A2(U_cr_n170), 
	.A1(U_cr_n544));
   NOR2_X2 U_cr_U184 (.ZN(U_cr_n270), 
	.A2(U_cr_n25), 
	.A1(U_cr_n544));
   NOR2_X2 U_cr_U183 (.ZN(U_cr_n194), 
	.A2(FE_PHN916_U_cr_cr_cs_2_), 
	.A1(FE_PHN837_U_cr_cr_cs_0_));
   NOR2_X2 U_cr_U182 (.ZN(U_cr_n193), 
	.A2(U_cr_n23), 
	.A1(U_cr_n178));
   NAND2_X1 U_cr_U181 (.ZN(U_cr_n503), 
	.A2(U_cr_n16), 
	.A1(FE_PHN916_U_cr_cr_cs_2_));
   NAND2_X2 U_cr_U180 (.ZN(U_cr_n526), 
	.A2(U_cr_n213), 
	.A1(U_cr_n217));
   NAND2_X1 U_cr_U179 (.ZN(U_cr_n242), 
	.A2(big_endian), 
	.A1(FE_PHN4616_n27));
   NOR2_X4 U_cr_U178 (.ZN(U_cr_n422), 
	.A2(U_cr_n263), 
	.A1(U_cr_n320));
   AOI222_X1 U_cr_U177 (.ZN(U_cr_n290), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[5]), 
	.B2(hiu_wr_data[21]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[13]), 
	.A1(FE_OFN357_U_addrdec_n40));
   AOI222_X1 U_cr_U176 (.ZN(U_cr_n314), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[4]), 
	.B2(hiu_wr_data[20]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[12]), 
	.A1(U_addrdec_n40));
   AOI222_X1 U_cr_U175 (.ZN(U_cr_n541), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[3]), 
	.B2(hiu_wr_data[19]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[11]), 
	.A1(U_addrdec_n40));
   AOI222_X1 U_cr_U174 (.ZN(U_cr_n293), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[7]), 
	.B2(hiu_wr_data[23]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[15]), 
	.A1(U_addrdec_n40));
   AOI222_X1 U_cr_U173 (.ZN(U_cr_n291), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[6]), 
	.B2(hiu_wr_data[22]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[14]), 
	.A1(FE_OFN357_U_addrdec_n40));
   AOI222_X1 U_cr_U172 (.ZN(U_cr_n516), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[9]), 
	.B2(hiu_wr_data[25]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[1]), 
	.A1(FE_OFN357_U_addrdec_n40));
   AOI222_X1 U_cr_U171 (.ZN(U_cr_n514), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[8]), 
	.B2(hiu_wr_data[24]), 
	.B1(U_cr_n168), 
	.A2(hiu_wr_data[0]), 
	.A1(FE_OFN357_U_addrdec_n40));
   NOR2_X2 U_cr_U170 (.ZN(U_cr_n190), 
	.A2(FE_PHN1401_U_cr_cr_cs_1_), 
	.A1(FE_PHN916_U_cr_cr_cs_2_));
   MUX2_X1 U_cr_U168 (.Z(U_cr_n95), 
	.S(FE_PHN1400_U_cr_n197), 
	.B(FE_PHN2432_n27), 
	.A(FE_PHN1475_cr_s_data_width_early_0_));
   NAND2_X2 U_cr_U167 (.ZN(U_cr_n200), 
	.A2(U_cr_n24), 
	.A1(U_cr_n191));
   INV_X1 U_cr_U166 (.ZN(U_cr_n192), 
	.A(U_cr_n191));
   OAI21_X1 U_cr_U165 (.ZN(U_cr_n207), 
	.B2(U_cr_n206), 
	.B1(FE_PHN1150_U_cr_sctlr_14_), 
	.A(U_cr_n208));
   INV_X2 U_cr_U164 (.ZN(U_cr_n209), 
	.A(U_cr_n208));
   INV_X2 U_cr_U162 (.ZN(U_cr_N572), 
	.A(U_cr_n207));
   NAND2_X1 U_cr_U161 (.ZN(U_cr_n179), 
	.A2(U_cr_n319), 
	.A1(U_cr_n193));
   NAND2_X1 U_cr_U160 (.ZN(U_cr_n360), 
	.A2(hiu_addr[6]), 
	.A1(hiu_haddr[2]));
   INV_X2 U_cr_U159 (.ZN(U_cr_n283), 
	.A(hiu_haddr[3]));
   NOR2_X1 U_cr_U158 (.ZN(U_cr_n284), 
	.A2(hiu_addr[7]), 
	.A1(hiu_addr[5]));
   NOR2_X1 U_cr_U157 (.ZN(U_cr_n300), 
	.A2(hiu_addr[4]), 
	.A1(hiu_addr[6]));
   INV_X2 U_cr_U156 (.ZN(U_cr_n320), 
	.A(hiu_haddr[2]));
   INV_X1 U_cr_U155 (.ZN(U_cr_n316), 
	.A(hiu_addr[6]));
   NAND3_X1 U_cr_U154 (.ZN(U_cr_n359), 
	.A3(hiu_addr[4]), 
	.A2(hiu_addr[7]), 
	.A1(hiu_addr[5]));
   NAND4_X1 U_cr_U153 (.ZN(U_cr_n308), 
	.A4(U_cr_n300), 
	.A3(hiu_addr[7]), 
	.A2(hiu_addr[5]), 
	.A1(hiu_haddr[3]));
   NOR2_X1 U_cr_U152 (.ZN(U_cr_n383), 
	.A2(U_cr_n21), 
	.A1(U_cr_n416));
   NOR2_X1 U_cr_U151 (.ZN(U_cr_n351), 
	.A2(U_cr_n36), 
	.A1(U_cr_n416));
   NAND3_X1 U_cr_U150 (.ZN(U_cr_n196), 
	.A3(FE_PHN837_U_cr_cr_cs_0_), 
	.A2(U_cr_n190), 
	.A1(U_cr_n550));
   AOI22_X1 U_cr_U149 (.ZN(U_cr_n353), 
	.B2(gpo[3]), 
	.B1(U_cr_n429), 
	.A2(U_cr_s_sda_d1), 
	.A1(U_cr_n407));
   INV_X2 U_cr_U148 (.ZN(U_cr_n377), 
	.A(U_cr_n412));
   AOI22_X1 U_cr_U147 (.ZN(U_cr_n401), 
	.B2(FE_PHN1855_cr_block_size1_7_), 
	.B1(U_cr_n525), 
	.A2(FE_PHN3054_cr_row_addr_width_2_), 
	.A1(U_cr_n407));
   OAI22_X1 U_cr_U146 (.ZN(U_cr_n222), 
	.B2(U_cr_n503), 
	.B1(FE_PHN1401_U_cr_cr_cs_1_), 
	.A2(U_cr_n200), 
	.A1(U_cr_n318));
   AOI21_X1 U_cr_U145 (.ZN(U_cr_n505), 
	.B2(U_cr_n504), 
	.B1(hiu_reg_req), 
	.A(FE_PHN837_U_cr_cr_cs_0_));
   AOI22_X1 U_cr_U144 (.ZN(U_cr_n380), 
	.B2(cr_t_init[5]), 
	.B1(U_cr_n171), 
	.A2(U_cr_n565), 
	.A1(U_cr_n424));
   AOI22_X1 U_cr_U143 (.ZN(U_cr_n388), 
	.B2(cr_t_init[6]), 
	.B1(U_cr_n171), 
	.A2(cr_t_rcd[0]), 
	.A1(U_cr_n430));
   OAI21_X2 U_cr_U142 (.ZN(U_cr_n217), 
	.B2(U_cr_n317), 
	.B1(U_cr_n200), 
	.A(U_cr_n17));
   NAND4_X1 U_cr_U141 (.ZN(U_cr_n96), 
	.A4(U_cr_n195), 
	.A3(U_cr_n198), 
	.A2(U_cr_n205), 
	.A1(U_cr_n196));
   AOI22_X1 U_cr_U140 (.ZN(U_cr_n400), 
	.B2(cr_t_init[7]), 
	.B1(U_cr_n171), 
	.A2(cr_t_rcd[1]), 
	.A1(U_cr_n430));
   OAI21_X1 U_cr_U139 (.ZN(U_cr_n98), 
	.B2(U_cr_n199), 
	.B1(U_cr_n505), 
	.A(U_cr_n198));
   INV_X2 U_cr_U138 (.ZN(U_cr_n403), 
	.A(U_cr_n484));
   INV_X1 U_cr_U137 (.ZN(U_cr_n189), 
	.A(U_cr_n188));
   AOI22_X1 U_cr_U136 (.ZN(U_cr_n404), 
	.B2(cr_t_init[15]), 
	.B1(U_cr_n171), 
	.A2(cr_t_rcar[1]), 
	.A1(U_cr_n430));
   AOI22_X1 U_cr_U135 (.ZN(U_cr_n394), 
	.B2(cr_t_init[14]), 
	.B1(U_cr_n171), 
	.A2(cr_t_rcar[0]), 
	.A1(U_cr_n430));
   AND2_X2 U_cr_U134 (.ZN(U_cr_n238), 
	.A2(U_cr_n17), 
	.A1(U_cr_n222));
   AOI21_X1 U_cr_U133 (.ZN(U_cr_n426), 
	.B2(U_cr_n422), 
	.B1(cr_do_self_ref_rp), 
	.A(U_cr_n421));
   AOI22_X1 U_cr_U132 (.ZN(U_cr_n348), 
	.B2(cr_t_init[3]), 
	.B1(U_cr_n171), 
	.A2(U_cr_n567), 
	.A1(U_cr_n424));
   NOR2_X1 U_cr_U131 (.ZN(U_cr_n335), 
	.A2(U_cr_n37), 
	.A1(U_cr_n334));
   AOI22_X1 U_cr_U130 (.ZN(U_cr_n375), 
	.B2(cr_t_init[13]), 
	.B1(U_cr_n171), 
	.A2(cr_t_wr[1]), 
	.A1(U_cr_n430));
   NAND2_X1 U_cr_U129 (.ZN(U_cr_n175), 
	.A2(U_addrdec_n40), 
	.A1(U_cr_n317));
   AOI21_X1 U_cr_U128 (.ZN(U_cr_n332), 
	.B2(U_cr_n430), 
	.B1(cr_t_xsr[0]), 
	.A(U_cr_n377));
   AOI22_X1 U_cr_U127 (.ZN(U_cr_n363), 
	.B2(cr_t_init[4]), 
	.B1(U_cr_n171), 
	.A2(cr_t_ras_min[2]), 
	.A1(U_cr_n430));
   AOI22_X1 U_cr_U126 (.ZN(U_cr_n428), 
	.B2(U_cr_n557), 
	.B1(U_cr_n525), 
	.A2(cr_t_ref[1]), 
	.A1(U_cr_n169));
   AND2_X2 U_cr_U125 (.ZN(U_cr_n344), 
	.A2(U_cr_stmg0r_26), 
	.A1(U_cr_n430));
   AOI22_X1 U_cr_U124 (.ZN(U_cr_n427), 
	.B2(cr_t_init[1]), 
	.B1(U_cr_n171), 
	.A2(U_cr_stmg0r_1_), 
	.A1(U_cr_n430));
   AOI22_X1 U_cr_U123 (.ZN(U_cr_n373), 
	.B2(U_cr_srefr[29]), 
	.B1(U_cr_n169), 
	.A2(cr_t_xsr[6]), 
	.A1(U_cr_n430));
   AOI22_X1 U_cr_U122 (.ZN(U_cr_n324), 
	.B2(cr_t_init[0]), 
	.B1(U_cr_n171), 
	.A2(FE_PHN1477_U_cr_stmg0r_0_), 
	.A1(U_cr_n430));
   AOI22_X1 U_cr_U121 (.ZN(U_cr_n410), 
	.B2(cr_t_init[9]), 
	.B1(U_cr_n171), 
	.A2(cr_t_rp[0]), 
	.A1(U_cr_n430));
   AOI21_X1 U_cr_U120 (.ZN(U_cr_n390), 
	.B2(U_cr_n169), 
	.B1(gpo[6]), 
	.A(U_cr_n392));
   NAND2_X1 U_cr_U119 (.ZN(U_cr_n237), 
	.A2(U_cr_n236), 
	.A1(U_cr_n430));
   AOI22_X1 U_cr_U118 (.ZN(U_cr_n389), 
	.B2(FE_PHN3126_cr_block_size1_6_), 
	.B1(U_cr_n525), 
	.A2(cr_t_ref[6]), 
	.A1(U_cr_n169));
   AOI22_X1 U_cr_U117 (.ZN(U_cr_n411), 
	.B2(U_cr_n552), 
	.B1(U_cr_n525), 
	.A2(cr_t_ref[9]), 
	.A1(U_cr_n169));
   AOI21_X1 U_cr_U116 (.ZN(U_cr_n327), 
	.B2(U_cr_n430), 
	.B1(cr_t_rcar[2]), 
	.A(U_cr_n377));
   OAI211_X1 U_cr_U115 (.ZN(U_cr_n414), 
	.C2(U_cr_n170), 
	.C1(U_cr_n29), 
	.B(U_cr_n412), 
	.A(U_cr_n413));
   AOI22_X1 U_cr_U114 (.ZN(U_cr_n325), 
	.B2(FE_PHN1088_U_cr_n558), 
	.B1(U_cr_n525), 
	.A2(cr_t_ref[0]), 
	.A1(U_cr_n169));
   AOI22_X1 U_cr_U113 (.ZN(U_cr_n381), 
	.B2(cr_block_size1[5]), 
	.B1(U_cr_n525), 
	.A2(cr_t_ref[5]), 
	.A1(U_cr_n169));
   OAI21_X1 U_cr_U112 (.ZN(cr_push_n), 
	.B2(FE_PHN1401_U_cr_cr_cs_1_), 
	.B1(U_cr_n189), 
	.A(U_cr_n194));
   AOI22_X1 U_cr_U111 (.ZN(U_cr_n349), 
	.B2(U_cr_n555), 
	.B1(U_cr_n525), 
	.A2(cr_t_ref[3]), 
	.A1(U_cr_n169));
   AOI22_X1 U_cr_U110 (.ZN(U_cr_n357), 
	.B2(U_cr_srefr[28]), 
	.B1(U_cr_n169), 
	.A2(cr_t_xsr[5]), 
	.A1(U_cr_n430));
   OAI211_X1 U_cr_U109 (.ZN(U_cr_n333), 
	.C2(U_cr_n30), 
	.C1(U_cr_n416), 
	.B(U_cr_n331), 
	.A(U_cr_n332));
   OAI211_X1 U_cr_U108 (.ZN(U_cr_n328), 
	.C2(U_cr_n28), 
	.C1(U_cr_n416), 
	.B(U_cr_n326), 
	.A(U_cr_n327));
   OAI211_X1 U_cr_U107 (.ZN(U_cr_n356), 
	.C2(U_cr_n391), 
	.C1(U_cr_n33), 
	.B(U_cr_n412), 
	.A(U_cr_n355));
   INV_X2 U_cr_U106 (.ZN(U_cr_n420), 
	.A(U_cr_n459));
   INV_X2 U_cr_U105 (.ZN(U_cr_n440), 
	.A(U_cr_n498));
   INV_X2 U_cr_U104 (.ZN(U_cr_n443), 
	.A(U_cr_n465));
   INV_X2 U_cr_U103 (.ZN(U_cr_n444), 
	.A(U_cr_n472));
   INV_X2 U_cr_U102 (.ZN(U_cr_n418), 
	.A(U_cr_n495));
   INV_X2 U_cr_U101 (.ZN(U_cr_n435), 
	.A(U_cr_n478));
   INV_X2 U_cr_U100 (.ZN(U_cr_n436), 
	.A(U_cr_n476));
   INV_X2 U_cr_U99 (.ZN(U_cr_n441), 
	.A(U_cr_n496));
   INV_X2 U_cr_U98 (.ZN(U_cr_n439), 
	.A(U_cr_n490));
   INV_X2 U_cr_U97 (.ZN(U_cr_n419), 
	.A(U_cr_n448));
   NAND2_X1 U_cr_U96 (.ZN(U_cr_n219), 
	.A2(U_cr_n221), 
	.A1(U_cr_n291));
   INV_X2 U_cr_U95 (.ZN(U_cr_n454), 
	.A(U_cr_n475));
   INV_X1 U_cr_U94 (.ZN(U_cr_n181), 
	.A(U_cr_n182));
   NAND2_X1 U_cr_U93 (.ZN(U_cr_n218), 
	.A2(FE_PHN1475_cr_s_data_width_early_0_), 
	.A1(U_cr_n219));
   NOR2_X1 U_cr_U92 (.ZN(cr_reg_data_out[31]), 
	.A2(U_cr_n185), 
	.A1(FE_PHN1103_U_cr_n455));
   INV_X2 U_cr_U91 (.ZN(U_cr_n477), 
	.A(U_cr_n452));
   INV_X2 U_cr_U90 (.ZN(U_cr_n417), 
	.A(U_cr_n494));
   OAI22_X1 U_cr_U89 (.ZN(U_cr_n286), 
	.B2(U_cr_n289), 
	.B1(cr_t_ref[1]), 
	.A2(U_cr_n534), 
	.A1(U_cr_n288));
   NAND2_X1 U_cr_U88 (.ZN(U_cr_n249), 
	.A2(U_cr_n259), 
	.A1(hiu_wr_data[3]));
   OAI22_X1 U_cr_U87 (.ZN(U_cr_n309), 
	.B2(U_cr_n313), 
	.B1(U_cr_n570), 
	.A2(U_cr_n537), 
	.A1(U_cr_n312));
   NAND2_X1 U_cr_U86 (.ZN(U_cr_n247), 
	.A2(U_cr_n259), 
	.A1(hiu_wr_data[2]));
   OAI22_X1 U_cr_U85 (.ZN(U_cr_n228), 
	.B2(U_cr_n230), 
	.B1(cr_t_ras_min[0]), 
	.A2(U_cr_n532), 
	.A1(U_cr_n229));
   OAI22_X1 U_cr_U84 (.ZN(U_cr_n310), 
	.B2(U_cr_n313), 
	.B1(U_cr_n569), 
	.A2(U_cr_n534), 
	.A1(U_cr_n312));
   NAND2_X1 U_cr_U83 (.ZN(U_cr_n245), 
	.A2(U_cr_n259), 
	.A1(hiu_wr_data[1]));
   OAI22_X1 U_cr_U82 (.ZN(U_cr_n266), 
	.B2(U_cr_n268), 
	.B1(cr_t_init[2]), 
	.A2(U_cr_n532), 
	.A1(U_cr_n267));
   NAND2_X1 U_cr_U81 (.ZN(U_cr_n243), 
	.A2(U_cr_n259), 
	.A1(hiu_wr_data[0]));
   OAI22_X1 U_cr_U80 (.ZN(U_cr_n265), 
	.B2(U_cr_n268), 
	.B1(cr_t_init[1]), 
	.A2(U_cr_n534), 
	.A1(U_cr_n267));
   OAI22_X1 U_cr_U79 (.ZN(U_cr_n264), 
	.B2(U_cr_n268), 
	.B1(FE_PHN3041_cr_t_init_0_), 
	.A2(U_cr_n537), 
	.A1(U_cr_n267));
   OAI22_X1 U_cr_U78 (.ZN(U_cr_n311), 
	.B2(U_cr_n313), 
	.B1(U_cr_n568), 
	.A2(U_cr_n532), 
	.A1(U_cr_n312));
   INV_X2 U_cr_U77 (.ZN(U_cr_n184), 
	.A(FE_PHN948_U_cr_n442));
   OAI22_X1 U_cr_U76 (.ZN(U_cr_n533), 
	.B2(U_cr_n536), 
	.B1(U_cr_n556), 
	.A2(U_cr_n532), 
	.A1(U_cr_n538));
   OAI22_X1 U_cr_U75 (.ZN(U_cr_n535), 
	.B2(U_cr_n536), 
	.B1(U_cr_n557), 
	.A2(U_cr_n534), 
	.A1(U_cr_n538));
   OAI22_X1 U_cr_U74 (.ZN(U_cr_n539), 
	.B2(U_cr_n536), 
	.B1(FE_PHN1088_U_cr_n558), 
	.A2(U_cr_n537), 
	.A1(U_cr_n538));
   AND2_X2 U_cr_U73 (.ZN(cr_reg_data_out[23]), 
	.A2(FE_PHN1163_U_cr_n482), 
	.A1(U_cr_n13));
   OAI21_X1 U_cr_U72 (.ZN(U_cr_N308), 
	.B2(U_cr_n219), 
	.B1(U_cr_n290), 
	.A(U_cr_n218));
   OAI22_X1 U_cr_U71 (.ZN(U_cr_n301), 
	.B2(U_cr_n305), 
	.B1(cr_exn_mode_value[0]), 
	.A2(U_cr_n537), 
	.A1(U_cr_n304));
   OAI22_X1 U_cr_U70 (.ZN(U_cr_n302), 
	.B2(U_cr_n305), 
	.B1(cr_exn_mode_value[1]), 
	.A2(U_cr_n534), 
	.A1(U_cr_n304));
   OAI22_X1 U_cr_U69 (.ZN(U_cr_n303), 
	.B2(U_cr_n305), 
	.B1(cr_exn_mode_value[2]), 
	.A2(U_cr_n532), 
	.A1(U_cr_n304));
   OAI22_X1 U_cr_U68 (.ZN(U_cr_n287), 
	.B2(U_cr_n289), 
	.B1(cr_t_ref[2]), 
	.A2(U_cr_n532), 
	.A1(U_cr_n288));
   OAI22_X1 U_cr_U67 (.ZN(U_cr_n285), 
	.B2(U_cr_n289), 
	.B1(cr_t_ref[0]), 
	.A2(U_cr_n537), 
	.A1(U_cr_n288));
   NAND2_X1 U_cr_U66 (.ZN(U_cr_n260), 
	.A2(U_cr_n259), 
	.A1(hiu_wr_data[7]));
   NAND2_X1 U_cr_U65 (.ZN(U_cr_n251), 
	.A2(U_cr_n259), 
	.A1(hiu_wr_data[4]));
   NAND2_X1 U_cr_U64 (.ZN(U_cr_n253), 
	.A2(U_cr_n259), 
	.A1(hiu_wr_data[5]));
   NAND2_X1 U_cr_U63 (.ZN(U_cr_n255), 
	.A2(U_cr_n259), 
	.A1(hiu_wr_data[6]));
   OAI22_X1 U_cr_U62 (.ZN(U_cr_n271), 
	.B2(U_cr_n273), 
	.B1(cr_do_power_down), 
	.A2(U_cr_n532), 
	.A1(U_cr_n272));
   INV_X2 U_cr_U61 (.ZN(U_cr_N464), 
	.A(U_cr_n264));
   OAI211_X1 U_cr_U60 (.ZN(U_cr_N417), 
	.C2(U_cr_n262), 
	.C1(FE_OFN0_U_cr_n314), 
	.B(U_cr_n251), 
	.A(U_cr_n252));
   NOR2_X1 U_cr_U59 (.ZN(cr_reg_data_out[27]), 
	.A2(U_cr_n185), 
	.A1(U_cr_n184));
   INV_X2 U_cr_U58 (.ZN(U_cr_N552), 
	.A(U_cr_n271));
   INV_X2 U_cr_U57 (.ZN(U_cr_N734), 
	.A(U_cr_n310));
   OAI211_X1 U_cr_U56 (.ZN(U_cr_N416), 
	.C2(U_cr_n262), 
	.C1(FE_OFN1_U_cr_n541), 
	.B(U_cr_n249), 
	.A(U_cr_n250));
   INV_X2 U_cr_U55 (.ZN(U_cr_n87), 
	.A(U_cr_n539));
   OAI211_X1 U_cr_U54 (.ZN(U_cr_N418), 
	.C2(U_cr_n262), 
	.C1(U_cr_n290), 
	.B(U_cr_n253), 
	.A(U_cr_n254));
   INV_X2 U_cr_U53 (.ZN(U_cr_N465), 
	.A(U_cr_n265));
   INV_X2 U_cr_U52 (.ZN(U_cr_N634), 
	.A(U_cr_n287));
   INV_X2 U_cr_U51 (.ZN(U_cr_N690), 
	.A(U_cr_n303));
   OAI211_X1 U_cr_U50 (.ZN(U_cr_N419), 
	.C2(U_cr_n262), 
	.C1(U_cr_n291), 
	.B(U_cr_n255), 
	.A(U_cr_n256));
   INV_X2 U_cr_U49 (.ZN(U_cr_N391), 
	.A(U_cr_n228));
   INV_X2 U_cr_U48 (.ZN(U_cr_N466), 
	.A(U_cr_n266));
   INV_X2 U_cr_U47 (.ZN(U_cr_N688), 
	.A(U_cr_n301));
   OAI211_X1 U_cr_U46 (.ZN(U_cr_N420), 
	.C2(U_cr_n262), 
	.C1(U_cr_n293), 
	.B(U_cr_n260), 
	.A(U_cr_n261));
   OAI211_X1 U_cr_U45 (.ZN(U_cr_N413), 
	.C2(U_cr_n262), 
	.C1(U_cr_n548), 
	.B(U_cr_n243), 
	.A(U_cr_n244));
   INV_X2 U_cr_U44 (.ZN(U_cr_n86), 
	.A(U_cr_n535));
   INV_X2 U_cr_U43 (.ZN(U_cr_N733), 
	.A(U_cr_n309));
   INV_X2 U_cr_U42 (.ZN(U_cr_N735), 
	.A(U_cr_n311));
   INV_X2 U_cr_U41 (.ZN(U_cr_N689), 
	.A(U_cr_n302));
   INV_X2 U_cr_U40 (.ZN(U_cr_n85), 
	.A(U_cr_n533));
   OAI21_X1 U_cr_U39 (.ZN(cr_reg_data_out[11]), 
	.B2(U_cr_n492), 
	.B1(U_cr_n456), 
	.A(U_cr_n354));
   OAI21_X1 U_cr_U38 (.ZN(cr_reg_data_out[7]), 
	.B2(U_cr_n487), 
	.B1(U_cr_n484), 
	.A(U_cr_n483));
   OAI21_X1 U_cr_U37 (.ZN(cr_reg_data_out[8]), 
	.B2(U_cr_n492), 
	.B1(U_cr_n493), 
	.A(U_cr_n491));
   OAI21_X1 U_cr_U36 (.ZN(cr_reg_data_out[10]), 
	.B2(U_cr_n487), 
	.B1(U_cr_n450), 
	.A(U_cr_n346));
   NOR2_X1 U_cr_U35 (.ZN(U_cr_n191), 
	.A2(U_cr_n16), 
	.A1(U_cr_n23));
   AOI22_X1 U_cr_U34 (.ZN(U_cr_N576), 
	.B2(FE_PHN2455_U_cr_n20), 
	.B1(FE_PHN3106_U_cr_n43), 
	.A2(U_cr_stmg0r_1_), 
	.A1(FE_PHN1477_U_cr_stmg0r_0_));
   INV_X4 U_cr_U33 (.ZN(U_cr_n178), 
	.A(U_cr_n194));
   NOR2_X1 U_cr_U32 (.ZN(U_cr_n198), 
	.A2(U_cr_n193), 
	.A1(U_cr_n201));
   NAND2_X1 U_cr_U31 (.ZN(U_cr_n502), 
	.A2(hiu_rw), 
	.A1(FE_PHN1401_U_cr_cr_cs_1_));
   NOR2_X1 U_cr_U30 (.ZN(U_cr_n211), 
	.A2(FE_OFN217_hiu_burst_size_2_), 
	.A1(FE_OFN214_hiu_burst_size_4_));
   NAND2_X1 U_cr_U29 (.ZN(U_cr_n188), 
	.A2(hiu_rw), 
	.A1(hiu_reg_req));
   OR2_X2 U_cr_U28 (.ZN(U_cr_n240), 
	.A2(U_cr_n222), 
	.A1(n27));
   AOI22_X1 U_cr_U27 (.ZN(U_cr_n413), 
	.B2(cr_num_init_ref[1]), 
	.B1(U_cr_n171), 
	.A2(cr_t_rcar[3]), 
	.A1(U_cr_n430));
   AOI22_X1 U_cr_U26 (.ZN(U_cr_n355), 
	.B2(gpo[4]), 
	.B1(U_cr_n169), 
	.A2(s_sda_oe_n), 
	.A1(U_cr_n407));
   AOI22_X1 U_cr_U25 (.ZN(U_cr_n432), 
	.B2(U_cr_srefr[25]), 
	.B1(U_cr_n169), 
	.A2(cr_t_rc[3]), 
	.A1(U_cr_n430));
   OAI21_X1 U_cr_U24 (.ZN(U_cr_n476), 
	.B2(FE_OFN23_U_cr_n64), 
	.B1(U_cr_n391), 
	.A(U_cr_n390));
   OAI21_X1 U_cr_U23 (.ZN(cr_reg_data_out[13]), 
	.B2(U_cr_n487), 
	.B1(U_cr_n474), 
	.A(U_cr_n385));
   OAI21_X1 U_cr_U22 (.ZN(cr_reg_data_out[3]), 
	.B2(U_cr_n492), 
	.B1(U_cr_n461), 
	.A(U_cr_n460));
   INV_X1 U_cr_U21 (.ZN(U_cr_n185), 
	.A(U_cr_n13));
   AOI21_X1 U_cr_U20 (.ZN(U_cr_n13), 
	.B2(U_cr_n17), 
	.B1(U_cr_n193), 
	.A(U_cr_n177));
   AOI211_X1 U_cr_U19 (.ZN(U_cr_n452), 
	.C2(cr_t_xsr[7]), 
	.C1(U_cr_n430), 
	.B(U_cr_n392), 
	.A(U_cr_n12));
   AND2_X1 U_cr_U18 (.ZN(U_cr_n12), 
	.A2(U_cr_srefr[30]), 
	.A1(U_cr_n169));
   NAND3_X1 U_cr_U17 (.ZN(U_cr_n99), 
	.A3(U_cr_n11), 
	.A2(U_cr_n10), 
	.A1(U_cr_n202));
   NAND4_X1 U_cr_U16 (.ZN(U_cr_n11), 
	.A4(hiu_reg_req), 
	.A3(U_cr_n17), 
	.A2(U_cr_n16), 
	.A1(U_cr_n23));
   AOI21_X1 U_cr_U15 (.ZN(U_cr_n10), 
	.B2(U_cr_n9), 
	.B1(U_cr_n550), 
	.A(U_cr_n201));
   INV_X1 U_cr_U14 (.ZN(U_cr_n9), 
	.A(U_cr_n200));
   AOI21_X1 U_cr_U13 (.ZN(U_cr_n456), 
	.B2(FE_OFN348_U_cr_n169), 
	.B1(cr_t_ref[11]), 
	.A(U_cr_n8));
   NAND4_X1 U_cr_U12 (.ZN(U_cr_n8), 
	.A4(U_cr_n378), 
	.A3(U_cr_n7), 
	.A2(U_cr_n6), 
	.A1(U_cr_n5));
   AOI22_X1 U_cr_U11 (.ZN(U_cr_n7), 
	.B2(U_cr_n422), 
	.B1(U_cr_sctlr_default_11), 
	.A2(U_cr_n407), 
	.A1(n[24]));
   AOI22_X1 U_cr_U10 (.ZN(U_cr_n6), 
	.B2(cr_t_rp[2]), 
	.B1(U_cr_n430), 
	.A2(cr_t_init[11]), 
	.A1(U_cr_n171));
   AOI22_X1 U_cr_U9 (.ZN(U_cr_n5), 
	.B2(U_cr_n423), 
	.B1(cr_exn_mode_value[11]), 
	.A2(U_cr_n560), 
	.A1(U_cr_n424));
   AOI222_X1 U_cr_U8 (.ZN(U_cr_n518), 
	.C2(U_cr_n319), 
	.C1(hiu_wr_data[10]), 
	.B2(U_cr_n168), 
	.B1(FE_OFN226_hiu_data_26_), 
	.A2(hiu_wr_data[2]), 
	.A1(FE_OFN357_U_addrdec_n40));
   AOI211_X1 U_cr_U7 (.ZN(U_cr_n493), 
	.C2(cr_t_ref[8]), 
	.C1(U_cr_n169), 
	.B(U_cr_n4), 
	.A(U_cr_n392));
   NAND3_X1 U_cr_U6 (.ZN(U_cr_n4), 
	.A3(U_cr_n3), 
	.A2(U_cr_n2), 
	.A1(U_cr_n1));
   AOI222_X1 U_cr_U5 (.ZN(U_cr_n3), 
	.C2(FE_PHN1064_cr_row_addr_width_3_), 
	.C1(U_cr_n407), 
	.B2(cr_exn_mode_value[8]), 
	.B1(U_cr_n423), 
	.A2(cr_t_rcd[2]), 
	.A1(U_cr_n430));
   AOI22_X1 U_cr_U4 (.ZN(U_cr_n2), 
	.B2(U_cr_n553), 
	.B1(U_cr_n525), 
	.A2(s_read_pipe[2]), 
	.A1(U_cr_n422));
   AOI22_X1 U_cr_U3 (.ZN(U_cr_n1), 
	.B2(U_cr_n562), 
	.B1(U_cr_n424), 
	.A2(cr_t_init[8]), 
	.A1(U_cr_n171));
   DFFR_X2 U_cr_smskr0_reg_8_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n154), 
	.Q(U_cr_n553), 
	.D(FE_PHN1522_U_cr_n94), 
	.CK(HCLK__L5_N35));
   DFFR_X2 U_cr_smskr0_reg_10_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n153), 
	.Q(U_cr_n551), 
	.D(FE_PHN1690_U_cr_n92), 
	.CK(HCLK__L5_N35));
   DFFR_X2 U_cr_cr_cs_reg_2_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_cr_n24), 
	.Q(U_cr_cr_cs_2_), 
	.D(FE_PHN800_U_cr_n96), 
	.CK(HCLK__L5_N17));
   DFFR_X2 U_cr_cr_cs_reg_0_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_cr_n16), 
	.Q(U_cr_cr_cs_0_), 
	.D(FE_PHN840_U_cr_n99), 
	.CK(HCLK__L5_N17));
   DFFR_X2 U_cr_cr_cs_reg_1_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_cr_n23), 
	.Q(U_cr_cr_cs_1_), 
	.D(FE_PHN926_U_cr_n98), 
	.CK(HCLK__L5_N17));
   DFFR_X2 U_cr_open_banks_o_reg_4_ (.RN(FE_OFN39_HRESETn), 
	.Q(cr_num_open_banks[4]), 
	.D(FE_PHN1661_U_cr_N574), 
	.CK(HCLK__L5_N11));
   DFFR_X2 U_cr_sctlr_reg_11_ (.RN(FE_OFN59_HRESETn), 
	.Q(U_cr_sctlr_default_11), 
	.D(FE_PHN3046_ctl_sd_in_sf_mode), 
	.CK(HCLK__L5_N11));
   DFFR_X2 U_cr_open_banks_o_reg_3_ (.RN(FE_OFN39_HRESETn), 
	.QN(n92), 
	.Q(cr_num_open_banks[3]), 
	.D(FE_PHN1256_U_cr_N573), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_cr_cas_latency_o_reg_2_ (.RN(FE_OFN188_HRESETn), 
	.QN(n91), 
	.Q(s_cas_latency[2]), 
	.D(FE_PHN1656_U_cr_N577), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_cr_open_banks_o_reg_2_ (.RN(FE_OFN39_HRESETn), 
	.Q(cr_num_open_banks[2]), 
	.D(U_cr_N572), 
	.CK(HCLK__L5_N11));
   DFFR_X2 U_cr_s_sda_d1_reg (.RN(FE_OFN51_HRESETn), 
	.Q(U_cr_s_sda_d1), 
	.D(FE_PHN2905_U_cr_s_sda_d), 
	.CK(hclk));
   DFFR_X2 U_cr_cas_latency_o_reg_0_ (.RN(FE_OFN188_HRESETn), 
	.QN(n90), 
	.Q(s_cas_latency[0]), 
	.D(FE_PHN2455_U_cr_n20), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_cr_syflash_opcode_reg_10_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n37), 
	.D(FE_PHN1378_U_cr_n90), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_srefr_reg_1_ (.SN(FE_OFN151_HRESETn), 
	.QN(cr_t_ref[1]), 
	.D(FE_PHN1628_U_cr_n286), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_srefr_reg_0_ (.SN(FE_OFN151_HRESETn), 
	.QN(cr_t_ref[0]), 
	.Q(n87), 
	.D(FE_PHN1918_U_cr_n285), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_srefr_reg_16_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n47), 
	.Q(gpo[0]), 
	.D(FE_PHN1376_U_cr_N648), 
	.CK(hclk));
   DFFR_X1 U_cr_srefr_reg_17_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n29), 
	.Q(gpo[1]), 
	.D(FE_PHN1375_U_cr_N649), 
	.CK(hclk));
   DFFR_X1 U_cr_srefr_reg_18_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_cr_n48), 
	.Q(gpo[2]), 
	.D(FE_PHN1083_U_cr_N650), 
	.CK(hclk));
   DFFR_X1 U_cr_srefr_reg_19_ (.RN(FE_OFN51_HRESETn), 
	.QN(U_cr_n49), 
	.Q(gpo[3]), 
	.D(FE_PHN1017_U_cr_N651), 
	.CK(hclk));
   DFFR_X1 U_cr_srefr_reg_20_ (.RN(FE_OFN51_HRESETn), 
	.QN(U_cr_n50), 
	.Q(gpo[4]), 
	.D(FE_PHN1044_U_cr_N652), 
	.CK(hclk));
   DFFR_X1 U_cr_srefr_reg_21_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_cr_n19), 
	.Q(gpo[5]), 
	.D(FE_PHN1119_U_cr_N653), 
	.CK(hclk));
   DFFR_X1 U_cr_srefr_reg_22_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_cr_n46), 
	.Q(gpo[6]), 
	.D(FE_PHN1118_U_cr_N654), 
	.CK(hclk));
   DFFR_X1 U_cr_srefr_reg_23_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_cr_n51), 
	.Q(gpo[7]), 
	.D(FE_PHN1243_U_cr_N655), 
	.CK(hclk));
   DFFR_X1 U_cr_sctlr_reg_18_ (.RN(FE_OFN63_HRESETn), 
	.Q(cr_exn_mode_reg_update), 
	.D(FE_PHN1014_U_cr_N567), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sctlr_reg_17_ (.RN(FE_OFN63_HRESETn), 
	.Q(cr_s_ready_valid), 
	.D(FE_PHN2915_U_cr_N566), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sctlr_reg_16_ (.RN(FE_OFN63_HRESETn), 
	.Q(U_cr_sctlr_16_), 
	.D(FE_PHN759_U_cr_N565), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sctlr_reg_19_ (.RN(FE_OFN51_HRESETn), 
	.Q(U_cr_n572), 
	.D(FE_PHN1013_U_cr_n73), 
	.CK(hclk));
   DFFS_X2 U_cr_stmg1r_reg_16_ (.SN(FE_OFN63_HRESETn), 
	.QN(U_cr_n115), 
	.Q(cr_num_init_ref[0]), 
	.D(FE_PHN1519_U_cr_n74), 
	.CK(hclk));
   DFFS_X2 U_cr_stmg1r_reg_17_ (.SN(FE_OFN63_HRESETn), 
	.QN(U_cr_n117), 
	.Q(cr_num_init_ref[1]), 
	.D(FE_PHN1520_U_cr_n75), 
	.CK(hclk));
   DFFS_X2 U_cr_stmg1r_reg_18_ (.SN(FE_OFN63_HRESETn), 
	.QN(U_cr_n116), 
	.Q(cr_num_init_ref[2]), 
	.D(FE_PHN1518_U_cr_n76), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg1r_reg_19_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n109), 
	.Q(cr_num_init_ref[3]), 
	.D(FE_PHN1082_U_cr_n77), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg1r_reg_20_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n53), 
	.Q(cr_t_wtr[0]), 
	.D(FE_PHN1517_U_cr_n78), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg1r_reg_21_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n60), 
	.Q(cr_t_wtr[1]), 
	.D(FE_PHN1516_U_cr_n79), 
	.CK(hclk));
   DFFS_X2 U_cr_stmg0r_reg_24_ (.SN(FE_OFN51_HRESETn), 
	.QN(n96), 
	.Q(cr_t_rc[2]), 
	.D(FE_PHN1168_U_cr_N413), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg0r_reg_25_ (.RN(FE_OFN51_HRESETn), 
	.Q(cr_t_rc[3]), 
	.D(FE_PHN698_U_cr_N414), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_stmg0r_reg_26_ (.RN(FE_OFN51_HRESETn), 
	.Q(U_cr_stmg0r_26), 
	.D(FE_PHN1116_U_cr_N415), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg0r_reg_27_ (.RN(FE_OFN28_HRESETn), 
	.Q(cr_t_xsr[4]), 
	.D(FE_PHN978_U_cr_N416), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_stmg0r_reg_28_ (.RN(FE_OFN28_HRESETn), 
	.Q(cr_t_xsr[5]), 
	.D(FE_PHN977_U_cr_N417), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_stmg0r_reg_29_ (.RN(FE_OFN53_HRESETn), 
	.Q(cr_t_xsr[6]), 
	.D(FE_PHN1076_U_cr_N418), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg0r_reg_30_ (.RN(FE_OFN53_HRESETn), 
	.Q(cr_t_xsr[7]), 
	.D(FE_PHN1040_U_cr_N419), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg0r_reg_31_ (.RN(FE_OFN53_HRESETn), 
	.Q(cr_t_xsr[8]), 
	.D(FE_PHN807_U_cr_N420), 
	.CK(HCLK__L5_N17));
   DFFS_X2 U_cr_stmg0r_reg_16_ (.SN(FE_OFN63_HRESETn), 
	.QN(U_cr_n104), 
	.Q(cr_t_rcar[2]), 
	.D(FE_PHN4627_U_cr_N405), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg0r_reg_17_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n72), 
	.Q(cr_t_rcar[3]), 
	.D(FE_PHN1617_U_cr_N406), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg0r_reg_18_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n108), 
	.Q(cr_t_xsr[0]), 
	.D(FE_PHN1526_U_cr_N407), 
	.CK(hclk));
   DFFS_X2 U_cr_stmg0r_reg_19_ (.SN(FE_OFN63_HRESETn), 
	.QN(U_cr_n32), 
	.Q(cr_t_xsr[1]), 
	.D(FE_PHN3220_U_cr_N408), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg0r_reg_20_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_cr_n33), 
	.Q(cr_t_xsr[2]), 
	.D(FE_PHN1523_U_cr_N409), 
	.CK(hclk));
   DFFS_X2 U_cr_stmg0r_reg_21_ (.SN(FE_OFN53_HRESETn), 
	.QN(U_cr_n34), 
	.Q(cr_t_xsr[3]), 
	.D(FE_PHN952_U_cr_N410), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg0r_reg_22_ (.RN(FE_OFN53_HRESETn), 
	.QN(U_cr_n64), 
	.D(FE_PHN889_U_cr_N411), 
	.CK(hclk));
   DFFS_X2 U_cr_stmg0r_reg_23_ (.SN(FE_OFN63_HRESETn), 
	.QN(U_cr_n106), 
	.Q(cr_t_rc[1]), 
	.D(FE_PHN1043_U_cr_N412), 
	.CK(hclk));
   DFFR_X1 U_cr_sconr_reg_16_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n28), 
	.Q(s_sa[1]), 
	.D(FE_PHN1514_U_cr_N311), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sconr_reg_17_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_cr_n31), 
	.Q(s_sa[2]), 
	.D(FE_PHN1240_U_cr_N312), 
	.CK(hclk));
   DFFS_X2 U_cr_sconr_reg_18_ (.SN(FE_OFN63_HRESETn), 
	.QN(U_cr_n30), 
	.Q(s_scl), 
	.D(FE_PHN1170_U_cr_N313), 
	.CK(hclk));
   DFFS_X2 U_cr_sconr_reg_20_ (.SN(FE_OFN51_HRESETn), 
	.QN(U_cr_n57), 
	.Q(s_sda_oe_n), 
	.D(FE_PHN2977_U_cr_N315), 
	.CK(hclk));
   DFFR_X1 U_cr_exn_mode_reg_reg_7_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_cr_n100), 
	.Q(cr_exn_mode_value[7]), 
	.D(FE_PHN1530_U_cr_N695), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_6_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_cr_n125), 
	.Q(cr_exn_mode_value[6]), 
	.D(FE_PHN1531_U_cr_N694), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_5_ (.RN(FE_OFN188_HRESETn), 
	.QN(U_cr_n124), 
	.Q(cr_exn_mode_value[5]), 
	.D(FE_PHN1702_U_cr_N693), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_4_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_cr_n26), 
	.Q(cr_exn_mode_value[4]), 
	.D(FE_PHN1382_U_cr_N692), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_3_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_cr_n97), 
	.Q(cr_exn_mode_value[3]), 
	.D(FE_PHN1703_U_cr_N691), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_2_ (.RN(FE_OFN35_HRESETn), 
	.Q(cr_exn_mode_value[2]), 
	.D(FE_PHN1567_U_cr_N690), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_1_ (.RN(FE_OFN151_HRESETn), 
	.Q(cr_exn_mode_value[1]), 
	.D(FE_PHN1638_U_cr_N689), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_0_ (.RN(FE_OFN35_HRESETn), 
	.Q(cr_exn_mode_value[0]), 
	.D(FE_PHN1643_U_cr_N688), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_smskr0_reg_7_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n167), 
	.Q(cr_block_size1[7]), 
	.D(FE_PHN3480_U_cr_n80), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_smskr0_reg_6_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n119), 
	.Q(cr_block_size1[6]), 
	.D(FE_PHN3230_U_cr_n81), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_smskr0_reg_5_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n110), 
	.Q(cr_block_size1[5]), 
	.D(FE_PHN1716_U_cr_n82), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_smskr0_reg_4_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n152), 
	.Q(U_cr_n554), 
	.D(FE_PHN1710_U_cr_n83), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_smskr0_reg_3_ (.SN(FE_OFN46_HRESETn), 
	.QN(U_cr_n165), 
	.Q(U_cr_n555), 
	.D(FE_PHN1176_U_cr_n84), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_smskr0_reg_2_ (.SN(FE_OFN46_HRESETn), 
	.Q(U_cr_n556), 
	.D(FE_PHN1409_U_cr_n85), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_smskr0_reg_1_ (.RN(FE_OFN46_HRESETn), 
	.Q(U_cr_n557), 
	.D(FE_PHN1647_U_cr_n86), 
	.CK(HCLK__L5_N35));
   DFFS_X2 U_cr_smskr0_reg_0_ (.SN(FE_OFN46_HRESETn), 
	.Q(U_cr_n558), 
	.D(FE_PHN3352_U_cr_n87), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_srefr_reg_7_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n113), 
	.Q(cr_t_ref[7]), 
	.D(FE_PHN1533_U_cr_N639), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_srefr_reg_6_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n121), 
	.Q(cr_t_ref[6]), 
	.D(FE_PHN1532_U_cr_N638), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_srefr_reg_5_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n112), 
	.Q(cr_t_ref[5]), 
	.D(FE_PHN1534_U_cr_N637), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_srefr_reg_4_ (.SN(FE_OFN46_HRESETn), 
	.QN(U_cr_n130), 
	.Q(cr_t_ref[4]), 
	.D(FE_PHN1713_U_cr_N636), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_srefr_reg_3_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n69), 
	.Q(cr_t_ref[3]), 
	.D(FE_PHN1714_U_cr_N635), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_srefr_reg_2_ (.RN(FE_OFN46_HRESETn), 
	.Q(cr_t_ref[2]), 
	.D(FE_PHN1412_U_cr_N634), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_sctlr_reg_7_ (.SN(FE_OFN59_HRESETn), 
	.QN(U_cr_n59), 
	.Q(s_read_pipe[1]), 
	.D(FE_PHN1745_U_cr_N557), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_sctlr_reg_6_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n40), 
	.Q(s_read_pipe[0]), 
	.D(FE_PHN1916_U_cr_N556), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_cr_sctlr_reg_5_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n132), 
	.Q(cr_ref_all_after_sr), 
	.D(FE_PHN1747_U_cr_N555), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_cr_sctlr_reg_4_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n139), 
	.Q(cr_ref_all_before_sr), 
	.D(FE_PHN1746_U_cr_N554), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_sctlr_reg_3_ (.SN(FE_OFN59_HRESETn), 
	.QN(U_cr_n58), 
	.Q(cr_delayed_precharge), 
	.D(FE_PHN1537_U_cr_N553), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sctlr_reg_2_ (.RN(FE_OFN148_HRESETn), 
	.Q(cr_do_power_down), 
	.D(FE_PHN1589_U_cr_N552), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sctlr_reg_1_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_cr_n39), 
	.Q(cr_do_self_ref_rp), 
	.D(FE_PHN3515_U_cr_N551), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_sctlr_reg_0_ (.SN(FE_OFN39_HRESETn), 
	.QN(U_cr_n56), 
	.Q(cr_do_initialize), 
	.D(FE_PHN1048_U_cr_N550), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg1r_reg_7_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n142), 
	.Q(cr_t_init[7]), 
	.D(FE_PHN1711_U_cr_N471), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg1r_reg_6_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_cr_n135), 
	.Q(cr_t_init[6]), 
	.D(FE_PHN1705_U_cr_N470), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_stmg1r_reg_5_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n141), 
	.Q(cr_t_init[5]), 
	.D(FE_PHN1704_U_cr_N469), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_stmg1r_reg_4_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_cr_n134), 
	.Q(cr_t_init[4]), 
	.D(FE_PHN1708_U_cr_N468), 
	.CK(HCLK__L5_N35));
   DFFS_X2 U_cr_stmg1r_reg_3_ (.SN(FE_OFN46_HRESETn), 
	.QN(U_cr_n150), 
	.Q(cr_t_init[3]), 
	.D(FE_PHN1384_U_cr_N467), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_stmg1r_reg_2_ (.RN(FE_OFN46_HRESETn), 
	.Q(cr_t_init[2]), 
	.D(FE_PHN1568_U_cr_N466), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_stmg1r_reg_1_ (.RN(FE_OFN172_HRESETn), 
	.Q(cr_t_init[1]), 
	.D(FE_PHN1845_U_cr_N465), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_stmg1r_reg_0_ (.RN(FE_OFN46_HRESETn), 
	.Q(cr_t_init[0]), 
	.D(FE_PHN1848_U_cr_N464), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_stmg0r_reg_7_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n133), 
	.Q(cr_t_rcd[1]), 
	.D(FE_PHN1734_U_cr_N396), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_stmg0r_reg_6_ (.SN(FE_OFN59_HRESETn), 
	.QN(U_cr_n149), 
	.Q(cr_t_rcd[0]), 
	.D(FE_PHN1735_U_cr_N395), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_cr_stmg0r_reg_5_ (.RN(FE_OFN187_HRESETn), 
	.QN(U_cr_n54), 
	.Q(cr_t_ras_min[3]), 
	.D(FE_PHN1736_U_cr_N394), 
	.CK(HCLK__L5_N28));
   DFFS_X2 U_cr_stmg0r_reg_4_ (.SN(FE_OFN188_HRESETn), 
	.QN(U_cr_n128), 
	.Q(cr_t_ras_min[2]), 
	.D(FE_PHN1388_U_cr_N393), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_cr_stmg0r_reg_3_ (.RN(FE_OFN36_HRESETn), 
	.QN(U_cr_n120), 
	.Q(cr_t_ras_min[1]), 
	.D(FE_PHN1739_U_cr_N392), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_cr_stmg0r_reg_2_ (.RN(FE_OFN36_HRESETn), 
	.QN(n95), 
	.Q(cr_t_ras_min[0]), 
	.D(FE_PHN1587_U_cr_N391), 
	.CK(HCLK__L5_N28));
   DFFS_X2 U_cr_cas_latency_o_reg_1_ (.SN(FE_OFN188_HRESETn), 
	.QN(n93), 
	.Q(s_cas_latency[1]), 
	.D(FE_PHN3287_U_cr_N576), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_cr_stmg0r_reg_1_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n43), 
	.Q(U_cr_stmg0r_1_), 
	.D(FE_PHN1737_U_cr_N390), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_stmg0r_reg_0_ (.SN(FE_OFN59_HRESETn), 
	.QN(U_cr_n20), 
	.Q(U_cr_stmg0r_0_), 
	.D(FE_PHN1913_U_cr_N389), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_sconr_reg_7_ (.SN(FE_OFN151_HRESETn), 
	.QN(U_cr_n55), 
	.Q(cr_row_addr_width[2]), 
	.D(FE_PHN4645_U_cr_N302), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_sconr_reg_6_ (.RN(FE_OFN36_HRESETn), 
	.QN(U_cr_n42), 
	.Q(cr_row_addr_width[1]), 
	.D(FE_PHN1706_U_cr_N301), 
	.CK(HCLK__L5_N28));
   DFFR_X1 U_cr_sconr_reg_5_ (.RN(FE_OFN188_HRESETn), 
	.QN(U_cr_n21), 
	.Q(cr_row_addr_width[0]), 
	.D(FE_PHN1700_U_cr_N300), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_sconr_reg_4_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_cr_n66), 
	.Q(cr_bank_addr_width[1]), 
	.D(FE_PHN1699_U_cr_N299), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_sconr_reg_3_ (.SN(FE_OFN35_HRESETn), 
	.QN(U_cr_n36), 
	.Q(cr_bank_addr_width[0]), 
	.D(FE_PHN988_U_cr_N298), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_7_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_cr_n159), 
	.Q(U_cr_n563), 
	.D(FE_PHN1707_U_cr_N740), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_6_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_cr_n158), 
	.Q(U_cr_n564), 
	.D(FE_PHN1709_U_cr_N739), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_5_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n157), 
	.Q(U_cr_n565), 
	.D(FE_PHN1712_U_cr_N738), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_4_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n164), 
	.Q(U_cr_n566), 
	.D(FE_PHN1701_U_cr_N737), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_3_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n156), 
	.Q(U_cr_n567), 
	.D(FE_PHN1383_U_cr_N736), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_2_ (.RN(FE_OFN151_HRESETn), 
	.Q(U_cr_n568), 
	.D(FE_PHN1569_U_cr_N735), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_1_ (.RN(FE_OFN151_HRESETn), 
	.Q(U_cr_n569), 
	.D(FE_PHN1637_U_cr_N734), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_0_ (.RN(FE_OFN151_HRESETn), 
	.Q(U_cr_n570), 
	.D(FE_PHN1639_U_cr_N733), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_8_ (.RN(FE_OFN188_HRESETn), 
	.QN(U_cr_n161), 
	.Q(U_cr_n562), 
	.D(FE_PHN1528_U_cr_n88), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_9_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n162), 
	.Q(U_cr_n561), 
	.D(FE_PHN1694_U_cr_n89), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_11_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n163), 
	.Q(U_cr_n560), 
	.D(FE_PHN1693_U_cr_n91), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_syflash_opcode_reg_12_ (.RN(FE_OFN188_HRESETn), 
	.QN(U_cr_n160), 
	.Q(U_cr_n571), 
	.D(FE_PHN1692_U_cr_N745), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_12_ (.RN(FE_OFN188_HRESETn), 
	.QN(U_cr_n103), 
	.Q(cr_exn_mode_value[12]), 
	.D(FE_PHN1695_U_cr_N700), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_11_ (.RN(FE_OFN188_HRESETn), 
	.QN(U_cr_n102), 
	.Q(cr_exn_mode_value[11]), 
	.D(FE_PHN1380_U_cr_N699), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_10_ (.RN(FE_OFN188_HRESETn), 
	.QN(U_cr_n71), 
	.Q(cr_exn_mode_value[10]), 
	.D(FE_PHN1696_U_cr_N698), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_9_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_cr_n101), 
	.Q(cr_exn_mode_value[9]), 
	.D(FE_PHN1697_U_cr_N697), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_exn_mode_reg_reg_8_ (.RN(FE_OFN189_HRESETn), 
	.QN(U_cr_n126), 
	.Q(cr_exn_mode_value[8]), 
	.D(FE_PHN1698_U_cr_N696), 
	.CK(HCLK__L5_N28));
   DFFS_X2 U_cr_smskr0_reg_9_ (.SN(FE_OFN46_HRESETn), 
	.QN(U_cr_n166), 
	.Q(U_cr_n552), 
	.D(FE_PHN982_U_cr_n93), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_srefr_reg_15_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_cr_n114), 
	.Q(cr_t_ref[15]), 
	.D(FE_PHN1722_U_cr_N647), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_srefr_reg_14_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_cr_n123), 
	.Q(cr_t_ref[14]), 
	.D(FE_PHN1444_U_cr_N646), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_srefr_reg_13_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_cr_n68), 
	.Q(cr_t_ref[13]), 
	.D(FE_PHN1124_U_cr_N645), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_srefr_reg_12_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_cr_n122), 
	.Q(cr_t_ref[12]), 
	.D(FE_PHN1723_U_cr_N644), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_srefr_reg_11_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_cr_n111), 
	.Q(cr_t_ref[11]), 
	.D(FE_PHN1720_U_cr_N643), 
	.CK(HCLK__L5_N35));
   DFFS_X2 U_cr_srefr_reg_10_ (.SN(FE_OFN31_HRESETn), 
	.QN(U_cr_n129), 
	.Q(cr_t_ref[10]), 
	.D(FE_PHN1715_U_cr_N642), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_srefr_reg_9_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n105), 
	.Q(cr_t_ref[9]), 
	.D(FE_PHN1721_U_cr_N641), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_srefr_reg_8_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_cr_n118), 
	.Q(cr_t_ref[8]), 
	.D(FE_PHN1718_U_cr_N640), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_cr_sctlr_reg_15_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_cr_n44), 
	.Q(U_cr_sctlr_15_), 
	.D(FE_PHN1740_U_cr_N564), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sctlr_reg_14_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_cr_n35), 
	.Q(U_cr_sctlr_14_), 
	.D(FE_PHN1733_U_cr_N563), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_sctlr_reg_13_ (.SN(FE_OFN39_HRESETn), 
	.QN(U_cr_n27), 
	.Q(U_cr_sctlr_13_), 
	.D(FE_PHN3237_U_cr_N562), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_sctlr_reg_12_ (.SN(FE_OFN59_HRESETn), 
	.QN(U_cr_n18), 
	.Q(U_cr_sctlr_12_), 
	.D(FE_PHN1449_U_cr_N561), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sctlr_reg_10_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n155), 
	.Q(U_cr_n559), 
	.D(FE_PHN1731_U_cr_N560), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sctlr_reg_9_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n61), 
	.Q(cr_mode_reg_update), 
	.D(FE_PHN957_U_cr_N559), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sctlr_reg_8_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n41), 
	.Q(s_read_pipe[2]), 
	.D(FE_PHN1726_U_cr_N558), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg1r_reg_15_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n146), 
	.Q(cr_t_init[15]), 
	.D(FE_PHN1732_U_cr_N479), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg1r_reg_14_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_cr_n138), 
	.Q(cr_t_init[14]), 
	.D(FE_PHN1536_U_cr_N478), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg1r_reg_13_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_cr_n145), 
	.Q(cr_t_init[13]), 
	.D(FE_PHN1535_U_cr_N477), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg1r_reg_12_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_cr_n131), 
	.Q(cr_t_init[12]), 
	.D(FE_PHN1719_U_cr_N476), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg1r_reg_11_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_cr_n144), 
	.Q(cr_t_init[11]), 
	.D(FE_PHN1728_U_cr_N475), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg1r_reg_10_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_cr_n137), 
	.Q(cr_t_init[10]), 
	.D(FE_PHN1386_U_cr_N474), 
	.CK(hclk));
   DFFR_X1 U_cr_stmg1r_reg_9_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_cr_n143), 
	.Q(cr_t_init[9]), 
	.D(FE_PHN1727_U_cr_N473), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg1r_reg_8_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_cr_n136), 
	.Q(cr_t_init[8]), 
	.D(FE_PHN1730_U_cr_N472), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_stmg0r_reg_15_ (.SN(FE_OFN63_HRESETn), 
	.QN(U_cr_n151), 
	.Q(cr_t_rcar[1]), 
	.D(FE_PHN4913_U_cr_N404), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_stmg0r_reg_14_ (.SN(FE_OFN63_HRESETn), 
	.QN(U_cr_n127), 
	.Q(cr_t_rcar[0]), 
	.D(FE_PHN4736_U_cr_N403), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg0r_reg_13_ (.RN(FE_OFN63_HRESETn), 
	.QN(U_cr_n67), 
	.Q(cr_t_wr[1]), 
	.D(FE_PHN1738_U_cr_N402), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_stmg0r_reg_12_ (.SN(FE_OFN39_HRESETn), 
	.QN(U_cr_n107), 
	.Q(cr_t_wr[0]), 
	.D(FE_PHN1387_U_cr_N401), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg0r_reg_11_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n148), 
	.Q(cr_t_rp[2]), 
	.D(FE_PHN1725_U_cr_N400), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_stmg0r_reg_10_ (.SN(FE_OFN59_HRESETn), 
	.QN(U_cr_n147), 
	.Q(cr_t_rp[1]), 
	.D(FE_PHN1911_U_cr_N399), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg0r_reg_9_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n45), 
	.Q(cr_t_rp[0]), 
	.D(FE_PHN1724_U_cr_N398), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_stmg0r_reg_8_ (.RN(FE_OFN59_HRESETn), 
	.QN(U_cr_n140), 
	.Q(cr_t_rcd[2]), 
	.D(FE_PHN1729_U_cr_N397), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_cr_sconr_reg_15_ (.RN(FE_OFN172_HRESETn), 
	.QN(U_cr_n52), 
	.Q(s_sa[0]), 
	.D(FE_PHN1456_U_cr_N310), 
	.CK(hclk));
   DFFS_X2 U_cr_sdram_data_width_reg_0_ (.SN(FE_OFN31_HRESETn), 
	.QN(U_cr_n17), 
	.Q(n27), 
	.D(U_cr_n95), 
	.CK(HCLK__L5_N17));
   DFFS_X2 U_cr_sconr_reg_13_ (.SN(FE_OFN51_HRESETn), 
	.QN(n85), 
	.Q(cr_s_data_width_early_0_), 
	.D(U_cr_N308), 
	.CK(hclk));
   DFFS_X2 U_cr_sconr_reg_12_ (.SN(FE_OFN35_HRESETn), 
	.QN(U_cr_n65), 
	.Q(n[23]), 
	.D(FE_PHN1252_U_cr_N307), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_sconr_reg_11_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_cr_n38), 
	.Q(n[24]), 
	.D(FE_PHN1253_U_cr_N306), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_sconr_reg_10_ (.SN(FE_OFN35_HRESETn), 
	.QN(U_cr_n22), 
	.Q(n[25]), 
	.D(FE_PHN1127_U_cr_N305), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_cr_sconr_reg_9_ (.SN(FE_OFN35_HRESETn), 
	.QN(U_cr_n63), 
	.Q(n[26]), 
	.D(FE_PHN1917_U_cr_N304), 
	.CK(HCLK__L5_N34));
   DFFS_X2 U_cr_sconr_reg_8_ (.SN(FE_OFN151_HRESETn), 
	.QN(U_cr_n70), 
	.Q(cr_row_addr_width[3]), 
	.D(FE_PHN1455_U_cr_N303), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_cr_s_sda_d_reg (.RN(FE_OFN51_HRESETn), 
	.Q(U_cr_s_sda_d), 
	.D(s_sda_in), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_srefr_reg_24_ (.RN(FE_OFN51_HRESETn), 
	.Q(U_cr_srefr[24]), 
	.D(gpi[0]), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_srefr_reg_25_ (.RN(FE_OFN51_HRESETn), 
	.Q(U_cr_srefr[25]), 
	.D(gpi[1]), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_srefr_reg_26_ (.RN(FE_OFN51_HRESETn), 
	.Q(U_cr_srefr[26]), 
	.D(gpi[2]), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_srefr_reg_27_ (.RN(FE_OFN28_HRESETn), 
	.Q(U_cr_srefr[27]), 
	.D(gpi[3]), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_srefr_reg_28_ (.RN(FE_OFN28_HRESETn), 
	.Q(U_cr_srefr[28]), 
	.D(gpi[4]), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_srefr_reg_29_ (.RN(FE_OFN28_HRESETn), 
	.Q(U_cr_srefr[29]), 
	.D(gpi[5]), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_srefr_reg_30_ (.RN(FE_OFN28_HRESETn), 
	.Q(U_cr_srefr[30]), 
	.D(gpi[6]), 
	.CK(HCLK__L5_N17));
   DFFR_X1 U_cr_srefr_reg_31_ (.RN(FE_OFN51_HRESETn), 
	.Q(U_cr_srefr[31]), 
	.D(gpi[7]), 
	.CK(HCLK__L5_N17));
   DFFS_X2 U_cr_open_banks_o_reg_0_ (.SN(FE_OFN59_HRESETn), 
	.Q(cr_num_open_banks[0]), 
	.D(FE_PHN4617_U_cr_n18), 
	.CK(HCLK__L5_N11));
   DFFS_X2 U_cr_open_banks_o_reg_1_ (.SN(FE_OFN39_HRESETn), 
	.Q(cr_num_open_banks[1]), 
	.D(FE_PHN1555_U_cr_N571), 
	.CK(HCLK__L5_N11));
   NAND2_X2 U_addrdec_U359 (.ZN(U_addrdec_n113), 
	.A2(U_addrdec_n21), 
	.A1(U_addrdec_n16));
   NAND2_X2 U_addrdec_U358 (.ZN(U_addrdec_n105), 
	.A2(U_addrdec_bcawp_1_), 
	.A1(U_addrdec_bcawp_2_));
   NAND2_X2 U_addrdec_U357 (.ZN(U_addrdec_n114), 
	.A2(U_addrdec_bcawp_3_), 
	.A1(U_addrdec_n101));
   MUX2_X2 U_addrdec_U356 (.Z(U_addrdec_n84), 
	.S(n[25]), 
	.B(debug_ad_col_addr_13_), 
	.A(U_addrdec_n79));
   AND2_X4 U_addrdec_U355 (.ZN(debug_ad_row_addr[13]), 
	.A2(U_addrdec_row_addr_mask[13]), 
	.A1(U_addrdec_n253));
   OAI211_X2 U_addrdec_U354 (.ZN(U_addrdec_n94), 
	.C2(U_addrdec_n80), 
	.C1(n[23]), 
	.B(U_addrdec_bank_addr_mask_1_), 
	.A(U_addrdec_n78));
   NOR2_X2 U_addrdec_U353 (.ZN(U_addrdec_n86), 
	.A2(n[26]), 
	.A1(U_addrdec_n80));
   AND2_X4 U_addrdec_U352 (.ZN(debug_ad_row_addr[15]), 
	.A2(U_addrdec_row_addr_mask[15]), 
	.A1(U_addrdec_n278));
   NAND2_X2 U_addrdec_U351 (.ZN(debug_ad_col_addr_8_), 
	.A2(U_addrdec_n43), 
	.A1(U_addrdec_n44));
   AND2_X4 U_addrdec_U350 (.ZN(U_addrdec_n32), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[12]));
   NOR2_X2 U_addrdec_U349 (.ZN(U_addrdec_n28), 
	.A2(U_addrdec_n113), 
	.A1(U_addrdec_n117));
   AND2_X4 U_addrdec_U348 (.ZN(U_addrdec_n27), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[13]));
   NOR2_X2 U_addrdec_U347 (.ZN(U_addrdec_n26), 
	.A2(U_addrdec_n105), 
	.A1(U_addrdec_n117));
   OR2_X4 U_addrdec_U346 (.ZN(U_addrdec_n24), 
	.A2(U_addrdec_n105), 
	.A1(U_addrdec_n114));
   OR2_X4 U_addrdec_U345 (.ZN(U_addrdec_n23), 
	.A2(U_addrdec_n113), 
	.A1(U_addrdec_n114));
   OR2_X4 U_addrdec_U344 (.ZN(U_addrdec_n22), 
	.A2(U_addrdec_n115), 
	.A1(U_addrdec_n117));
   NOR3_X2 U_addrdec_U343 (.ZN(U_addrdec_n18), 
	.A3(U_addrdec_bcawp_3_), 
	.A2(U_addrdec_n105), 
	.A1(U_addrdec_n106));
   AND2_X4 U_addrdec_U342 (.ZN(U_addrdec_n13), 
	.A2(U_addrdec_n103), 
	.A1(U_addrdec_n104));
   NOR2_X2 U_addrdec_U341 (.ZN(U_addrdec_n272), 
	.A2(U_addrdec_n115), 
	.A1(U_addrdec_n114));
   NOR3_X2 U_addrdec_U340 (.ZN(U_addrdec_n74), 
	.A3(U_cr_n63), 
	.A2(n[23]), 
	.A1(U_addrdec_n67));
   NOR2_X2 U_addrdec_U339 (.ZN(U_addrdec_n81), 
	.A2(n[25]), 
	.A1(U_cr_n38));
   NOR2_X2 U_addrdec_U338 (.ZN(U_addrdec_n92), 
	.A2(U_addrdec_n90), 
	.A1(U_addrdec_n91));
   AOI21_X2 U_addrdec_U337 (.ZN(U_addrdec_n73), 
	.B2(n[26]), 
	.B1(U_addrdec_n59), 
	.A(U_addrdec_n57));
   AOI22_X2 U_addrdec_U336 (.ZN(U_addrdec_n70), 
	.B2(U_addrdec_n75), 
	.B1(debug_ad_col_addr_15_), 
	.A2(debug_ad_col_addr_8_), 
	.A1(U_addrdec_n74));
   AND2_X4 U_addrdec_U335 (.ZN(debug_ad_row_addr[14]), 
	.A2(U_addrdec_row_addr_mask[14]), 
	.A1(U_addrdec_n263));
   AOI22_X1 U_addrdec_U332 (.ZN(U_addrdec_n100), 
	.B2(U_addrdec_n39), 
	.B1(hiu_addr[7]), 
	.A2(hiu_addr[8]), 
	.A1(U_addrdec_n220));
   XNOR2_X2 U_addrdec_U331 (.ZN(U_addrdec_N108), 
	.B(U_addrdec_n286), 
	.A(FE_PHN1034_cr_bank_addr_width_1_));
   NAND2_X2 U_addrdec_U329 (.ZN(U_addrdec_n106), 
	.A2(U_addrdec_bcawp_0_), 
	.A1(U_addrdec_n15));
   NAND2_X2 U_addrdec_U328 (.ZN(U_addrdec_n115), 
	.A2(U_addrdec_bcawp_1_), 
	.A1(U_addrdec_n16));
   INV_X4 U_addrdec_U325 (.ZN(U_addrdec_n180), 
	.A(U_addrdec_n102));
   NAND3_X2 U_addrdec_U324 (.ZN(U_addrdec_n117), 
	.A3(U_addrdec_bcawp_3_), 
	.A2(U_addrdec_n15), 
	.A1(U_addrdec_n20));
   NAND2_X2 U_addrdec_U323 (.ZN(U_addrdec_n116), 
	.A2(U_addrdec_bcawp_2_), 
	.A1(U_addrdec_n21));
   NOR2_X2 U_addrdec_U322 (.ZN(U_addrdec_n17), 
	.A2(U_addrdec_n116), 
	.A1(U_addrdec_n117));
   INV_X4 U_addrdec_U321 (.ZN(U_addrdec_n161), 
	.A(U_addrdec_n17));
   OAI22_X2 U_addrdec_U320 (.ZN(U_addrdec_n136), 
	.B2(U_addrdec_n130), 
	.B1(U_addrdec_n13), 
	.A2(U_addrdec_n161), 
	.A1(U_addrdec_n180));
   NAND2_X2 U_addrdec_U319 (.ZN(U_addrdec_n107), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[20]));
   NAND2_X2 U_addrdec_U318 (.ZN(U_addrdec_n181), 
	.A2(U_addrdec_n107), 
	.A1(U_addrdec_n108));
   INV_X4 U_addrdec_U317 (.ZN(U_addrdec_n35), 
	.A(U_addrdec_n24));
   AOI22_X2 U_addrdec_U316 (.ZN(U_addrdec_n134), 
	.B2(U_addrdec_n35), 
	.B1(U_addrdec_n181), 
	.A2(U_addrdec_n34), 
	.A1(FE_OFN360_U_addrdec_n26));
   NAND2_X2 U_addrdec_U315 (.ZN(U_addrdec_n132), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[22]));
   NAND2_X2 U_addrdec_U314 (.ZN(U_addrdec_n131), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[21]));
   NAND2_X2 U_addrdec_U313 (.ZN(U_addrdec_n232), 
	.A2(U_addrdec_n131), 
	.A1(U_addrdec_n132));
   NAND2_X2 U_addrdec_U312 (.ZN(U_addrdec_n122), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[20]));
   NAND2_X2 U_addrdec_U311 (.ZN(U_addrdec_n121), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[21]));
   INV_X4 U_addrdec_U310 (.ZN(U_addrdec_n36), 
	.A(U_addrdec_n25));
   AOI22_X2 U_addrdec_U309 (.ZN(U_addrdec_n133), 
	.B2(U_addrdec_n36), 
	.B1(U_addrdec_n219), 
	.A2(U_addrdec_n232), 
	.A1(U_addrdec_n30));
   NAND2_X2 U_addrdec_U308 (.ZN(U_addrdec_n135), 
	.A2(U_addrdec_n133), 
	.A1(U_addrdec_n134));
   AOI211_X2 U_addrdec_U307 (.ZN(U_addrdec_n139), 
	.C2(debug_ad_col_addr_15_), 
	.C1(U_addrdec_n272), 
	.B(U_addrdec_n135), 
	.A(U_addrdec_n136));
   INV_X4 U_addrdec_U306 (.ZN(debug_ad_col_addr_12__BAR_BAR), 
	.A(debug_ad_col_addr_12_));
   NAND2_X2 U_addrdec_U305 (.ZN(U_addrdec_n54), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[12]));
   AOI22_X2 U_addrdec_U304 (.ZN(U_addrdec_n138), 
	.B2(U_addrdec_n18), 
	.B1(debug_ad_col_addr_11_), 
	.A2(U_addrdec_n28), 
	.A1(debug_ad_col_addr_12__BAR_BAR));
   INV_X4 U_addrdec_U303 (.ZN(U_addrdec_n37), 
	.A(U_addrdec_n23));
   INV_X4 U_addrdec_U299 (.ZN(U_addrdec_n38), 
	.A(U_addrdec_n22));
   AOI22_X2 U_addrdec_U298 (.ZN(U_addrdec_n137), 
	.B2(U_addrdec_n38), 
	.B1(debug_ad_col_addr_14_), 
	.A2(U_addrdec_n37), 
	.A1(debug_ad_col_addr_13__BAR_BAR));
   NAND3_X2 U_addrdec_U297 (.ZN(debug_ad_row_addr[2]), 
	.A3(U_addrdec_n137), 
	.A2(U_addrdec_n138), 
	.A1(U_addrdec_n139));
   INV_X4 U_addrdec_U296 (.ZN(U_addrdec_n310), 
	.A(hiu_mem_req));
   OAI22_X2 U_addrdec_U295 (.ZN(U_addrdec_n126), 
	.B2(U_addrdec_n256), 
	.B1(U_addrdec_n13), 
	.A2(U_addrdec_n130), 
	.A1(U_addrdec_n180));
   AOI22_X2 U_addrdec_U294 (.ZN(U_addrdec_n124), 
	.B2(U_addrdec_n30), 
	.B1(U_addrdec_n219), 
	.A2(U_addrdec_n34), 
	.A1(U_addrdec_n35));
   AOI22_X2 U_addrdec_U293 (.ZN(U_addrdec_n123), 
	.B2(U_addrdec_n36), 
	.B1(U_addrdec_n181), 
	.A2(debug_ad_col_addr_11_), 
	.A1(U_addrdec_n28));
   NAND2_X2 U_addrdec_U292 (.ZN(U_addrdec_n125), 
	.A2(U_addrdec_n123), 
	.A1(U_addrdec_n124));
   AOI211_X2 U_addrdec_U291 (.ZN(U_addrdec_n129), 
	.C2(debug_ad_col_addr_15_), 
	.C1(U_addrdec_n17), 
	.B(U_addrdec_n125), 
	.A(U_addrdec_n126));
   AOI22_X2 U_addrdec_U288 (.ZN(U_addrdec_n128), 
	.B2(U_addrdec_n18), 
	.B1(debug_ad_col_addr_10_), 
	.A2(U_addrdec_n37), 
	.A1(debug_ad_col_addr_12__BAR_BAR));
   AOI22_X2 U_addrdec_U287 (.ZN(U_addrdec_n127), 
	.B2(U_addrdec_n272), 
	.B1(debug_ad_col_addr_14_), 
	.A2(U_addrdec_n38), 
	.A1(FE_OFN211_debug_ad_col_addr_13_));
   NAND3_X2 U_addrdec_U286 (.ZN(debug_ad_row_addr[1]), 
	.A3(U_addrdec_n127), 
	.A2(U_addrdec_n128), 
	.A1(U_addrdec_n129));
   INV_X4 U_addrdec_U285 (.ZN(U_addrdec_n79), 
	.A(debug_ad_col_addr_11_));
   NAND2_X2 U_addrdec_U282 (.ZN(U_addrdec_n67), 
	.A2(n[25]), 
	.A1(n[24]));
   NAND2_X2 U_addrdec_U280 (.ZN(U_addrdec_n77), 
	.A2(U_addrdec_n74), 
	.A1(debug_ad_col_addr_9_));
   NAND2_X2 U_addrdec_U276 (.ZN(U_addrdec_n76), 
	.A2(U_addrdec_n75), 
	.A1(U_addrdec_n102));
   NAND2_X2 U_addrdec_U275 (.ZN(U_addrdec_n80), 
	.A2(U_addrdec_n76), 
	.A1(U_addrdec_n77));
   NOR2_X2 U_addrdec_U274 (.ZN(U_addrdec_n83), 
	.A2(U_cr_n63), 
	.A1(U_addrdec_n80));
   NAND2_X2 U_addrdec_U273 (.ZN(U_addrdec_n82), 
	.A2(U_addrdec_n81), 
	.A1(debug_ad_col_addr_15_));
   INV_X4 U_addrdec_U272 (.ZN(U_addrdec_n93), 
	.A(U_addrdec_n85));
   NAND2_X2 U_addrdec_U271 (.ZN(U_addrdec_n88), 
	.A2(U_addrdec_n81), 
	.A1(debug_ad_col_addr_14_));
   NAND3_X2 U_addrdec_U270 (.ZN(U_addrdec_n78), 
	.A3(U_addrdec_n88), 
	.A2(n[24]), 
	.A1(U_addrdec_n86));
   NAND2_X2 U_addrdec_U269 (.ZN(U_addrdec_n87), 
	.A2(U_cr_n22), 
	.A1(debug_ad_col_addr_10_));
   OAI211_X2 U_addrdec_U268 (.ZN(U_addrdec_n90), 
	.C2(U_cr_n22), 
	.C1(debug_ad_col_addr_12_), 
	.B(U_addrdec_n87), 
	.A(U_addrdec_n88));
   NOR3_X2 U_addrdec_U267 (.ZN(n44), 
	.A3(U_addrdec_n92), 
	.A2(U_addrdec_n94), 
	.A1(U_addrdec_n93));
   NOR3_X2 U_addrdec_U266 (.ZN(U_addrdec_n57), 
	.A3(U_addrdec_n56), 
	.A2(n[26]), 
	.A1(debug_ad_col_addr_13_));
   NOR3_X2 U_addrdec_U265 (.ZN(U_addrdec_n60), 
	.A3(U_cr_n22), 
	.A2(U_cr_n63), 
	.A1(debug_ad_col_addr_12__BAR_BAR));
   NOR3_X2 U_addrdec_U264 (.ZN(U_addrdec_n66), 
	.A3(FE_PHN1645_U_cr_n65), 
	.A2(n[24]), 
	.A1(U_addrdec_n60));
   NAND3_X2 U_addrdec_U263 (.ZN(U_addrdec_n65), 
	.A3(U_cr_n63), 
	.A2(n[25]), 
	.A1(U_addrdec_n79));
   NAND3_X2 U_addrdec_U262 (.ZN(U_addrdec_n64), 
	.A3(U_cr_n22), 
	.A2(U_cr_n63), 
	.A1(U_addrdec_n61));
   NAND3_X2 U_addrdec_U261 (.ZN(U_addrdec_n63), 
	.A3(U_cr_n22), 
	.A2(n[26]), 
	.A1(U_addrdec_n62));
   NAND4_X2 U_addrdec_U260 (.ZN(U_addrdec_n71), 
	.A4(U_addrdec_n63), 
	.A3(U_addrdec_n64), 
	.A2(U_addrdec_n65), 
	.A1(U_addrdec_n66));
   NAND2_X2 U_addrdec_U259 (.ZN(U_addrdec_n44), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[9]));
   NAND2_X2 U_addrdec_U258 (.ZN(U_addrdec_n43), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[8]));
   NAND2_X2 U_addrdec_U257 (.ZN(U_addrdec_n141), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[23]));
   NAND2_X2 U_addrdec_U256 (.ZN(U_addrdec_n140), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[22]));
   NAND2_X2 U_addrdec_U255 (.ZN(U_addrdec_n242), 
	.A2(U_addrdec_n140), 
	.A1(U_addrdec_n141));
   AOI22_X2 U_addrdec_U254 (.ZN(U_addrdec_n226), 
	.B2(U_addrdec_n37), 
	.B1(U_addrdec_n242), 
	.A2(U_addrdec_n219), 
	.A1(U_addrdec_n18));
   NAND2_X2 U_addrdec_U253 (.ZN(U_addrdec_n156), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[24]));
   NAND2_X2 U_addrdec_U252 (.ZN(U_addrdec_n155), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[23]));
   NAND2_X2 U_addrdec_U251 (.ZN(U_addrdec_n254), 
	.A2(U_addrdec_n155), 
	.A1(U_addrdec_n156));
   NAND2_X2 U_addrdec_U250 (.ZN(U_addrdec_n167), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[25]));
   NAND2_X2 U_addrdec_U249 (.ZN(U_addrdec_n166), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[24]));
   NAND2_X2 U_addrdec_U248 (.ZN(U_addrdec_n264), 
	.A2(U_addrdec_n166), 
	.A1(U_addrdec_n167));
   AOI22_X2 U_addrdec_U247 (.ZN(U_addrdec_n225), 
	.B2(U_addrdec_n272), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n254), 
	.A1(U_addrdec_n38));
   NAND2_X2 U_addrdec_U246 (.ZN(U_addrdec_n270), 
	.A2(U_addrdec_n221), 
	.A1(U_addrdec_n222));
   AOI22_X2 U_addrdec_U245 (.ZN(U_addrdec_n224), 
	.B2(U_addrdec_n30), 
	.B1(U_addrdec_n270), 
	.A2(U_addrdec_n28), 
	.A1(U_addrdec_n232));
   NAND4_X2 U_addrdec_U244 (.ZN(U_addrdec_n230), 
	.A4(U_addrdec_n223), 
	.A3(U_addrdec_n224), 
	.A2(U_addrdec_n225), 
	.A1(U_addrdec_n226));
   NAND2_X2 U_addrdec_U243 (.ZN(U_addrdec_n176), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[25]));
   NAND2_X2 U_addrdec_U242 (.ZN(U_addrdec_n265), 
	.A2(U_addrdec_n175), 
	.A1(U_addrdec_n176));
   NAND2_X2 U_addrdec_U241 (.ZN(U_addrdec_n267), 
	.A2(U_addrdec_n195), 
	.A1(U_addrdec_n196));
   AOI22_X2 U_addrdec_U240 (.ZN(U_addrdec_n228), 
	.B2(U_addrdec_n26), 
	.B1(U_addrdec_n267), 
	.A2(U_addrdec_n265), 
	.A1(U_addrdec_n17));
   NAND2_X2 U_addrdec_U239 (.ZN(U_addrdec_n273), 
	.A2(U_addrdec_n205), 
	.A1(U_addrdec_n206));
   NAND2_X2 U_addrdec_U238 (.ZN(U_addrdec_n266), 
	.A2(U_addrdec_n186), 
	.A1(U_addrdec_n187));
   AOI22_X2 U_addrdec_U237 (.ZN(U_addrdec_n227), 
	.B2(U_addrdec_n269), 
	.B1(U_addrdec_n266), 
	.A2(U_addrdec_n273), 
	.A1(U_addrdec_n35));
   NAND2_X2 U_addrdec_U236 (.ZN(U_addrdec_n229), 
	.A2(U_addrdec_n227), 
	.A1(U_addrdec_n228));
   OAI21_X2 U_addrdec_U235 (.ZN(U_addrdec_n231), 
	.B2(U_addrdec_n229), 
	.B1(U_addrdec_n230), 
	.A(U_addrdec_row_addr_mask[11]));
   INV_X4 U_addrdec_U234 (.ZN(debug_ad_row_addr[11]), 
	.A(U_addrdec_n231));
   INV_X4 U_addrdec_U233 (.ZN(U_addrdec_n245), 
	.A(U_addrdec_n18));
   INV_X4 U_addrdec_U232 (.ZN(U_addrdec_n210), 
	.A(U_addrdec_n181));
   INV_X4 U_addrdec_U231 (.ZN(U_addrdec_n243), 
	.A(U_addrdec_n28));
   OAI22_X2 U_addrdec_U230 (.ZN(U_addrdec_n204), 
	.B2(U_addrdec_n243), 
	.B1(U_addrdec_n210), 
	.A2(U_addrdec_n245), 
	.A1(U_addrdec_n200));
   AOI22_X2 U_addrdec_U229 (.ZN(U_addrdec_n202), 
	.B2(U_addrdec_n272), 
	.B1(U_addrdec_n242), 
	.A2(U_addrdec_n219), 
	.A1(U_addrdec_n37));
   AOI22_X2 U_addrdec_U228 (.ZN(U_addrdec_n201), 
	.B2(U_addrdec_n17), 
	.B1(U_addrdec_n254), 
	.A2(U_addrdec_n232), 
	.A1(U_addrdec_n38));
   NAND2_X2 U_addrdec_U227 (.ZN(U_addrdec_n203), 
	.A2(U_addrdec_n201), 
	.A1(U_addrdec_n202));
   AOI211_X2 U_addrdec_U226 (.ZN(U_addrdec_n209), 
	.C2(U_addrdec_n267), 
	.C1(U_addrdec_n36), 
	.B(U_addrdec_n203), 
	.A(U_addrdec_n204));
   AOI22_X2 U_addrdec_U225 (.ZN(U_addrdec_n208), 
	.B2(U_addrdec_n269), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n265), 
	.A1(U_addrdec_n26));
   AOI22_X2 U_addrdec_U224 (.ZN(U_addrdec_n207), 
	.B2(U_addrdec_n35), 
	.B1(U_addrdec_n266), 
	.A2(U_addrdec_n273), 
	.A1(U_addrdec_n30));
   NAND3_X2 U_addrdec_U223 (.ZN(debug_ad_row_addr[9]), 
	.A3(U_addrdec_n207), 
	.A2(U_addrdec_n208), 
	.A1(U_addrdec_n209));
   OAI22_X2 U_addrdec_U222 (.ZN(U_addrdec_n165), 
	.B2(U_addrdec_n161), 
	.B1(U_addrdec_n210), 
	.A2(U_addrdec_n23), 
	.A1(U_addrdec_n180));
   AOI22_X2 U_addrdec_U221 (.ZN(U_addrdec_n163), 
	.B2(U_addrdec_n269), 
	.B1(U_addrdec_n219), 
	.A2(U_addrdec_n232), 
	.A1(U_addrdec_n26));
   OAI211_X2 U_addrdec_U220 (.ZN(U_addrdec_n164), 
	.C2(U_addrdec_n22), 
	.C1(U_addrdec_n13), 
	.B(U_addrdec_n162), 
	.A(U_addrdec_n163));
   AOI22_X2 U_addrdec_U219 (.ZN(U_addrdec_n169), 
	.B2(U_addrdec_n30), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n242), 
	.A1(U_addrdec_n35));
   AOI22_X2 U_addrdec_U218 (.ZN(U_addrdec_n168), 
	.B2(U_addrdec_n36), 
	.B1(U_addrdec_n254), 
	.A2(debug_ad_col_addr_15_), 
	.A1(U_addrdec_n28));
   NAND3_X2 U_addrdec_U217 (.ZN(debug_ad_row_addr[5]), 
	.A3(U_addrdec_n168), 
	.A2(U_addrdec_n169), 
	.A1(U_addrdec_n170));
   AOI22_X2 U_addrdec_U216 (.ZN(U_addrdec_n277), 
	.B2(U_addrdec_n18), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n265), 
	.A1(U_addrdec_n28));
   AOI22_X2 U_addrdec_U215 (.ZN(U_addrdec_n276), 
	.B2(U_addrdec_n37), 
	.B1(U_addrdec_n266), 
	.A2(U_addrdec_n267), 
	.A1(U_addrdec_n38));
   NAND2_X2 U_addrdec_U214 (.ZN(U_addrdec_n255), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[31]));
   AOI22_X2 U_addrdec_U213 (.ZN(U_addrdec_n275), 
	.B2(U_addrdec_n26), 
	.B1(U_addrdec_n268), 
	.A2(U_addrdec_n269), 
	.A1(U_addrdec_n270));
   AOI22_X2 U_addrdec_U212 (.ZN(U_addrdec_n274), 
	.B2(U_addrdec_n17), 
	.B1(U_addrdec_n271), 
	.A2(U_addrdec_n272), 
	.A1(U_addrdec_n273));
   NAND4_X2 U_addrdec_U211 (.ZN(U_addrdec_n278), 
	.A4(U_addrdec_n274), 
	.A3(U_addrdec_n275), 
	.A2(U_addrdec_n276), 
	.A1(U_addrdec_n277));
   NOR2_X2 U_addrdec_U210 (.ZN(U_addrdec_n248), 
	.A2(U_addrdec_n25), 
	.A1(U_addrdec_n255));
   OAI22_X2 U_addrdec_U209 (.ZN(U_addrdec_n247), 
	.B2(U_addrdec_n243), 
	.B1(U_addrdec_n244), 
	.A2(U_addrdec_n245), 
	.A1(U_addrdec_n246));
   AOI211_X2 U_addrdec_U208 (.ZN(U_addrdec_n252), 
	.C2(U_addrdec_n270), 
	.C1(U_addrdec_n35), 
	.B(U_addrdec_n247), 
	.A(U_addrdec_n248));
   AOI22_X2 U_addrdec_U207 (.ZN(U_addrdec_n251), 
	.B2(U_addrdec_n37), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n266), 
	.A1(U_addrdec_n272));
   AOI22_X2 U_addrdec_U206 (.ZN(U_addrdec_n250), 
	.B2(U_addrdec_n269), 
	.B1(U_addrdec_n273), 
	.A2(U_addrdec_n265), 
	.A1(U_addrdec_n38));
   AOI22_X2 U_addrdec_U205 (.ZN(U_addrdec_n249), 
	.B2(U_addrdec_n26), 
	.B1(U_addrdec_n271), 
	.A2(U_addrdec_n17), 
	.A1(U_addrdec_n267));
   NAND4_X2 U_addrdec_U204 (.ZN(U_addrdec_n253), 
	.A4(U_addrdec_n249), 
	.A3(U_addrdec_n250), 
	.A2(U_addrdec_n251), 
	.A1(U_addrdec_n252));
   OAI22_X2 U_addrdec_U203 (.ZN(U_addrdec_n185), 
	.B2(U_addrdec_n243), 
	.B1(U_addrdec_n13), 
	.A2(U_addrdec_n245), 
	.A1(U_addrdec_n180));
   AOI22_X2 U_addrdec_U202 (.ZN(U_addrdec_n183), 
	.B2(FE_OFN353_U_addrdec_n272), 
	.B1(U_addrdec_n219), 
	.A2(U_addrdec_n181), 
	.A1(U_addrdec_n38));
   AOI22_X2 U_addrdec_U201 (.ZN(U_addrdec_n182), 
	.B2(U_addrdec_n37), 
	.B1(U_addrdec_n34), 
	.A2(U_addrdec_n232), 
	.A1(U_addrdec_n17));
   NAND2_X2 U_addrdec_U200 (.ZN(U_addrdec_n184), 
	.A2(U_addrdec_n182), 
	.A1(U_addrdec_n183));
   AOI211_X2 U_addrdec_U199 (.ZN(U_addrdec_n190), 
	.C2(U_addrdec_n265), 
	.C1(U_addrdec_n36), 
	.B(U_addrdec_n184), 
	.A(U_addrdec_n185));
   AOI22_X2 U_addrdec_U198 (.ZN(U_addrdec_n189), 
	.B2(U_addrdec_n269), 
	.B1(U_addrdec_n242), 
	.A2(U_addrdec_n254), 
	.A1(U_addrdec_n26));
   AOI22_X2 U_addrdec_U197 (.ZN(U_addrdec_n188), 
	.B2(U_addrdec_n35), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n266), 
	.A1(U_addrdec_n30));
   NAND3_X2 U_addrdec_U196 (.ZN(debug_ad_row_addr[7]), 
	.A3(U_addrdec_n188), 
	.A2(U_addrdec_n189), 
	.A1(U_addrdec_n190));
   AOI22_X2 U_addrdec_U195 (.ZN(U_addrdec_n236), 
	.B2(U_addrdec_n18), 
	.B1(U_addrdec_n232), 
	.A2(U_addrdec_n242), 
	.A1(U_addrdec_n28));
   AOI22_X2 U_addrdec_U194 (.ZN(U_addrdec_n235), 
	.B2(U_addrdec_n272), 
	.B1(U_addrdec_n265), 
	.A2(U_addrdec_n254), 
	.A1(U_addrdec_n37));
   AOI22_X2 U_addrdec_U193 (.ZN(U_addrdec_n234), 
	.B2(U_addrdec_n30), 
	.B1(U_addrdec_n268), 
	.A2(U_addrdec_n36), 
	.A1(U_addrdec_n270));
   NAND4_X2 U_addrdec_U192 (.ZN(U_addrdec_n240), 
	.A4(U_addrdec_n233), 
	.A3(U_addrdec_n234), 
	.A2(U_addrdec_n235), 
	.A1(U_addrdec_n236));
   AOI22_X2 U_addrdec_U191 (.ZN(U_addrdec_n238), 
	.B2(U_addrdec_n38), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n266), 
	.A1(U_addrdec_n17));
   AOI22_X2 U_addrdec_U190 (.ZN(U_addrdec_n237), 
	.B2(U_addrdec_n269), 
	.B1(U_addrdec_n267), 
	.A2(U_addrdec_n273), 
	.A1(U_addrdec_n26));
   NAND2_X2 U_addrdec_U189 (.ZN(U_addrdec_n239), 
	.A2(U_addrdec_n237), 
	.A1(U_addrdec_n238));
   OAI21_X2 U_addrdec_U188 (.ZN(U_addrdec_n241), 
	.B2(U_addrdec_n239), 
	.B1(U_addrdec_n240), 
	.A(U_addrdec_row_addr_mask[12]));
   INV_X4 U_addrdec_U187 (.ZN(debug_ad_row_addr[12]), 
	.A(U_addrdec_n241));
   OAI22_X2 U_addrdec_U186 (.ZN(U_addrdec_n145), 
	.B2(U_addrdec_n161), 
	.B1(U_addrdec_n13), 
	.A2(U_addrdec_n150), 
	.A1(U_addrdec_n180));
   AOI22_X2 U_addrdec_U185 (.ZN(U_addrdec_n143), 
	.B2(U_addrdec_n269), 
	.B1(U_addrdec_n34), 
	.A2(U_addrdec_n181), 
	.A1(U_addrdec_n26));
   AOI22_X2 U_addrdec_U184 (.ZN(U_addrdec_n142), 
	.B2(U_addrdec_n30), 
	.B1(U_addrdec_n242), 
	.A2(U_addrdec_n219), 
	.A1(U_addrdec_n35));
   NAND2_X2 U_addrdec_U183 (.ZN(U_addrdec_n144), 
	.A2(U_addrdec_n142), 
	.A1(U_addrdec_n143));
   AOI211_X2 U_addrdec_U182 (.ZN(U_addrdec_n149), 
	.C2(debug_ad_col_addr_15_), 
	.C1(U_addrdec_n38), 
	.B(U_addrdec_n144), 
	.A(U_addrdec_n145));
   AOI22_X2 U_addrdec_U181 (.ZN(U_addrdec_n148), 
	.B2(U_addrdec_n36), 
	.B1(U_addrdec_n232), 
	.A2(U_addrdec_n28), 
	.A1(debug_ad_col_addr_13__BAR_BAR));
   AOI22_X2 U_addrdec_U180 (.ZN(U_addrdec_n147), 
	.B2(U_addrdec_n37), 
	.B1(debug_ad_col_addr_14_), 
	.A2(U_addrdec_n18), 
	.A1(debug_ad_col_addr_12__BAR_BAR));
   NAND3_X2 U_addrdec_U179 (.ZN(debug_ad_row_addr[3]), 
	.A3(U_addrdec_n147), 
	.A2(U_addrdec_n148), 
	.A1(U_addrdec_n149));
   OAI22_X2 U_addrdec_U178 (.ZN(U_addrdec_n174), 
	.B2(U_addrdec_n23), 
	.B1(U_addrdec_n13), 
	.A2(U_addrdec_n243), 
	.A1(U_addrdec_n180));
   AOI22_X2 U_addrdec_U177 (.ZN(U_addrdec_n172), 
	.B2(FE_OFN353_U_addrdec_n272), 
	.B1(U_addrdec_n181), 
	.A2(U_addrdec_n34), 
	.A1(U_addrdec_n38));
   AOI22_X2 U_addrdec_U176 (.ZN(U_addrdec_n171), 
	.B2(U_addrdec_n26), 
	.B1(U_addrdec_n242), 
	.A2(U_addrdec_n219), 
	.A1(U_addrdec_n17));
   NAND2_X2 U_addrdec_U175 (.ZN(U_addrdec_n173), 
	.A2(U_addrdec_n171), 
	.A1(U_addrdec_n172));
   AOI211_X2 U_addrdec_U174 (.ZN(U_addrdec_n179), 
	.C2(debug_ad_col_addr_15_), 
	.C1(U_addrdec_n18), 
	.B(U_addrdec_n173), 
	.A(U_addrdec_n174));
   AOI22_X2 U_addrdec_U173 (.ZN(U_addrdec_n178), 
	.B2(U_addrdec_n35), 
	.B1(U_addrdec_n254), 
	.A2(U_addrdec_n232), 
	.A1(U_addrdec_n269));
   AOI22_X2 U_addrdec_U172 (.ZN(U_addrdec_n177), 
	.B2(U_addrdec_n36), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n265), 
	.A1(U_addrdec_n30));
   NAND3_X2 U_addrdec_U171 (.ZN(debug_ad_row_addr[6]), 
	.A3(U_addrdec_n177), 
	.A2(U_addrdec_n178), 
	.A1(U_addrdec_n179));
   OAI22_X2 U_addrdec_U170 (.ZN(U_addrdec_n194), 
	.B2(U_addrdec_n245), 
	.B1(U_addrdec_n13), 
	.A2(U_addrdec_n23), 
	.A1(U_addrdec_n210));
   AOI22_X2 U_addrdec_U169 (.ZN(U_addrdec_n192), 
	.B2(U_addrdec_n272), 
	.B1(U_addrdec_n232), 
	.A2(U_addrdec_n34), 
	.A1(U_addrdec_n28));
   AOI22_X2 U_addrdec_U168 (.ZN(U_addrdec_n191), 
	.B2(U_addrdec_n17), 
	.B1(U_addrdec_n242), 
	.A2(U_addrdec_n219), 
	.A1(U_addrdec_n38));
   NAND2_X2 U_addrdec_U167 (.ZN(U_addrdec_n193), 
	.A2(U_addrdec_n191), 
	.A1(U_addrdec_n192));
   AOI211_X2 U_addrdec_U166 (.ZN(U_addrdec_n199), 
	.C2(U_addrdec_n266), 
	.C1(U_addrdec_n36), 
	.B(U_addrdec_n193), 
	.A(U_addrdec_n194));
   AOI22_X2 U_addrdec_U165 (.ZN(U_addrdec_n198), 
	.B2(U_addrdec_n26), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n254), 
	.A1(U_addrdec_n269));
   AOI22_X2 U_addrdec_U164 (.ZN(U_addrdec_n197), 
	.B2(U_addrdec_n30), 
	.B1(U_addrdec_n267), 
	.A2(U_addrdec_n265), 
	.A1(U_addrdec_n35));
   NAND3_X2 U_addrdec_U163 (.ZN(debug_ad_row_addr[8]), 
	.A3(U_addrdec_n197), 
	.A2(U_addrdec_n198), 
	.A1(U_addrdec_n199));
   OAI22_X2 U_addrdec_U162 (.ZN(U_addrdec_n154), 
	.B2(U_addrdec_n150), 
	.B1(U_addrdec_n13), 
	.A2(U_addrdec_n22), 
	.A1(U_addrdec_n180));
   AOI22_X2 U_addrdec_U161 (.ZN(U_addrdec_n152), 
	.B2(U_addrdec_n269), 
	.B1(U_addrdec_n181), 
	.A2(U_addrdec_n219), 
	.A1(U_addrdec_n26));
   AOI22_X2 U_addrdec_U160 (.ZN(U_addrdec_n151), 
	.B2(U_addrdec_n35), 
	.B1(U_addrdec_n232), 
	.A2(U_addrdec_n34), 
	.A1(U_addrdec_n17));
   NAND2_X2 U_addrdec_U159 (.ZN(U_addrdec_n153), 
	.A2(U_addrdec_n151), 
	.A1(U_addrdec_n152));
   AOI211_X2 U_addrdec_U158 (.ZN(U_addrdec_n160), 
	.C2(debug_ad_col_addr_15_), 
	.C1(U_addrdec_n37), 
	.B(U_addrdec_n153), 
	.A(U_addrdec_n154));
   AOI22_X2 U_addrdec_U157 (.ZN(U_addrdec_n159), 
	.B2(U_addrdec_n36), 
	.B1(U_addrdec_n242), 
	.A2(U_addrdec_n254), 
	.A1(U_addrdec_n30));
   AOI22_X2 U_addrdec_U156 (.ZN(U_addrdec_n158), 
	.B2(U_addrdec_n28), 
	.B1(debug_ad_col_addr_14_), 
	.A2(U_addrdec_n18), 
	.A1(debug_ad_col_addr_13__BAR_BAR));
   NAND3_X2 U_addrdec_U155 (.ZN(debug_ad_row_addr[4]), 
	.A3(U_addrdec_n158), 
	.A2(U_addrdec_n159), 
	.A1(U_addrdec_n160));
   OAI22_X2 U_addrdec_U154 (.ZN(U_addrdec_n112), 
	.B2(U_addrdec_n24), 
	.B1(U_addrdec_n13), 
	.A2(U_addrdec_n256), 
	.A1(U_addrdec_n180));
   AOI22_X2 U_addrdec_U153 (.ZN(U_addrdec_n109), 
	.B2(U_addrdec_n36), 
	.B1(U_addrdec_n34), 
	.A2(U_addrdec_n181), 
	.A1(U_addrdec_n30));
   NAND2_X2 U_addrdec_U152 (.ZN(U_addrdec_n111), 
	.A2(U_addrdec_n109), 
	.A1(U_addrdec_n110));
   AOI211_X2 U_addrdec_U151 (.ZN(U_addrdec_n120), 
	.C2(debug_ad_col_addr_13__BAR_BAR), 
	.C1(U_addrdec_n272), 
	.B(U_addrdec_n111), 
	.A(U_addrdec_n112));
   AOI22_X2 U_addrdec_U150 (.ZN(U_addrdec_n119), 
	.B2(U_addrdec_n269), 
	.B1(debug_ad_col_addr_15_), 
	.A2(debug_ad_col_addr_11_), 
	.A1(U_addrdec_n37));
   AOI22_X2 U_addrdec_U149 (.ZN(U_addrdec_n118), 
	.B2(U_addrdec_n17), 
	.B1(debug_ad_col_addr_14_), 
	.A2(U_addrdec_n38), 
	.A1(debug_ad_col_addr_12__BAR_BAR));
   NAND3_X2 U_addrdec_U148 (.ZN(debug_ad_row_addr[0]), 
	.A3(U_addrdec_n118), 
	.A2(U_addrdec_n119), 
	.A1(U_addrdec_n120));
   INV_X4 U_addrdec_U147 (.ZN(U_addrdec_n211), 
	.A(U_addrdec_n219));
   OAI22_X2 U_addrdec_U146 (.ZN(U_addrdec_n215), 
	.B2(U_addrdec_n245), 
	.B1(U_addrdec_n210), 
	.A2(U_addrdec_n243), 
	.A1(U_addrdec_n211));
   AOI22_X2 U_addrdec_U145 (.ZN(U_addrdec_n213), 
	.B2(U_addrdec_n37), 
	.B1(U_addrdec_n232), 
	.A2(U_addrdec_n254), 
	.A1(U_addrdec_n272));
   AOI22_X2 U_addrdec_U144 (.ZN(U_addrdec_n212), 
	.B2(U_addrdec_n17), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n242), 
	.A1(U_addrdec_n38));
   NAND2_X2 U_addrdec_U143 (.ZN(U_addrdec_n214), 
	.A2(U_addrdec_n212), 
	.A1(U_addrdec_n213));
   AOI211_X2 U_addrdec_U142 (.ZN(U_addrdec_n218), 
	.C2(U_addrdec_n273), 
	.C1(U_addrdec_n36), 
	.B(U_addrdec_n214), 
	.A(U_addrdec_n215));
   AOI22_X2 U_addrdec_U141 (.ZN(U_addrdec_n217), 
	.B2(U_addrdec_n26), 
	.B1(U_addrdec_n266), 
	.A2(U_addrdec_n265), 
	.A1(U_addrdec_n269));
   AOI22_X2 U_addrdec_U140 (.ZN(U_addrdec_n216), 
	.B2(U_addrdec_n30), 
	.B1(U_addrdec_n271), 
	.A2(U_addrdec_n35), 
	.A1(U_addrdec_n267));
   NAND3_X2 U_addrdec_U139 (.ZN(debug_ad_row_addr[10]), 
	.A3(U_addrdec_n216), 
	.A2(U_addrdec_n217), 
	.A1(U_addrdec_n218));
   AOI22_X2 U_addrdec_U138 (.ZN(U_addrdec_n262), 
	.B2(U_addrdec_n28), 
	.B1(U_addrdec_n264), 
	.A2(U_addrdec_n254), 
	.A1(U_addrdec_n18));
   OAI22_X2 U_addrdec_U137 (.ZN(U_addrdec_n258), 
	.B2(U_addrdec_n24), 
	.B1(U_addrdec_n255), 
	.A2(U_addrdec_n256), 
	.A1(U_addrdec_n257));
   AOI21_X2 U_addrdec_U136 (.ZN(U_addrdec_n261), 
	.B2(U_addrdec_n271), 
	.B1(U_addrdec_n269), 
	.A(U_addrdec_n258));
   AOI22_X2 U_addrdec_U135 (.ZN(U_addrdec_n260), 
	.B2(U_addrdec_n37), 
	.B1(U_addrdec_n265), 
	.A2(U_addrdec_n266), 
	.A1(U_addrdec_n38));
   AOI22_X2 U_addrdec_U134 (.ZN(U_addrdec_n259), 
	.B2(U_addrdec_n272), 
	.B1(U_addrdec_n267), 
	.A2(U_addrdec_n273), 
	.A1(U_addrdec_n17));
   NAND4_X2 U_addrdec_U133 (.ZN(U_addrdec_n263), 
	.A4(U_addrdec_n259), 
	.A3(U_addrdec_n260), 
	.A2(U_addrdec_n261), 
	.A1(U_addrdec_n262));
   NOR3_X2 U_addrdec_U132 (.ZN(U_addrdec_n311), 
	.A3(U_addrdec_sram_select_0_), 
	.A2(U_addrdec_rom_select_0_), 
	.A1(U_addrdec_flash_select_0_));
   NOR3_X2 U_addrdec_U131 (.ZN(ad_static_mem_req), 
	.A3(U_addrdec_n310), 
	.A2(ad_sdram_type_0_), 
	.A1(U_addrdec_n311));
   AOI22_X2 U_addrdec_U130 (.ZN(U_addrdec_n295), 
	.B2(U_addrdec_n293), 
	.B1(hiu_haddr[1]), 
	.A2(hiu_hsize[0]), 
	.A1(hiu_haddr[0]));
   NOR2_X2 U_addrdec_U129 (.ZN(U_addrdec_n300), 
	.A2(hiu_hsize[0]), 
	.A1(hiu_haddr[0]));
   AOI22_X2 U_addrdec_U128 (.ZN(U_addrdec_n294), 
	.B2(U_addrdec_n40), 
	.B1(U_addrdec_n296), 
	.A2(U_addrdec_n295), 
	.A1(big_endian));
   NAND2_X2 U_addrdec_U127 (.ZN(U_addrdec_n297), 
	.A2(hiu_haddr[0]), 
	.A1(hiu_haddr[1]));
   AOI21_X2 U_addrdec_U126 (.ZN(ad_cr_data_mask[1]), 
	.B2(U_addrdec_n297), 
	.B1(U_addrdec_n294), 
	.A(U_addrdec_n301));
   AOI22_X2 U_addrdec_U125 (.ZN(U_addrdec_n299), 
	.B2(U_addrdec_n40), 
	.B1(U_addrdec_n291), 
	.A2(hiu_haddr[1]), 
	.A1(big_endian));
   AOI221_X2 U_addrdec_U124 (.ZN(U_addrdec_n302), 
	.C2(U_addrdec_n40), 
	.C1(U_addrdec_n300), 
	.B2(big_endian), 
	.B1(hiu_haddr[0]), 
	.A(U_addrdec_n303));
   NOR2_X2 U_addrdec_U123 (.ZN(ad_cr_data_mask[3]), 
	.A2(U_addrdec_n301), 
	.A1(U_addrdec_n302));
   AOI221_X2 U_addrdec_U122 (.ZN(U_addrdec_n292), 
	.C2(U_addrdec_n40), 
	.C1(hiu_haddr[0]), 
	.B2(big_endian), 
	.B1(U_addrdec_n300), 
	.A(U_addrdec_n299));
   NOR2_X2 U_addrdec_U121 (.ZN(ad_cr_data_mask[0]), 
	.A2(U_addrdec_n301), 
	.A1(U_addrdec_n292));
   AOI22_X2 U_addrdec_U120 (.ZN(U_addrdec_n298), 
	.B2(U_addrdec_n40), 
	.B1(U_addrdec_n295), 
	.A2(U_addrdec_n296), 
	.A1(big_endian));
   AOI21_X2 U_addrdec_U119 (.ZN(ad_cr_data_mask[2]), 
	.B2(U_addrdec_n297), 
	.B1(U_addrdec_n298), 
	.A(U_addrdec_n301));
   INV_X4 U_addrdec_U118 (.ZN(debug_ad_col_addr_1_), 
	.A(U_addrdec_n96));
   INV_X4 U_addrdec_U117 (.ZN(debug_ad_col_addr_4_), 
	.A(U_addrdec_n97));
   INV_X4 U_addrdec_U116 (.ZN(debug_ad_col_addr_6_), 
	.A(U_addrdec_n99));
   INV_X4 U_addrdec_U115 (.ZN(debug_ad_col_addr_5_), 
	.A(U_addrdec_n98));
   INV_X4 U_addrdec_U114 (.ZN(debug_ad_col_addr_7_), 
	.A(U_addrdec_n100));
   NAND2_X2 U_addrdec_U113 (.ZN(U_addrdec_n283), 
	.A2(U_addrdec_n281), 
	.A1(U_addrdec_n282));
   NAND2_X2 U_addrdec_U112 (.ZN(U_addrdec_n286), 
	.A2(U_addrdec_n280), 
	.A1(U_addrdec_n281));
   OAI221_X2 U_addrdec_U111 (.ZN(U_addrdec_N133), 
	.C2(U_cr_n21), 
	.C1(U_addrdec_n290), 
	.B2(cr_row_addr_width[1]), 
	.B1(FE_PHN3054_cr_row_addr_width_2_), 
	.A(FE_PHN1064_cr_row_addr_width_3_));
   NOR3_X2 U_addrdec_U110 (.ZN(U_addrdec_n347), 
	.A3(FE_PHN3126_cr_block_size1_6_), 
	.A2(cr_block_size1[5]), 
	.A1(FE_PHN1855_cr_block_size1_7_));
   NAND2_X2 U_addrdec_U109 (.ZN(U_addrdec_n309), 
	.A2(FE_PHN1634_U_cr_n167), 
	.A1(cr_block_size1[5]));
   NOR2_X2 U_addrdec_U108 (.ZN(U_addrdec_n348), 
	.A2(FE_PHN1868_U_addrdec_n309), 
	.A1(FE_PHN3126_cr_block_size1_6_));
   NOR3_X2 U_addrdec_U107 (.ZN(U_addrdec_n346), 
	.A3(FE_PHN1642_U_cr_n119), 
	.A2(cr_block_size1[5]), 
	.A1(FE_PHN1855_cr_block_size1_7_));
   NOR2_X2 U_addrdec_U106 (.ZN(U_addrdec_n345), 
	.A2(FE_PHN1642_U_cr_n119), 
	.A1(FE_PHN1868_U_addrdec_n309));
   NOR2_X2 U_addrdec_U105 (.ZN(U_addrdec_n269), 
	.A2(U_addrdec_n116), 
	.A1(U_addrdec_n114));
   NAND2_X2 U_addrdec_U104 (.ZN(debug_ad_col_addr_11_), 
	.A2(U_addrdec_n53), 
	.A1(U_addrdec_n54));
   NOR2_X1 U_addrdec_U103 (.ZN(debug_ad_col_addr_0_), 
	.A2(U_addrdec_n95), 
	.A1(U_addrdec_n39));
   NAND2_X2 U_addrdec_U101 (.ZN(U_addrdec_n53), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[11]));
   AOI22_X2 U_addrdec_U98 (.ZN(U_addrdec_n110), 
	.B2(U_addrdec_n18), 
	.B1(debug_ad_col_addr_9_), 
	.A2(debug_ad_col_addr_10_), 
	.A1(U_addrdec_n28));
   INV_X1 U_addrdec_U97 (.ZN(debug_ad_col_addr_13__BAR_BAR), 
	.A(debug_ad_col_addr_13_));
   AOI211_X2 U_addrdec_U90 (.ZN(U_addrdec_n170), 
	.C2(debug_ad_col_addr_14_), 
	.C1(U_addrdec_n18), 
	.B(U_addrdec_n164), 
	.A(U_addrdec_n165));
   NAND2_X1 U_addrdec_U89 (.ZN(U_addrdec_n42), 
	.A2(FE_PHN918_cr_bank_addr_width_0_), 
	.A1(n[26]));
   OR2_X2 U_addrdec_U87 (.ZN(U_addrdec_N119), 
	.A2(FE_PHN918_cr_bank_addr_width_0_), 
	.A1(FE_PHN1034_cr_bank_addr_width_1_));
   NAND2_X1 U_addrdec_U84 (.ZN(U_addrdec_n287), 
	.A2(FE_PHN1064_cr_row_addr_width_3_), 
	.A1(FE_PHN3054_cr_row_addr_width_2_));
   NAND2_X1 U_addrdec_U81 (.ZN(U_addrdec_n290), 
	.A2(cr_row_addr_width[1]), 
	.A1(FE_PHN3054_cr_row_addr_width_2_));
   NAND3_X1 U_addrdec_U79 (.ZN(U_addrdec_N130), 
	.A3(FE_PHN1254_U_cr_n55), 
	.A2(FE_PHN1064_cr_row_addr_width_3_), 
	.A1(cr_row_addr_width[1]));
   NAND2_X1 U_addrdec_U77 (.ZN(U_addrdec_n280), 
	.A2(U_cr_n22), 
	.A1(U_addrdec_n42));
   INV_X2 U_addrdec_U76 (.ZN(U_addrdec_n101), 
	.A(U_addrdec_n106));
   OAI21_X1 U_addrdec_U75 (.ZN(U_addrdec_n58), 
	.B2(U_addrdec_n287), 
	.B1(cr_row_addr_width[1]), 
	.A(U_addrdec_N130));
   OR2_X2 U_addrdec_U74 (.ZN(U_addrdec_N129), 
	.A2(cr_row_addr_width[0]), 
	.A1(U_addrdec_N130));
   NAND2_X1 U_addrdec_U73 (.ZN(U_addrdec_n281), 
	.A2(n[25]), 
	.A1(U_addrdec_n41));
   INV_X1 U_addrdec_U72 (.ZN(U_addrdec_n56), 
	.A(U_addrdec_n81));
   NAND2_X1 U_addrdec_U71 (.ZN(U_addrdec_n205), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[28]));
   NAND2_X1 U_addrdec_U70 (.ZN(U_addrdec_n206), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[29]));
   NAND2_X1 U_addrdec_U69 (.ZN(U_addrdec_n196), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[28]));
   OAI21_X1 U_addrdec_U68 (.ZN(U_addrdec_N131), 
	.B2(FE_PHN1254_U_cr_n55), 
	.B1(U_cr_n21), 
	.A(FE_PHN1662_U_addrdec_n58));
   INV_X2 U_addrdec_U67 (.ZN(U_addrdec_n95), 
	.A(hiu_addr[1]));
   NAND2_X1 U_addrdec_U66 (.ZN(U_addrdec_n285), 
	.A2(n[24]), 
	.A1(U_addrdec_n283));
   INV_X1 U_addrdec_U65 (.ZN(U_addrdec_n293), 
	.A(hiu_haddr[0]));
   NAND2_X1 U_addrdec_U64 (.ZN(U_addrdec_n104), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[18]));
   NAND2_X1 U_addrdec_U63 (.ZN(U_addrdec_n103), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[17]));
   NAND2_X1 U_addrdec_U62 (.ZN(U_addrdec_n108), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[19]));
   INV_X2 U_addrdec_U59 (.ZN(U_addrdec_n268), 
	.A(U_addrdec_n255));
   INV_X2 U_addrdec_U58 (.ZN(U_addrdec_n150), 
	.A(U_addrdec_n272));
   INV_X2 U_addrdec_U57 (.ZN(U_addrdec_n130), 
	.A(U_addrdec_n269));
   INV_X2 U_addrdec_U56 (.ZN(U_addrdec_n244), 
	.A(U_addrdec_n254));
   INV_X2 U_addrdec_U55 (.ZN(U_addrdec_n246), 
	.A(U_addrdec_n242));
   NAND2_X1 U_addrdec_U54 (.ZN(U_addrdec_n233), 
	.A2(U_addrdec_n35), 
	.A1(U_addrdec_n271));
   NAND2_X1 U_addrdec_U53 (.ZN(U_addrdec_n223), 
	.A2(U_addrdec_n36), 
	.A1(U_addrdec_n271));
   NOR2_X2 U_addrdec_U49 (.ZN(debug_ad_col_addr_12_), 
	.A2(U_addrdec_n27), 
	.A1(U_addrdec_n32));
   INV_X2 U_addrdec_U48 (.ZN(U_addrdec_n257), 
	.A(U_addrdec_n270));
   OR2_X2 U_addrdec_U47 (.ZN(U_addrdec_n296), 
	.A2(U_addrdec_n300), 
	.A1(hiu_haddr[1]));
   OAI21_X1 U_addrdec_U46 (.ZN(U_addrdec_n284), 
	.B2(U_addrdec_n283), 
	.B1(n[24]), 
	.A(U_addrdec_n285));
   XOR2_X1 U_addrdec_U45 (.Z(U_addrdec_N110), 
	.B(FE_PHN1645_U_cr_n65), 
	.A(U_addrdec_n285));
   NOR2_X1 U_addrdec_U44 (.ZN(U_addrdec_N111), 
	.A2(FE_PHN1645_U_cr_n65), 
	.A1(U_addrdec_n285));
   INV_X2 U_addrdec_U43 (.ZN(U_addrdec_n62), 
	.A(debug_ad_col_addr_10_));
   INV_X2 U_addrdec_U42 (.ZN(U_addrdec_n61), 
	.A(debug_ad_col_addr_9_));
   INV_X2 U_addrdec_U41 (.ZN(U_addrdec_n200), 
	.A(U_addrdec_n34));
   NAND2_X1 U_addrdec_U40 (.ZN(U_addrdec_n162), 
	.A2(FE_OFN353_U_addrdec_n272), 
	.A1(U_addrdec_n34));
   INV_X2 U_addrdec_U39 (.ZN(U_addrdec_n303), 
	.A(U_addrdec_n299));
   INV_X2 U_addrdec_U38 (.ZN(U_addrdec_N109), 
	.A(U_addrdec_n284));
   INV_X1 U_addrdec_U37 (.ZN(U_addrdec_n59), 
	.A(U_addrdec_n88));
   NOR2_X2 U_addrdec_U36 (.ZN(sdram_req_i), 
	.A2(U_addrdec_n310), 
	.A1(ad_sdram_chip_select_0_));
   INV_X2 U_addrdec_U33 (.ZN(U_addrdec_n91), 
	.A(U_addrdec_n86));
   INV_X1 U_addrdec_U32 (.ZN(U_addrdec_n41), 
	.A(U_addrdec_n42));
   NAND2_X2 U_addrdec_U31 (.ZN(U_addrdec_n282), 
	.A2(FE_PHN1034_cr_bank_addr_width_1_), 
	.A1(U_addrdec_n280));
   INV_X2 U_addrdec_U30 (.ZN(U_addrdec_n256), 
	.A(U_addrdec_n26));
   NAND2_X1 U_addrdec_U29 (.ZN(U_addrdec_n221), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[31]));
   NAND2_X1 U_addrdec_U28 (.ZN(U_addrdec_n222), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[30]));
   NAND2_X1 U_addrdec_U27 (.ZN(U_addrdec_n175), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[26]));
   NAND2_X1 U_addrdec_U26 (.ZN(U_addrdec_n195), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[27]));
   NAND2_X1 U_addrdec_U25 (.ZN(U_addrdec_n187), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[27]));
   NAND2_X1 U_addrdec_U24 (.ZN(U_addrdec_n186), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[26]));
   INV_X2 U_addrdec_U23 (.ZN(U_addrdec_n291), 
	.A(hiu_haddr[1]));
   XNOR2_X1 U_addrdec_U21 (.ZN(U_addrdec_N107), 
	.B(FE_PHN918_cr_bank_addr_width_0_), 
	.A(FE_PHN3113_U_cr_n63));
   INV_X1 U_addrdec_U20 (.ZN(U_addrdec_n271), 
	.A(U_addrdec_n11));
   AOI22_X1 U_addrdec_U19 (.ZN(U_addrdec_n11), 
	.B2(hiu_addr[29]), 
	.B1(U_addrdec_n39), 
	.A2(hiu_addr[30]), 
	.A1(U_addrdec_n220));
   INV_X1 U_addrdec_U18 (.ZN(U_addrdec_n34), 
	.A(U_addrdec_n10));
   AOI22_X1 U_addrdec_U17 (.ZN(U_addrdec_n10), 
	.B2(hiu_addr[19]), 
	.B1(U_addrdec_n220), 
	.A2(hiu_addr[18]), 
	.A1(U_addrdec_n39));
   INV_X1 U_addrdec_U16 (.ZN(debug_ad_col_addr_3_), 
	.A(U_addrdec_n9));
   AOI22_X1 U_addrdec_U15 (.ZN(U_addrdec_n9), 
	.B2(U_addrdec_n39), 
	.B1(hiu_addr[3]), 
	.A2(U_addrdec_n220), 
	.A1(hiu_addr[4]));
   AOI22_X2 U_addrdec_U14 (.ZN(U_addrdec_n30), 
	.B2(U_addrdec_n7), 
	.B1(U_addrdec_n5), 
	.A2(U_addrdec_n15), 
	.A1(U_addrdec_bcawp_3_));
   AOI22_X2 U_addrdec_U13 (.ZN(U_addrdec_n7), 
	.B2(U_addrdec_n21), 
	.B1(U_addrdec_bcawp_0_), 
	.A2(U_addrdec_n20), 
	.A1(U_addrdec_n15));
   AOI221_X2 U_addrdec_U12 (.ZN(U_addrdec_n5), 
	.C2(U_addrdec_bcawp_4_), 
	.C1(U_addrdec_bcawp_2_), 
	.B2(U_addrdec_bcawp_4_), 
	.B1(U_addrdec_bcawp_3_), 
	.A(U_addrdec_n4));
   INV_X4 U_addrdec_U11 (.ZN(U_addrdec_n4), 
	.A(U_addrdec_n115));
   NAND4_X1 U_addrdec_U10 (.ZN(U_addrdec_n25), 
	.A4(U_addrdec_n3), 
	.A3(U_addrdec_n20), 
	.A2(U_addrdec_bcawp_4_), 
	.A1(U_addrdec_n14));
   INV_X1 U_addrdec_U9 (.ZN(U_addrdec_n3), 
	.A(U_addrdec_n113));
   OR2_X1 U_addrdec_U8 (.ZN(U_addrdec_n301), 
	.A2(hiu_hsize[1]), 
	.A1(hiu_hsize[2]));
   INV_X1 U_addrdec_U7 (.ZN(debug_ad_col_addr_2_), 
	.A(U_addrdec_n2));
   AOI22_X1 U_addrdec_U6 (.ZN(U_addrdec_n2), 
	.B2(U_addrdec_n220), 
	.B1(hiu_addr[3]), 
	.A2(U_addrdec_n39), 
	.A1(hiu_addr[2]));
   INV_X1 U_addrdec_U5 (.ZN(U_addrdec_n102), 
	.A(U_addrdec_n1));
   AOI22_X2 U_addrdec_U4 (.ZN(U_addrdec_n1), 
	.B2(hiu_addr[16]), 
	.B1(U_addrdec_n39), 
	.A2(hiu_addr[17]), 
	.A1(U_addrdec_n220));
   NAND2_X2 U_addrdec_U3 (.ZN(U_addrdec_n219), 
	.A2(U_addrdec_n121), 
	.A1(U_addrdec_n122));
   DFFR_X2 U_addrdec_bcawp_reg_3_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_addrdec_n14), 
	.Q(U_addrdec_bcawp_3_), 
	.D(U_addrdec_N110), 
	.CK(HCLK__L5_N34));
   DFFR_X2 U_addrdec_bcawp_reg_2_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_addrdec_n16), 
	.Q(U_addrdec_bcawp_2_), 
	.D(U_addrdec_N109), 
	.CK(HCLK__L5_N34));
   DFFR_X2 U_addrdec_bcawp_reg_1_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_addrdec_n21), 
	.Q(U_addrdec_bcawp_1_), 
	.D(FE_PHN927_U_addrdec_N108), 
	.CK(HCLK__L5_N34));
   DFFR_X2 U_addrdec_bcawp_reg_4_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_addrdec_n15), 
	.Q(U_addrdec_bcawp_4_), 
	.D(U_addrdec_N111), 
	.CK(HCLK__L5_N34));
   DFFR_X2 U_addrdec_bcawp_reg_0_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_addrdec_n20), 
	.Q(U_addrdec_bcawp_0_), 
	.D(FE_PHN2025_U_addrdec_N107), 
	.CK(HCLK__L5_N34));
   DFFR_X2 U_addrdec_sdram_select_reg_0_ (.RN(FE_OFN44_HRESETn), 
	.QN(ad_sdram_chip_select_0_), 
	.Q(ad_sdram_type_0_), 
	.D(FE_PHN3373_U_addrdec_n347), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_addrdec_s_data_width_prog_buf_reg_0_ (.RN(FE_OFN35_HRESETn), 
	.QN(U_addrdec_n39), 
	.Q(U_addrdec_n220), 
	.D(FE_PHN5171_n27), 
	.CK(HCLK__L5_N32));
   DFFR_X2 U_addrdec_sram_select_reg_0_ (.RN(FE_OFN188_HRESETn), 
	.Q(U_addrdec_sram_select_0_), 
	.D(FE_PHN2422_U_addrdec_n348), 
	.CK(HCLK__L5_N28));
   DFFR_X2 U_addrdec_rom_select_reg_0_ (.RN(FE_OFN188_HRESETn), 
	.Q(U_addrdec_rom_select_0_), 
	.D(FE_PHN1641_U_addrdec_n345), 
	.CK(HCLK__L5_N32));
   DFFR_X2 U_addrdec_flash_select_reg_0_ (.RN(FE_OFN188_HRESETn), 
	.Q(U_addrdec_flash_select_0_), 
	.D(FE_PHN1854_U_addrdec_n346), 
	.CK(HCLK__L5_N32));
   DFFS_X2 U_addrdec_row_addr_mask_hi_reg_0_ (.SN(FE_OFN50_HRESETn), 
	.Q(U_addrdec_row_addr_mask[11]), 
	.D(FE_PHN2431_U_addrdec_N129), 
	.CK(HCLK__L5_N33));
   DFFS_X2 U_addrdec_row_addr_mask_hi_reg_1_ (.SN(FE_OFN50_HRESETn), 
	.Q(U_addrdec_row_addr_mask[12]), 
	.D(FE_PHN3164_U_addrdec_N130), 
	.CK(HCLK__L5_N34));
   DFFS_X2 U_addrdec_row_addr_mask_hi_reg_2_ (.SN(FE_OFN50_HRESETn), 
	.Q(U_addrdec_row_addr_mask[13]), 
	.D(FE_PHN2146_U_addrdec_N131), 
	.CK(HCLK__L5_N34));
   DFFR_X1 U_addrdec_row_addr_mask_hi_reg_3_ (.RN(FE_OFN50_HRESETn), 
	.QN(U_addrdec_row_addr_mask[14]), 
	.D(FE_PHN1662_U_addrdec_n58), 
	.CK(HCLK__L5_N34));
   DFFS_X2 U_addrdec_row_addr_mask_hi_reg_4_ (.SN(FE_OFN50_HRESETn), 
	.Q(U_addrdec_row_addr_mask[15]), 
	.D(FE_PHN5102_U_addrdec_N133), 
	.CK(HCLK__L5_N34));
   DFFS_X2 U_addrdec_bank_addr_mask_reg_1_ (.SN(FE_OFN35_HRESETn), 
	.Q(U_addrdec_bank_addr_mask_1_), 
	.D(FE_PHN3188_U_addrdec_N119), 
	.CK(HCLK__L5_N34));
   OAI221_X2 U_refctl_U142 (.ZN(U_refctl_n112), 
	.C2(U_refctl_n97), 
	.C1(U_refctl_current_state_1_), 
	.B2(U_refctl_current_state_0_), 
	.B1(U_refctl_current_state_1_), 
	.A(ctl_auto_ref_en));
   NOR2_X2 U_refctl_U141 (.ZN(U_refctl_count_next_0_), 
	.A2(FE_PHN1663_U_refctl_count_0_), 
	.A1(U_refctl_n112));
   NOR2_X2 U_refctl_U140 (.ZN(U_refctl_n119), 
	.A2(FE_PHN1411_U_refctl_n91), 
	.A1(U_refctl_N27));
   OAI22_X2 U_refctl_U139 (.ZN(U_refctl_n120), 
	.B2(U_refctl_n86), 
	.B1(U_refctl_N28), 
	.A2(U_refctl_n81), 
	.A1(U_refctl_N29));
   AOI22_X2 U_refctl_U138 (.ZN(U_refctl_n115), 
	.B2(FE_PHN1574_U_refctl_n78), 
	.B1(U_refctl_N23), 
	.A2(U_refctl_n87), 
	.A1(U_refctl_N22));
   AOI211_X2 U_refctl_U137 (.ZN(U_refctl_n122), 
	.C2(FE_PHN1424_U_refctl_count_12_), 
	.C1(U_refctl_n121), 
	.B(U_refctl_n119), 
	.A(U_refctl_n120));
   INV_X4 U_refctl_U136 (.ZN(U_refctl_n127), 
	.A(U_refctl_n124));
   AOI221_X2 U_refctl_U135 (.ZN(U_refctl_ref_req_next), 
	.C2(U_refctl_n126), 
	.C1(U_refctl_n92), 
	.B2(U_refctl_n127), 
	.B1(U_refctl_current_state_1_), 
	.A(n94));
   NAND4_X2 U_refctl_U134 (.ZN(U_refctl_n106), 
	.A4(FE_PHN1663_U_refctl_count_0_), 
	.A3(U_refctl_count_1_), 
	.A2(U_refctl_count_2_), 
	.A1(U_refctl_count_3_));
   NOR2_X2 U_refctl_U133 (.ZN(U_refctl_n105), 
	.A2(U_refctl_n106), 
	.A1(U_refctl_n84));
   INV_X4 U_refctl_U132 (.ZN(U_refctl_n107), 
	.A(U_refctl_n105));
   NOR2_X2 U_refctl_U131 (.ZN(U_refctl_n108), 
	.A2(U_refctl_n107), 
	.A1(FE_PHN1548_U_refctl_n85));
   NAND2_X2 U_refctl_U130 (.ZN(U_refctl_n109), 
	.A2(U_refctl_n108), 
	.A1(FE_PHN1419_U_refctl_count_6_));
   NOR2_X2 U_refctl_U129 (.ZN(U_refctl_n110), 
	.A2(U_refctl_n109), 
	.A1(FE_PHN1549_U_refctl_n89));
   NAND2_X2 U_refctl_U128 (.ZN(U_refctl_n113), 
	.A2(U_refctl_n110), 
	.A1(FE_PHN1420_U_refctl_count_8_));
   NOR2_X2 U_refctl_U127 (.ZN(U_refctl_n111), 
	.A2(U_refctl_n113), 
	.A1(FE_PHN1574_U_refctl_n78));
   NAND2_X2 U_refctl_U126 (.ZN(U_refctl_n98), 
	.A2(U_refctl_n111), 
	.A1(FE_PHN1421_U_refctl_count_10_));
   NOR2_X2 U_refctl_U125 (.ZN(U_refctl_n99), 
	.A2(U_refctl_n98), 
	.A1(FE_PHN1583_U_refctl_n80));
   NAND2_X2 U_refctl_U124 (.ZN(U_refctl_n100), 
	.A2(U_refctl_n99), 
	.A1(FE_PHN1424_U_refctl_count_12_));
   NOR2_X2 U_refctl_U123 (.ZN(U_refctl_n101), 
	.A2(U_refctl_n100), 
	.A1(FE_PHN1411_U_refctl_n91));
   AOI211_X2 U_refctl_U122 (.ZN(U_refctl_count_next_13_), 
	.C2(U_refctl_n100), 
	.C1(FE_PHN1411_U_refctl_n91), 
	.B(U_refctl_n101), 
	.A(U_refctl_n112));
   AOI211_X2 U_refctl_U121 (.ZN(U_refctl_count_next_9_), 
	.C2(U_refctl_n113), 
	.C1(FE_PHN1574_U_refctl_n78), 
	.B(U_refctl_n111), 
	.A(U_refctl_n112));
   AOI211_X2 U_refctl_U120 (.ZN(U_refctl_count_next_4_), 
	.C2(U_refctl_n106), 
	.C1(U_refctl_n84), 
	.B(U_refctl_n105), 
	.A(U_refctl_n112));
   AOI211_X2 U_refctl_U119 (.ZN(U_refctl_count_next_11_), 
	.C2(U_refctl_n98), 
	.C1(FE_PHN1583_U_refctl_n80), 
	.B(U_refctl_n99), 
	.A(U_refctl_n112));
   AOI211_X2 U_refctl_U118 (.ZN(U_refctl_count_next_7_), 
	.C2(U_refctl_n109), 
	.C1(FE_PHN1549_U_refctl_n89), 
	.B(U_refctl_n110), 
	.A(U_refctl_n112));
   AOI211_X2 U_refctl_U117 (.ZN(U_refctl_count_next_5_), 
	.C2(U_refctl_n107), 
	.C1(FE_PHN1548_U_refctl_n85), 
	.B(U_refctl_n108), 
	.A(U_refctl_n112));
   INV_X4 U_refctl_U116 (.ZN(U_refctl_n102), 
	.A(U_refctl_n101));
   NOR2_X2 U_refctl_U115 (.ZN(U_refctl_n104), 
	.A2(U_refctl_n102), 
	.A1(FE_PHN1415_U_refctl_n86));
   AOI211_X2 U_refctl_U114 (.ZN(U_refctl_count_next_14_), 
	.C2(U_refctl_n102), 
	.C1(FE_PHN1415_U_refctl_n86), 
	.B(U_refctl_n104), 
	.A(U_refctl_n112));
   AOI21_X2 U_refctl_U113 (.ZN(U_refctl_next_state_0_), 
	.B2(U_refctl_n124), 
	.B1(U_refctl_current_state_1_), 
	.A(U_refctl_n123));
   AOI221_X2 U_refctl_U112 (.ZN(U_refctl_count_next_1_), 
	.C2(U_refctl_n83), 
	.C1(U_refctl_n73), 
	.B2(FE_PHN1663_U_refctl_count_0_), 
	.B1(U_refctl_count_1_), 
	.A(U_refctl_n112));
   AOI221_X2 U_refctl_U111 (.ZN(U_refctl_count_next_15_), 
	.C2(U_refctl_n103), 
	.C1(U_refctl_n81), 
	.B2(U_refctl_n104), 
	.B1(U_refctl_count_15_), 
	.A(U_refctl_n112));
   NOR4_X2 U_refctl_U110 (.ZN(U_refctl_N31), 
	.A4(U_refctl_n64), 
	.A3(U_refctl_n65), 
	.A2(U_refctl_n66), 
	.A1(U_refctl_N30));
   NAND4_X2 U_refctl_U109 (.ZN(U_refctl_n64), 
	.A4(U_refctl_n60), 
	.A3(U_refctl_n61), 
	.A2(U_refctl_n62), 
	.A1(U_refctl_n63));
   NOR4_X2 U_refctl_U108 (.ZN(U_refctl_n63), 
	.A4(U_refctl_n56), 
	.A3(U_refctl_n57), 
	.A2(U_refctl_n58), 
	.A1(U_refctl_n59));
   NAND4_X2 U_refctl_U107 (.ZN(U_refctl_n56), 
	.A4(U_refctl_n52), 
	.A3(U_refctl_n53), 
	.A2(U_refctl_n54), 
	.A1(U_refctl_n55));
   NOR4_X2 U_refctl_U106 (.ZN(U_refctl_n55), 
	.A4(U_refctl_n48), 
	.A3(U_refctl_n49), 
	.A2(U_refctl_n50), 
	.A1(U_refctl_n51));
   OAI221_X2 U_refctl_U105 (.ZN(U_refctl_n48), 
	.C2(FE_PHN1663_U_refctl_count_0_), 
	.C1(cr_t_ref[0]), 
	.B2(U_refctl_n47), 
	.B1(U_refctl_count_1_), 
	.A(U_refctl_n46));
   AOI22_X2 U_refctl_U104 (.ZN(U_refctl_n46), 
	.B2(FE_PHN1663_U_refctl_count_0_), 
	.B1(cr_t_ref[0]), 
	.A2(U_refctl_n47), 
	.A1(U_refctl_count_1_));
   NOR3_X2 U_refctl_U103 (.ZN(U_refctl_n33), 
	.A3(cr_t_ref[0]), 
	.A2(cr_t_ref[1]), 
	.A1(cr_t_ref[2]));
   NOR2_X2 U_refctl_U102 (.ZN(U_refctl_n32), 
	.A2(cr_t_ref[0]), 
	.A1(cr_t_ref[1]));
   NOR2_X2 U_refctl_U101 (.ZN(U_refctl_N30), 
	.A2(U_refctl_n45), 
	.A1(cr_t_ref[15]));
   NAND2_X2 U_refctl_U100 (.ZN(U_refctl_n45), 
	.A2(U_cr_n123), 
	.A1(U_refctl_n44));
   NOR2_X2 U_refctl_U98 (.ZN(U_refctl_n44), 
	.A2(U_refctl_n43), 
	.A1(cr_t_ref[13]));
   NAND2_X2 U_refctl_U97 (.ZN(U_refctl_n43), 
	.A2(U_cr_n122), 
	.A1(U_refctl_n42));
   NOR2_X2 U_refctl_U95 (.ZN(U_refctl_n42), 
	.A2(U_refctl_n41), 
	.A1(cr_t_ref[11]));
   NAND2_X2 U_refctl_U94 (.ZN(U_refctl_n41), 
	.A2(U_cr_n129), 
	.A1(U_refctl_n40));
   NOR2_X2 U_refctl_U92 (.ZN(U_refctl_n40), 
	.A2(U_refctl_n39), 
	.A1(cr_t_ref[9]));
   NAND2_X2 U_refctl_U91 (.ZN(U_refctl_n39), 
	.A2(U_cr_n118), 
	.A1(U_refctl_n38));
   NOR2_X2 U_refctl_U89 (.ZN(U_refctl_n38), 
	.A2(U_refctl_n37), 
	.A1(cr_t_ref[7]));
   NAND2_X2 U_refctl_U88 (.ZN(U_refctl_n37), 
	.A2(U_cr_n121), 
	.A1(U_refctl_n36));
   NOR2_X2 U_refctl_U86 (.ZN(U_refctl_n36), 
	.A2(U_refctl_n35), 
	.A1(cr_t_ref[5]));
   NAND2_X2 U_refctl_U85 (.ZN(U_refctl_n35), 
	.A2(U_cr_n130), 
	.A1(U_refctl_n34));
   NOR4_X2 U_refctl_U83 (.ZN(U_refctl_n34), 
	.A4(cr_t_ref[0]), 
	.A3(cr_t_ref[1]), 
	.A2(cr_t_ref[2]), 
	.A1(cr_t_ref[3]));
   XNOR2_X2 U_refctl_U82 (.ZN(U_refctl_n61), 
	.B(U_refctl_N26), 
	.A(FE_PHN1424_U_refctl_count_12_));
   XNOR2_X2 U_refctl_U81 (.ZN(U_refctl_N26), 
	.B(U_cr_n122), 
	.A(U_refctl_n42));
   XNOR2_X2 U_refctl_U80 (.ZN(U_refctl_n62), 
	.B(U_refctl_N25), 
	.A(U_refctl_count_11_));
   XNOR2_X2 U_refctl_U79 (.ZN(U_refctl_N25), 
	.B(U_refctl_n41), 
	.A(cr_t_ref[11]));
   XNOR2_X2 U_refctl_U78 (.ZN(U_refctl_n52), 
	.B(U_refctl_N21), 
	.A(U_refctl_count_7_));
   XNOR2_X2 U_refctl_U77 (.ZN(U_refctl_N21), 
	.B(U_refctl_n37), 
	.A(cr_t_ref[7]));
   XNOR2_X2 U_refctl_U76 (.ZN(U_refctl_n53), 
	.B(U_refctl_N19), 
	.A(U_refctl_count_5_));
   XNOR2_X2 U_refctl_U75 (.ZN(U_refctl_N19), 
	.B(U_refctl_n35), 
	.A(cr_t_ref[5]));
   XNOR2_X2 U_refctl_U74 (.ZN(U_refctl_N20), 
	.B(U_cr_n121), 
	.A(U_refctl_n36));
   XOR2_X2 U_refctl_U73 (.Z(U_refctl_n47), 
	.B(cr_t_ref[0]), 
	.A(cr_t_ref[1]));
   XOR2_X2 U_refctl_U72 (.Z(U_refctl_N17), 
	.B(U_refctl_n33), 
	.A(cr_t_ref[3]));
   XOR2_X2 U_refctl_U71 (.Z(U_refctl_N16), 
	.B(U_refctl_n32), 
	.A(cr_t_ref[2]));
   XOR2_X2 U_refctl_U70 (.Z(U_refctl_n51), 
	.B(U_refctl_N18), 
	.A(U_refctl_count_4_));
   XNOR2_X2 U_refctl_U69 (.ZN(U_refctl_N18), 
	.B(U_cr_n130), 
	.A(U_refctl_n34));
   XOR2_X2 U_refctl_U68 (.Z(U_refctl_n57), 
	.B(U_refctl_N23), 
	.A(U_refctl_count_9_));
   XNOR2_X2 U_refctl_U67 (.ZN(U_refctl_N23), 
	.B(U_refctl_n39), 
	.A(cr_t_ref[9]));
   XOR2_X2 U_refctl_U66 (.Z(U_refctl_n58), 
	.B(U_refctl_N24), 
	.A(U_refctl_count_10_));
   XNOR2_X2 U_refctl_U65 (.ZN(U_refctl_N24), 
	.B(U_cr_n129), 
	.A(U_refctl_n40));
   XOR2_X2 U_refctl_U64 (.Z(U_refctl_n59), 
	.B(U_refctl_N22), 
	.A(U_refctl_count_8_));
   XNOR2_X2 U_refctl_U63 (.ZN(U_refctl_N22), 
	.B(U_cr_n118), 
	.A(U_refctl_n38));
   XOR2_X2 U_refctl_U62 (.Z(U_refctl_n65), 
	.B(U_refctl_N28), 
	.A(U_refctl_count_14_));
   XNOR2_X2 U_refctl_U61 (.ZN(U_refctl_N28), 
	.B(U_cr_n123), 
	.A(U_refctl_n44));
   XOR2_X2 U_refctl_U60 (.Z(U_refctl_n66), 
	.B(U_refctl_N29), 
	.A(U_refctl_count_15_));
   XNOR2_X2 U_refctl_U59 (.ZN(U_refctl_N29), 
	.B(U_refctl_n45), 
	.A(cr_t_ref[15]));
   XNOR2_X2 U_refctl_U58 (.ZN(U_refctl_n60), 
	.B(U_refctl_N27), 
	.A(U_refctl_count_13_));
   XNOR2_X2 U_refctl_U57 (.ZN(U_refctl_N27), 
	.B(U_refctl_n43), 
	.A(cr_t_ref[13]));
   XOR2_X1 U_refctl_U55 (.Z(U_refctl_n50), 
	.B(U_refctl_N16), 
	.A(U_refctl_count_2_));
   XOR2_X1 U_refctl_U54 (.Z(U_refctl_n49), 
	.B(U_refctl_N17), 
	.A(U_refctl_count_3_));
   XNOR2_X1 U_refctl_U53 (.ZN(U_refctl_n54), 
	.B(U_refctl_N20), 
	.A(U_refctl_count_6_));
   INV_X2 U_refctl_U52 (.ZN(U_refctl_n118), 
	.A(U_refctl_N21));
   OAI21_X1 U_refctl_U51 (.ZN(U_refctl_n95), 
	.B2(FE_PHN1419_U_refctl_count_6_), 
	.B1(U_refctl_n108), 
	.A(U_refctl_n109));
   OAI21_X1 U_refctl_U50 (.ZN(U_refctl_n96), 
	.B2(FE_PHN1420_U_refctl_count_8_), 
	.B1(U_refctl_n110), 
	.A(U_refctl_n113));
   OAI211_X1 U_refctl_U49 (.ZN(U_refctl_n114), 
	.C2(U_refctl_n80), 
	.C1(U_refctl_N25), 
	.B(U_refctl_n90), 
	.A(U_refctl_N24));
   OAI21_X1 U_refctl_U48 (.ZN(U_refctl_n93), 
	.B2(FE_PHN1421_U_refctl_count_10_), 
	.B1(U_refctl_n111), 
	.A(U_refctl_n98));
   INV_X1 U_refctl_U47 (.ZN(U_refctl_n121), 
	.A(U_refctl_N26));
   OAI21_X1 U_refctl_U46 (.ZN(U_refctl_n94), 
	.B2(FE_PHN1424_U_refctl_count_12_), 
	.B1(U_refctl_n99), 
	.A(U_refctl_n100));
   INV_X2 U_refctl_U45 (.ZN(U_refctl_n103), 
	.A(U_refctl_n104));
   NAND2_X1 U_refctl_U44 (.ZN(U_refctl_n126), 
	.A2(U_refctl_N31), 
	.A1(U_refctl_current_state_0_));
   INV_X2 U_refctl_U43 (.ZN(U_refctl_n97), 
	.A(U_refctl_N31));
   OAI21_X1 U_refctl_U42 (.ZN(U_refctl_n123), 
	.B2(U_refctl_current_state_1_), 
	.B1(U_refctl_n126), 
	.A(ctl_auto_ref_en));
   NOR2_X1 U_refctl_U41 (.ZN(U_refctl_n76), 
	.A2(U_refctl_n96), 
	.A1(U_refctl_n112));
   NOR2_X1 U_refctl_U40 (.ZN(U_refctl_n75), 
	.A2(U_refctl_n95), 
	.A1(U_refctl_n112));
   NOR2_X1 U_refctl_U39 (.ZN(U_refctl_n79), 
	.A2(U_refctl_n93), 
	.A1(U_refctl_n112));
   NOR2_X1 U_refctl_U38 (.ZN(U_refctl_n82), 
	.A2(U_refctl_n94), 
	.A1(U_refctl_n112));
   AOI22_X1 U_refctl_U37 (.ZN(U_refctl_count_next_3_), 
	.B2(U_refctl_n30), 
	.B1(U_refctl_n74), 
	.A2(U_refctl_count_3_), 
	.A1(U_refctl_n28));
   NAND4_X1 U_refctl_U36 (.ZN(U_refctl_n30), 
	.A4(U_refctl_n29), 
	.A3(U_refctl_count_1_), 
	.A2(U_refctl_count_2_), 
	.A1(FE_PHN1663_U_refctl_count_0_));
   INV_X1 U_refctl_U35 (.ZN(U_refctl_n29), 
	.A(U_refctl_n112));
   NOR2_X1 U_refctl_U34 (.ZN(U_refctl_n28), 
	.A2(U_refctl_n27), 
	.A1(U_refctl_count_next_0_));
   AOI21_X1 U_refctl_U33 (.ZN(U_refctl_n27), 
	.B2(U_refctl_count_2_), 
	.B1(U_refctl_count_1_), 
	.A(U_refctl_n112));
   OAI222_X1 U_refctl_U32 (.ZN(U_refctl_n116), 
	.C2(U_refctl_n80), 
	.C1(U_refctl_N25), 
	.B2(U_refctl_n90), 
	.B1(U_refctl_N24), 
	.A2(U_refctl_N23), 
	.A1(FE_PHN1574_U_refctl_n78));
   AOI221_X1 U_refctl_U30 (.ZN(U_refctl_count_next_2_), 
	.C2(U_refctl_n25), 
	.C1(U_refctl_n77), 
	.B2(U_refctl_n25), 
	.B1(U_refctl_n23), 
	.A(U_refctl_n112));
   NAND3_X1 U_refctl_U29 (.ZN(U_refctl_n25), 
	.A3(U_refctl_n77), 
	.A2(U_refctl_count_1_), 
	.A1(FE_PHN1663_U_refctl_count_0_));
   NOR2_X1 U_refctl_U27 (.ZN(U_refctl_n23), 
	.A2(U_refctl_n73), 
	.A1(U_refctl_n83));
   OAI221_X1 U_refctl_U26 (.ZN(U_refctl_n117), 
	.C2(U_refctl_n22), 
	.C1(U_refctl_n88), 
	.B2(U_refctl_n21), 
	.B1(U_refctl_N20), 
	.A(U_refctl_n11));
   AND2_X1 U_refctl_U25 (.ZN(U_refctl_n22), 
	.A2(U_refctl_n21), 
	.A1(U_refctl_N20));
   AOI222_X1 U_refctl_U24 (.ZN(U_refctl_n21), 
	.C2(U_refctl_n20), 
	.C1(U_refctl_n19), 
	.B2(U_refctl_n20), 
	.B1(U_refctl_count_5_), 
	.A2(U_refctl_n19), 
	.A1(U_refctl_count_5_));
   INV_X1 U_refctl_U23 (.ZN(U_refctl_n20), 
	.A(U_refctl_N19));
   AOI21_X1 U_refctl_U22 (.ZN(U_refctl_n19), 
	.B2(U_refctl_N18), 
	.B1(U_refctl_n84), 
	.A(U_refctl_n18));
   AOI221_X1 U_refctl_U21 (.ZN(U_refctl_n18), 
	.C2(U_refctl_n15), 
	.C1(U_refctl_n16), 
	.B2(U_refctl_n15), 
	.B1(U_refctl_n14), 
	.A(U_refctl_n17));
   OAI22_X1 U_refctl_U20 (.ZN(U_refctl_n17), 
	.B2(U_refctl_n84), 
	.B1(U_refctl_N18), 
	.A2(U_refctl_n74), 
	.A1(U_refctl_N17));
   OAI22_X1 U_refctl_U19 (.ZN(U_refctl_n16), 
	.B2(U_refctl_n12), 
	.B1(U_refctl_n73), 
	.A2(U_refctl_n77), 
	.A1(U_refctl_N16));
   AOI22_X1 U_refctl_U18 (.ZN(U_refctl_n15), 
	.B2(U_refctl_n77), 
	.B1(U_refctl_N16), 
	.A2(U_refctl_n74), 
	.A1(U_refctl_N17));
   AOI22_X1 U_refctl_U17 (.ZN(U_refctl_n14), 
	.B2(n87), 
	.B1(U_refctl_n83), 
	.A2(U_refctl_n12), 
	.A1(U_refctl_n73));
   INV_X1 U_refctl_U15 (.ZN(U_refctl_n12), 
	.A(U_refctl_n47));
   NAND2_X1 U_refctl_U14 (.ZN(U_refctl_n11), 
	.A2(U_refctl_count_7_), 
	.A1(U_refctl_n118));
   OAI221_X1 U_refctl_U13 (.ZN(U_refctl_n124), 
	.C2(U_refctl_n10), 
	.C1(U_refctl_n5), 
	.B2(U_refctl_n122), 
	.B1(U_refctl_n5), 
	.A(ctl_ref_ack));
   OAI21_X1 U_refctl_U12 (.ZN(U_refctl_n10), 
	.B2(U_refctl_n7), 
	.B1(U_refctl_n116), 
	.A(U_refctl_n9));
   AOI21_X1 U_refctl_U11 (.ZN(U_refctl_n9), 
	.B2(U_refctl_n80), 
	.B1(U_refctl_N25), 
	.A(U_refctl_n8));
   OAI21_X1 U_refctl_U10 (.ZN(U_refctl_n8), 
	.B2(U_refctl_n115), 
	.B1(U_refctl_n116), 
	.A(U_refctl_n114));
   OAI21_X1 U_refctl_U9 (.ZN(U_refctl_n7), 
	.B2(U_refctl_n87), 
	.B1(U_refctl_N22), 
	.A(U_refctl_n6));
   OAI21_X1 U_refctl_U8 (.ZN(U_refctl_n6), 
	.B2(U_refctl_n118), 
	.B1(U_refctl_count_7_), 
	.A(U_refctl_n117));
   OAI211_X1 U_refctl_U7 (.ZN(U_refctl_n5), 
	.C2(U_refctl_n2), 
	.C1(U_refctl_n120), 
	.B(U_refctl_n4), 
	.A(U_refctl_n3));
   OAI211_X1 U_refctl_U6 (.ZN(U_refctl_n4), 
	.C2(U_refctl_n81), 
	.C1(U_refctl_N29), 
	.B(U_refctl_n86), 
	.A(U_refctl_N28));
   AOI21_X1 U_refctl_U5 (.ZN(U_refctl_n3), 
	.B2(U_refctl_N29), 
	.B1(U_refctl_n81), 
	.A(U_refctl_N30));
   AOI22_X1 U_refctl_U4 (.ZN(U_refctl_n2), 
	.B2(U_refctl_n1), 
	.B1(U_refctl_N26), 
	.A2(FE_PHN1411_U_refctl_n91), 
	.A1(U_refctl_N27));
   NOR2_X1 U_refctl_U3 (.ZN(U_refctl_n1), 
	.A2(U_refctl_n119), 
	.A1(FE_PHN1424_U_refctl_count_12_));
   DFFR_X1 U_refctl_count_reg_0_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_refctl_n83), 
	.Q(U_refctl_count_0_), 
	.D(FE_PHN4543_U_refctl_count_next_0_), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_refctl_count_reg_10_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_refctl_n90), 
	.Q(U_refctl_count_10_), 
	.D(U_refctl_n79), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_refctl_count_reg_11_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_refctl_n80), 
	.Q(U_refctl_count_11_), 
	.D(FE_PHN1207_U_refctl_count_next_11_), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_refctl_count_reg_12_ (.RN(FE_OFN31_HRESETn), 
	.Q(U_refctl_count_12_), 
	.D(U_refctl_n82), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_refctl_count_reg_13_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_refctl_n91), 
	.Q(U_refctl_count_13_), 
	.D(FE_PHN1201_U_refctl_count_next_13_), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_refctl_count_reg_14_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_refctl_n86), 
	.Q(U_refctl_count_14_), 
	.D(FE_PHN1414_U_refctl_count_next_14_), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_refctl_count_reg_15_ (.RN(FE_OFN31_HRESETn), 
	.QN(U_refctl_n81), 
	.Q(U_refctl_count_15_), 
	.D(FE_PHN1476_U_refctl_count_next_15_), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_refctl_count_reg_1_ (.RN(FE_OFN151_HRESETn), 
	.QN(U_refctl_n73), 
	.Q(U_refctl_count_1_), 
	.D(FE_PHN1557_U_refctl_count_next_1_), 
	.CK(HCLK__L5_N32));
   DFFR_X1 U_refctl_count_reg_2_ (.RN(FE_OFN57_HRESETn), 
	.QN(U_refctl_n77), 
	.Q(U_refctl_count_2_), 
	.D(FE_PHN3607_U_refctl_count_next_2_), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_refctl_count_reg_3_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_refctl_n74), 
	.Q(U_refctl_count_3_), 
	.D(FE_PHN1091_U_refctl_count_next_3_), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_refctl_count_reg_4_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_refctl_n84), 
	.Q(U_refctl_count_4_), 
	.D(FE_PHN1089_U_refctl_count_next_4_), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_refctl_count_reg_5_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_refctl_n85), 
	.Q(U_refctl_count_5_), 
	.D(FE_PHN1403_U_refctl_count_next_5_), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_refctl_count_reg_6_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_refctl_n88), 
	.Q(U_refctl_count_6_), 
	.D(U_refctl_n75), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_refctl_count_reg_7_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_refctl_n89), 
	.Q(U_refctl_count_7_), 
	.D(FE_PHN1185_U_refctl_count_next_7_), 
	.CK(HCLK__L5_N36));
   DFFR_X1 U_refctl_count_reg_8_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_refctl_n87), 
	.Q(U_refctl_count_8_), 
	.D(U_refctl_n76), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_refctl_count_reg_9_ (.RN(FE_OFN46_HRESETn), 
	.QN(U_refctl_n78), 
	.Q(U_refctl_count_9_), 
	.D(FE_PHN1203_U_refctl_count_next_9_), 
	.CK(HCLK__L5_N35));
   DFFR_X1 U_refctl_current_state_reg_1_ (.RN(FE_OFN39_HRESETn), 
	.QN(U_refctl_n92), 
	.Q(U_refctl_current_state_1_), 
	.D(FE_PHN4727_U_refctl_ref_req_next), 
	.CK(HCLK__L5_N11));
   DFFR_X1 U_refctl_ref_req_reg (.RN(FE_OFN183_HRESETn), 
	.QN(n84), 
	.Q(debug_ref_req), 
	.D(FE_PHN4727_U_refctl_ref_req_next), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_refctl_current_state_reg_0_ (.RN(FE_OFN39_HRESETn), 
	.Q(U_refctl_current_state_0_), 
	.D(FE_PHN1494_U_refctl_next_state_0_), 
	.CK(HCLK__L5_N11));
   AND3_X4 U_dmc_U76 (.ZN(U_dmc_n52), 
	.A3(U_dmc_n19), 
	.A2(U_dmc_n8), 
	.A1(U_dmc_n63));
   AND2_X4 U_dmc_U75 (.ZN(U_dmc_n8), 
	.A2(U_dmc_n6), 
	.A1(U_dmc_n62));
   NOR2_X2 U_dmc_U73 (.ZN(U_dmc_n39), 
	.A2(U_dmc_n33), 
	.A1(U_dmc_n70));
   AND4_X4 U_dmc_U72 (.ZN(U_dmc_n12), 
	.A4(U_dmc_n63), 
	.A3(U_dmc_n62), 
	.A2(hiu_wrapped_burst), 
	.A1(FE_PHN1056_U_dmc_terminate));
   NOR3_X2 U_dmc_U69 (.ZN(U_dmc_n18), 
	.A3(U_dmc_n58), 
	.A2(U_dmc_data_cnt_5_), 
	.A1(FE_PHN902_U_dmc_data_cnt_4_));
   NAND2_X2 U_dmc_U68 (.ZN(U_dmc_n20), 
	.A2(U_dmc_n18), 
	.A1(U_dmc_n63));
   NAND2_X2 U_dmc_U67 (.ZN(U_dmc_n59), 
	.A2(U_dmc_n6), 
	.A1(U_dmc_n20));
   NAND2_X2 U_dmc_U66 (.ZN(U_dmc_n15), 
	.A2(U_dmc_dmc_cs_1_), 
	.A1(FE_PHN967_U_dmc_n4));
   NOR2_X2 U_dmc_U65 (.ZN(U_dmc_n53), 
	.A2(U_dmc_dmc_cs_2_), 
	.A1(U_dmc_n15));
   INV_X4 U_dmc_U64 (.ZN(U_dmc_n27), 
	.A(U_dmc_n53));
   NAND2_X2 U_dmc_U63 (.ZN(U_dmc_n10), 
	.A2(U_dmc_dmc_cs_0_), 
	.A1(U_dmc_dmc_cs_1_));
   NOR2_X2 U_dmc_U62 (.ZN(U_dmc_n55), 
	.A2(U_dmc_dmc_cs_2_), 
	.A1(U_dmc_n10));
   AOI211_X2 U_dmc_U61 (.ZN(U_dmc_n30), 
	.C2(U_dmc_n24), 
	.C1(U_dmc_n25), 
	.B(hiu_terminate), 
	.A(U_dmc_n23));
   NAND2_X2 U_dmc_U60 (.ZN(U_dmc_n11), 
	.A2(U_dmc_dmc_cs_0_), 
	.A1(FE_PHN943_U_dmc_n7));
   NOR2_X2 U_dmc_U59 (.ZN(U_dmc_n54), 
	.A2(U_dmc_dmc_cs_2_), 
	.A1(U_dmc_n11));
   OAI211_X2 U_dmc_U58 (.ZN(U_dmc_N23), 
	.C2(U_dmc_n27), 
	.C1(U_dmc_n32), 
	.B(U_dmc_n26), 
	.A(U_dmc_n30));
   INV_X4 U_dmc_U57 (.ZN(U_dmc_n31), 
	.A(FE_PHN944_U_dmc_n54));
   OAI211_X2 U_dmc_U56 (.ZN(U_dmc_N24), 
	.C2(U_dmc_n31), 
	.C1(U_dmc_n32), 
	.B(U_dmc_n29), 
	.A(U_dmc_n30));
   NAND2_X2 U_dmc_U55 (.ZN(U_dmc_n61), 
	.A2(FE_PHN943_U_dmc_n7), 
	.A1(FE_PHN967_U_dmc_n4));
   NAND2_X2 U_dmc_U54 (.ZN(U_dmc_n62), 
	.A2(U_dmc_n27), 
	.A1(U_dmc_n31));
   AOI22_X2 U_dmc_U53 (.ZN(U_dmc_n60), 
	.B2(U_dmc_n59), 
	.B1(U_dmc_n62), 
	.A2(U_dmc_n55), 
	.A1(FE_PHN1056_U_dmc_terminate));
   AOI21_X2 U_dmc_U51 (.ZN(U_dmc_n70), 
	.B2(U_dmc_n25), 
	.B1(N28), 
	.A(U_dmc_n21));
   NAND2_X2 U_dmc_U50 (.ZN(U_dmc_n48), 
	.A2(U_dmc_n34), 
	.A1(U_dmc_n35));
   NOR2_X2 U_dmc_U49 (.ZN(U_dmc_n47), 
	.A2(FE_PHN1160_U_dmc_n48), 
	.A1(U_dmc_n51));
   NAND2_X2 U_dmc_U47 (.ZN(U_dmc_n46), 
	.A2(U_dmc_n45), 
	.A1(U_dmc_n47));
   NOR2_X2 U_dmc_U45 (.ZN(U_dmc_n42), 
	.A2(U_dmc_n43), 
	.A1(U_dmc_n46));
   NAND2_X2 U_dmc_U44 (.ZN(U_dmc_n41), 
	.A2(U_dmc_n40), 
	.A1(U_dmc_n42));
   NOR2_X2 U_dmc_U43 (.ZN(U_dmc_n50), 
	.A2(U_dmc_n52), 
	.A1(U_dmc_n39));
   AOI21_X2 U_dmc_U42 (.ZN(U_dmc_n44), 
	.B2(U_dmc_n46), 
	.B1(U_dmc_n43), 
	.A(U_dmc_n42));
   NOR2_X2 U_dmc_U41 (.ZN(U_dmc_data_cnt_nxt[3]), 
	.A2(U_dmc_n50), 
	.A1(U_dmc_n44));
   AOI21_X2 U_dmc_U40 (.ZN(U_dmc_n49), 
	.B2(FE_PHN1160_U_dmc_n48), 
	.B1(U_dmc_n51), 
	.A(U_dmc_n47));
   NOR2_X2 U_dmc_U39 (.ZN(U_dmc_data_cnt_nxt[1]), 
	.A2(U_dmc_n50), 
	.A1(U_dmc_n49));
   NAND3_X2 U_dmc_U38 (.ZN(U_dmc_n69), 
	.A3(U_dmc_n64), 
	.A2(hiu_wrapped_burst), 
	.A1(U_dmc_n8));
   AOI21_X2 U_dmc_U37 (.ZN(U_dmc_n67), 
	.B2(U_dmc_n66), 
	.B1(FE_PHN944_U_dmc_n54), 
	.A(U_dmc_n52));
   AOI21_X1 U_dmc_U36 (.ZN(U_dmc_n26), 
	.B2(U_dmc_n28), 
	.B1(hiu_rw), 
	.A(FE_PHN944_U_dmc_n54));
   INV_X1 U_dmc_U35 (.ZN(U_dmc_n19), 
	.A(U_dmc_n18));
   AOI22_X2 U_dmc_U34 (.ZN(U_dmc_n40), 
	.B2(U_dmc_n52), 
	.B1(FE_PHN902_U_dmc_data_cnt_4_), 
	.A2(FE_OFN215_hiu_burst_size_4_), 
	.A1(U_dmc_n39));
   INV_X1 U_dmc_U33 (.ZN(U_dmc_n64), 
	.A(U_dmc_n20));
   OAI211_X1 U_dmc_U32 (.ZN(U_dmc_n13), 
	.C2(hiu_rw), 
	.C1(U_dmc_n70), 
	.B(U_dmc_n69), 
	.A(U_dmc_n65));
   INV_X1 U_dmc_U31 (.ZN(U_dmc_n32), 
	.A(FE_PHN3197_U_dmc_n59));
   INV_X1 U_dmc_U30 (.ZN(U_dmc_n33), 
	.A(U_dmc_n63));
   NOR3_X1 U_dmc_U29 (.ZN(U_dmc_n25), 
	.A3(U_dmc_dmc_cs_0_), 
	.A2(U_dmc_dmc_cs_1_), 
	.A1(U_dmc_dmc_cs_2_));
   OR4_X2 U_dmc_U28 (.ZN(U_dmc_n58), 
	.A4(U_dmc_data_cnt_3_), 
	.A3(U_dmc_data_cnt_0_), 
	.A2(U_dmc_data_cnt_2_), 
	.A1(U_dmc_data_cnt_1_));
   INV_X1 U_dmc_U27 (.ZN(U_dmc_n22), 
	.A(U_dmc_n55));
   NOR2_X1 U_dmc_U26 (.ZN(U_dmc_n21), 
	.A2(FE_PHN1056_U_dmc_terminate), 
	.A1(U_dmc_n22));
   OAI21_X1 U_dmc_U25 (.ZN(U_dmc_n23), 
	.B2(U_dmc_n6), 
	.B1(U_dmc_n22), 
	.A(U_dmc_n5));
   AOI21_X1 U_dmc_U24 (.ZN(U_dmc_n29), 
	.B2(U_dmc_n28), 
	.B1(U_dsdc_n1438), 
	.A(U_dmc_n53));
   AOI22_X1 U_dmc_U22 (.ZN(U_dmc_n65), 
	.B2(U_dmc_n66), 
	.B1(U_dmc_n53), 
	.A2(U_dmc_n52), 
	.A1(U_dmc_dmc_cs_1_));
   NAND2_X1 U_dmc_U21 (.ZN(U_dmc_n34), 
	.A2(U_dmc_data_cnt_1_), 
	.A1(U_dmc_n52));
   OR2_X1 U_dmc_U18 (.ZN(U_dmc_n68), 
	.A2(U_dmc_n67), 
	.A1(FE_PHN967_U_dmc_n4));
   INV_X2 U_dmc_U17 (.ZN(U_dmc_n24), 
	.A(N28));
   NAND2_X1 U_dmc_U15 (.ZN(U_dmc_n35), 
	.A2(hiu_burst_size[1]), 
	.A1(U_dmc_n39));
   NOR2_X1 U_dmc_U14 (.ZN(U_dmc_data_cnt_nxt[0]), 
	.A2(U_dmc_n50), 
	.A1(U_dmc_n51));
   OR2_X1 U_dmc_U13 (.ZN(U_dmc_n28), 
	.A2(U_dmc_n55), 
	.A1(U_dmc_n25));
   INV_X4 U_dmc_U12 (.ZN(U_dmc_n16), 
	.A(FE_OFN215_hiu_burst_size_4_));
   NOR2_X1 U_dmc_U11 (.ZN(U_dmc_n66), 
	.A2(U_dmc_n63), 
	.A1(FE_PHN1056_U_dmc_terminate));
   OAI211_X1 U_dmc_U10 (.ZN(U_dmc_n14), 
	.C2(U_dsdc_n1438), 
	.C1(U_dmc_n70), 
	.B(U_dmc_n68), 
	.A(U_dmc_n69));
   AOI221_X1 U_dmc_U9 (.ZN(U_dmc_data_cnt_nxt[2]), 
	.C2(U_dmc_n46), 
	.C1(U_dmc_n45), 
	.B2(U_dmc_n46), 
	.B1(U_dmc_n47), 
	.A(U_dmc_n50));
   AOI221_X1 U_dmc_U8 (.ZN(U_dmc_data_cnt_nxt[4]), 
	.C2(U_dmc_n41), 
	.C1(FE_PHN3454_U_dmc_n40), 
	.B2(U_dmc_n41), 
	.B1(U_dmc_n42), 
	.A(U_dmc_n50));
   AOI211_X1 U_dmc_U7 (.ZN(U_dmc_data_cnt_nxt[5]), 
	.C2(U_dmc_n2), 
	.C1(U_dmc_n41), 
	.B(U_dmc_n3), 
	.A(U_dmc_n50));
   NOR2_X1 U_dmc_U6 (.ZN(U_dmc_n3), 
	.A2(U_dmc_n2), 
	.A1(U_dmc_n41));
   AOI22_X1 U_dmc_U5 (.ZN(U_dmc_n2), 
	.B2(U_dmc_n39), 
	.B1(hiu_burst_size[5]), 
	.A2(U_dmc_data_cnt_5_), 
	.A1(U_dmc_n52));
   INV_X1 U_dmc_U4 (.ZN(U_dmc_n51), 
	.A(FE_PHN3193_U_dmc_n1));
   AOI22_X1 U_dmc_U3 (.ZN(U_dmc_n1), 
	.B2(U_dmc_n52), 
	.B1(U_dmc_data_cnt_0_), 
	.A2(U_dmc_n39), 
	.A1(FE_OFN221_hiu_burst_size_0_));
   DFFR_X2 U_dmc_terminate_reg (.RN(FE_OFN183_HRESETn), 
	.QN(U_dmc_n6), 
	.Q(U_dmc_terminate), 
	.D(hiu_terminate), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dmc_dmc_cs_reg_0_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dmc_n4), 
	.Q(U_dmc_dmc_cs_0_), 
	.D(FE_PHN1000_U_dmc_n14), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dmc_dmc_cs_reg_1_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dmc_n7), 
	.Q(U_dmc_dmc_cs_1_), 
	.D(FE_PHN3345_U_dmc_n13), 
	.CK(HCLK__L5_N12));
   DFFR_X2 U_dmc_dmc_cs_reg_2_ (.RN(FE_OFN183_HRESETn), 
	.QN(U_dmc_n5), 
	.Q(U_dmc_dmc_cs_2_), 
	.D(FE_PHN3870_U_dmc_n12), 
	.CK(HCLK__L5_N12));
   DFFS_X2 U_dmc_miu_pop_n_reg (.SN(FE_OFN183_HRESETn), 
	.Q(dmc_pop_n), 
	.D(FE_PHN777_U_dmc_N23), 
	.CK(HCLK__L5_N12));
   DFFS_X2 U_dmc_miu_push_n_reg (.SN(FE_OFN183_HRESETn), 
	.Q(dmc_push_n), 
	.D(FE_PHN713_U_dmc_N24), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dmc_data_cnt_reg_5_ (.RN(FE_OFN183_HRESETn), 
	.Q(U_dmc_data_cnt_5_), 
	.D(FE_PHN4713_U_dmc_data_cnt_nxt_5_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dmc_data_cnt_reg_4_ (.RN(FE_OFN183_HRESETn), 
	.Q(U_dmc_data_cnt_4_), 
	.D(U_dmc_data_cnt_nxt[4]), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dmc_data_cnt_reg_3_ (.RN(FE_OFN183_HRESETn), 
	.Q(U_dmc_data_cnt_3_), 
	.D(U_dmc_data_cnt_nxt[3]), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dmc_data_cnt_reg_2_ (.RN(FE_OFN183_HRESETn), 
	.Q(U_dmc_data_cnt_2_), 
	.D(FE_PHN1217_U_dmc_data_cnt_nxt_2_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dmc_data_cnt_reg_1_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dmc_data_cnt_1_), 
	.D(FE_PHN1340_U_dmc_data_cnt_nxt_1_), 
	.CK(HCLK__L5_N12));
   DFFR_X1 U_dmc_data_cnt_reg_0_ (.RN(FE_OFN64_HRESETn), 
	.Q(U_dmc_data_cnt_0_), 
	.D(U_dmc_data_cnt_nxt[0]), 
	.CK(HCLK__L5_N12));
   NAND2_X2 U_dsdc_U_minmax1_dwbb_U40 (.ZN(U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_1_), 
	.A2(U_dsdc_U_minmax1_dwbb_n2), 
	.A1(U_dsdc_U_minmax1_dwbb_n26));
   NAND4_X2 U_dsdc_U_minmax1_dwbb_U39 (.ZN(U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_0_), 
	.A4(U_dsdc_U_minmax1_dwbb_n19), 
	.A3(U_dsdc_U_minmax1_dwbb_n20), 
	.A2(U_dsdc_U_minmax1_dwbb_n21), 
	.A1(U_dsdc_U_minmax1_dwbb_n22));
   MUX2_X2 U_dsdc_U_minmax1_dwbb_U37 (.Z(U_dsdc_oldest_bank_0_), 
	.S(U_dsdc_oldest_bank_1_), 
	.B(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_), 
	.A(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_));
   OR2_X1 U_dsdc_U_minmax1_dwbb_U32 (.ZN(U_dsdc_U_minmax1_dwbb_n21), 
	.A2(U_dsdc_bm_bank_age_0__0_), 
	.A1(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_));
   NAND2_X1 U_dsdc_U_minmax1_dwbb_U31 (.ZN(U_dsdc_U_minmax1_dwbb_n20), 
	.A2(FE_PHN897_U_dsdc_n352), 
	.A1(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_));
   NAND2_X1 U_dsdc_U_minmax1_dwbb_U30 (.ZN(U_dsdc_U_minmax1_dwbb_n19), 
	.A2(U_dsdc_bm_bank_age_3__0_), 
	.A1(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_));
   NAND2_X1 U_dsdc_U_minmax1_dwbb_U29 (.ZN(U_dsdc_U_minmax1_dwbb_n22), 
	.A2(U_dsdc_bm_bank_age_2__0_), 
	.A1(U_dsdc_U_minmax1_dwbb_n24));
   AND2_X2 U_dsdc_U_minmax1_dwbb_U28 (.ZN(U_dsdc_U_minmax1_dwbb_n32), 
	.A2(U_dsdc_U_minmax1_dwbb_n31), 
	.A1(U_dsdc_U_minmax1_dwbb_n33));
   OR2_X2 U_dsdc_U_minmax1_dwbb_U27 (.ZN(U_dsdc_U_minmax1_dwbb_n34), 
	.A2(U_dsdc_U_minmax1_dwbb_n31), 
	.A1(U_dsdc_U_minmax1_dwbb_n33));
   INV_X2 U_dsdc_U_minmax1_dwbb_U26 (.ZN(U_dsdc_U_minmax1_dwbb_n26), 
	.A(U_dsdc_U_minmax1_dwbb_n30));
   AND2_X2 U_dsdc_U_minmax1_dwbb_U25 (.ZN(U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_PI_1_), 
	.A2(U_dsdc_U_minmax1_dwbb_n29), 
	.A1(U_dsdc_U_minmax1_dwbb_n30));
   INV_X1 U_dsdc_U_minmax1_dwbb_U22 (.ZN(U_dsdc_U_minmax1_dwbb_n24), 
	.A(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_));
   OAI21_X1 U_dsdc_U_minmax1_dwbb_U21 (.ZN(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_), 
	.B2(U_dsdc_n303), 
	.B1(U_dsdc_bm_bank_age_2__2_), 
	.A(U_dsdc_U_minmax1_dwbb_n15));
   OAI211_X1 U_dsdc_U_minmax1_dwbb_U20 (.ZN(U_dsdc_U_minmax1_dwbb_n15), 
	.C2(U_dsdc_n336), 
	.C1(U_dsdc_bm_bank_age_3__2_), 
	.B(U_dsdc_U_minmax1_dwbb_n11), 
	.A(U_dsdc_U_minmax1_dwbb_n12));
   NAND2_X1 U_dsdc_U_minmax1_dwbb_U17 (.ZN(U_dsdc_U_minmax1_dwbb_n12), 
	.A2(U_dsdc_n302), 
	.A1(U_dsdc_bm_bank_age_2__1_));
   OAI211_X1 U_dsdc_U_minmax1_dwbb_U16 (.ZN(U_dsdc_U_minmax1_dwbb_n11), 
	.C2(U_dsdc_n302), 
	.C1(U_dsdc_bm_bank_age_2__1_), 
	.B(U_dsdc_bm_bank_age_2__0_), 
	.A(U_dsdc_n304));
   AOI22_X1 U_dsdc_U_minmax1_dwbb_U15 (.ZN(U_dsdc_U_minmax1_dwbb_n33), 
	.B2(U_dsdc_U_minmax1_dwbb_n24), 
	.B1(U_dsdc_bm_bank_age_2__2_), 
	.A2(U_dsdc_bm_bank_age_3__2_), 
	.A1(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_));
   OAI21_X1 U_dsdc_U_minmax1_dwbb_U13 (.ZN(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_), 
	.B2(U_dsdc_n337), 
	.B1(U_dsdc_bm_bank_age_0__2_), 
	.A(U_dsdc_U_minmax1_dwbb_n9));
   OAI211_X1 U_dsdc_U_minmax1_dwbb_U12 (.ZN(U_dsdc_U_minmax1_dwbb_n9), 
	.C2(U_dsdc_n334), 
	.C1(U_dsdc_bm_bank_age_1__2_), 
	.B(U_dsdc_U_minmax1_dwbb_n5), 
	.A(U_dsdc_U_minmax1_dwbb_n6));
   NAND2_X1 U_dsdc_U_minmax1_dwbb_U9 (.ZN(U_dsdc_U_minmax1_dwbb_n6), 
	.A2(U_dsdc_n335), 
	.A1(U_dsdc_bm_bank_age_0__1_));
   OAI211_X1 U_dsdc_U_minmax1_dwbb_U8 (.ZN(U_dsdc_U_minmax1_dwbb_n5), 
	.C2(U_dsdc_n335), 
	.C1(U_dsdc_bm_bank_age_0__1_), 
	.B(U_dsdc_bm_bank_age_0__0_), 
	.A(FE_PHN897_U_dsdc_n352));
   AOI22_X2 U_dsdc_U_minmax1_dwbb_U7 (.ZN(U_dsdc_U_minmax1_dwbb_n30), 
	.B2(U_dsdc_U_minmax1_dwbb_n4), 
	.B1(U_dsdc_bm_bank_age_0__1_), 
	.A2(U_dsdc_bm_bank_age_1__1_), 
	.A1(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_));
   INV_X4 U_dsdc_U_minmax1_dwbb_U6 (.ZN(U_dsdc_U_minmax1_dwbb_n4), 
	.A(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_));
   INV_X1 U_dsdc_U_minmax1_dwbb_U4 (.ZN(U_dsdc_U_minmax1_dwbb_n29), 
	.A(U_dsdc_U_minmax1_dwbb_n2));
   AOI22_X1 U_dsdc_U_minmax1_dwbb_U3 (.ZN(U_dsdc_U_minmax1_dwbb_n2), 
	.B2(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_), 
	.B1(U_dsdc_bm_bank_age_3__1_), 
	.A2(U_dsdc_U_minmax1_dwbb_n24), 
	.A1(U_dsdc_bm_bank_age_2__1_));
   OAI21_X2 U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_UGT1_1_0_0 (.ZN(U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_GT_4_), 
	.B2(U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_0_), 
	.B1(U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_PI_1_), 
	.A(U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_1_));
   AOI21_X2 U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_UGT0_2_0_0 (.ZN(U_dsdc_oldest_bank_1_), 
	.B2(U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_GT_4_), 
	.B1(U_dsdc_U_minmax1_dwbb_n34), 
	.A(U_dsdc_U_minmax1_dwbb_n32));
   OAI33_X1 U17 (.ZN(n45), 
	.B3(U_dsdc_n741), 
	.B2(U_dsdc_n739), 
	.B1(U_dsdc_n740), 
	.A3(U_dsdc_n934), 
	.A2(U_dsdc_n903), 
	.A1(U_dsdc_n165));
   INV_X4 U22 (.ZN(U_dsdc_n744), 
	.A(n45));
   AOI22_X1 U23 (.ZN(U_dmc_n45), 
	.B2(U_dmc_n52), 
	.B1(FE_PHN1418_U_dmc_data_cnt_2_), 
	.A2(U_dmc_n39), 
	.A1(FE_OFN218_hiu_burst_size_2_));
   OAI22_X1 U28 (.ZN(n46), 
	.B2(U_dsdc_n1421), 
	.B1(U_dsdc_n1426), 
	.A2(U_dsdc_n1628), 
	.A1(U_dsdc_n1424));
   NOR3_X1 U46 (.ZN(n47), 
	.A3(n46), 
	.A2(U_dsdc_n967), 
	.A1(U_dsdc_n1872));
   INV_X1 U47 (.ZN(n48), 
	.A(U_dsdc_n1591));
   NAND3_X1 U57 (.ZN(U_dsdc_n1383), 
	.A3(n48), 
	.A2(n47), 
	.A1(U_dsdc_n705));
   AOI22_X2 U58 (.ZN(debug_ad_col_addr_13_), 
	.B2(hiu_addr[14]), 
	.B1(U_addrdec_n220), 
	.A2(hiu_addr[13]), 
	.A1(U_addrdec_n39));
   NOR4_X1 U59 (.ZN(n49), 
	.A4(hiu_burst_size[1]), 
	.A3(FE_OFN221_hiu_burst_size_0_), 
	.A2(hiu_burst_size[3]), 
	.A1(FE_OFN218_hiu_burst_size_2_));
   INV_X1 U60 (.ZN(n50), 
	.A(hiu_burst_size[5]));
   NAND3_X1 U61 (.ZN(U_dmc_n63), 
	.A3(n50), 
	.A2(n49), 
	.A1(U_dmc_n16));
   NOR4_X2 U62 (.ZN(n51), 
	.A4(U_dsdc_r_burst_size_0_), 
	.A3(FE_PHN1890_U_dsdc_r_burst_size_5_), 
	.A2(FE_PHN1892_U_dsdc_r_burst_size_3_), 
	.A1(FE_PHN1888_U_dsdc_r_burst_size_4_));
   NAND2_X1 U63 (.ZN(U_dsdc_n1312), 
	.A2(n51), 
	.A1(U_dsdc_n687));
   NAND2_X1 U64 (.ZN(n52), 
	.A2(hiu_rw), 
	.A1(U_dsdc_n1284));
   NOR3_X1 U65 (.ZN(U_dsdc_n1124), 
	.A3(U_dsdc_n1053), 
	.A2(U_dsdc_n1286), 
	.A1(n52));
   AOI22_X2 U66 (.ZN(n53), 
	.B2(hiu_addr[9]), 
	.B1(U_addrdec_n39), 
	.A2(hiu_addr[10]), 
	.A1(U_addrdec_n220));
   INV_X4 U67 (.ZN(debug_ad_col_addr_9_), 
	.A(n53));
   AOI22_X2 U68 (.ZN(n54), 
	.B2(hiu_addr[14]), 
	.B1(U_addrdec_n39), 
	.A2(hiu_addr[15]), 
	.A1(U_addrdec_n220));
   INV_X4 U69 (.ZN(debug_ad_col_addr_14_), 
	.A(n54));
   AOI22_X2 U70 (.ZN(U_dsdc_n558), 
	.B2(U_dsdc_n998), 
	.B1(U_dsdc_bm_row_addr_0__0_), 
	.A2(U_dsdc_bm_row_addr_1__0_), 
	.A1(U_dsdc_n604));
   AOI22_X1 U71 (.ZN(n55), 
	.B2(U_dmc_n52), 
	.B1(FE_PHN1228_U_dmc_data_cnt_3_), 
	.A2(U_dmc_n39), 
	.A1(hiu_burst_size[3]));
   INV_X1 U72 (.ZN(U_dmc_n43), 
	.A(n55));
   AND2_X1 U73 (.ZN(n56), 
	.A2(U_dsdc_n1253), 
	.A1(U_dsdc_n1254));
   OAI221_X1 U74 (.ZN(U_dsdc_n1270), 
	.C2(U_dsdc_n2013), 
	.C1(n56), 
	.B2(U_dsdc_n1546), 
	.B1(n56), 
	.A(U_dsdc_n1409));
   AOI211_X1 U75 (.ZN(n57), 
	.C2(U_dsdc_n1416), 
	.C1(U_dsdc_n1876), 
	.B(U_dsdc_n1872), 
	.A(U_dsdc_n1412));
   OAI211_X1 U76 (.ZN(n58), 
	.C2(U_dsdc_n2071), 
	.C1(U_dsdc_n1414), 
	.B(n57), 
	.A(U_dsdc_n705));
   OAI21_X1 U77 (.ZN(n59), 
	.B2(U_dsdc_n856), 
	.B1(U_dsdc_n991), 
	.A(U_dsdc_n2072));
   AOI211_X1 U78 (.ZN(U_dsdc_n183), 
	.C2(U_dsdc_n708), 
	.C1(U_dsdc_n721), 
	.B(n59), 
	.A(n58));
   AOI22_X2 U79 (.ZN(n60), 
	.B2(hiu_addr[10]), 
	.B1(U_addrdec_n39), 
	.A2(hiu_addr[11]), 
	.A1(U_addrdec_n220));
   INV_X4 U80 (.ZN(debug_ad_col_addr_10_), 
	.A(n60));
   AOI222_X1 U81 (.ZN(n61), 
	.C2(U_dsdc_bm_row_addr_2__3_), 
	.C1(U_dsdc_n159), 
	.B2(U_dsdc_bm_row_addr_3__3_), 
	.B1(U_dsdc_n978), 
	.A2(U_dsdc_bm_row_addr_1__3_), 
	.A1(U_dsdc_n604));
   INV_X1 U82 (.ZN(U_dsdc_n798), 
	.A(n61));
   AOI22_X1 U83 (.ZN(n62), 
	.B2(U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_), 
	.B1(U_dsdc_bm_bank_age_1__2_), 
	.A2(U_dsdc_bm_bank_age_0__2_), 
	.A1(U_dsdc_U_minmax1_dwbb_n4));
   INV_X1 U84 (.ZN(U_dsdc_U_minmax1_dwbb_n31), 
	.A(n62));
   OAI21_X2 U85 (.ZN(n63), 
	.B2(U_dsdc_n1836), 
	.B1(U_dsdc_n1945), 
	.A(U_dsdc_n1837));
   AOI222_X1 U86 (.ZN(n64), 
	.C2(n63), 
	.C1(U_dsdc_bm_bank_age_2__3_), 
	.B2(n63), 
	.B1(U_dsdc_n1953), 
	.A2(U_dsdc_bm_bank_age_2__3_), 
	.A1(U_dsdc_n1953));
   AOI222_X1 U87 (.ZN(U_dsdc_n1849), 
	.C2(n64), 
	.C1(U_dsdc_n350), 
	.B2(n64), 
	.B1(U_dsdc_n1954), 
	.A2(U_dsdc_n350), 
	.A1(U_dsdc_n1954));
   AOI22_X2 U88 (.ZN(n65), 
	.B2(hiu_addr[15]), 
	.B1(U_addrdec_n39), 
	.A2(hiu_addr[16]), 
	.A1(U_addrdec_n220));
   INV_X4 U89 (.ZN(debug_ad_col_addr_15_), 
	.A(n65));
   NAND3_X1 U90 (.ZN(n66), 
	.A3(FE_PHN1212_U_dsdc_cas_latency_cnt_1_), 
	.A2(FE_PHN2036_U_dsdc_cas_latency_cnt_0_), 
	.A1(U_dsdc_n1393));
   INV_X1 U91 (.ZN(n67), 
	.A(U_dsdc_n1393));
   NAND2_X1 U92 (.ZN(n68), 
	.A2(n67), 
	.A1(U_dsdc_cas_latency_1_));
   OAI211_X1 U93 (.ZN(U_dsdc_N4127), 
	.C2(U_dsdc_n1087), 
	.C1(U_dsdc_n1090), 
	.B(n68), 
	.A(n66));
   OAI33_X1 U94 (.ZN(n69), 
	.B3(U_dsdc_bm_row_addr_0__11_), 
	.B2(U_dsdc_n812), 
	.B1(U_addrdec_n231), 
	.A3(U_dsdc_n814), 
	.A2(U_dsdc_bm_row_addr_0__1_), 
	.A1(U_dsdc_n815));
   INV_X1 U95 (.ZN(U_dsdc_n536), 
	.A(n69));
   OAI211_X1 U96 (.ZN(n70), 
	.C2(U_dsdc_n816), 
	.C1(U_dsdc_n602), 
	.B(U_dsdc_n51), 
	.A(U_dsdc_n488));
   INV_X1 U97 (.ZN(U_dsdc_n499), 
	.A(n70));
   NAND2_X1 U98 (.ZN(n71), 
	.A2(U_dsdc_n753), 
	.A1(U_dsdc_r_cas_latency_3_));
   XNOR2_X1 U99 (.ZN(U_dsdc_DP_OP_1642_126_2028_n19), 
	.B(U_dsdc_DP_OP_1642_126_2028_n85), 
	.A(n71));
   INV_X1 U100 (.ZN(n72), 
	.A(FE_PHN1645_U_cr_n65));
   AOI21_X1 U101 (.ZN(U_addrdec_n75), 
	.B2(n72), 
	.B1(U_addrdec_n67), 
	.A(U_addrdec_n74));
   OAI21_X1 U102 (.ZN(n73), 
	.B2(U_dsdc_n1948), 
	.B1(U_dsdc_bm_bank_age_0__1_), 
	.A(U_dsdc_n1947));
   OAI21_X1 U103 (.ZN(n74), 
	.B2(U_dsdc_n334), 
	.B1(U_dsdc_n1951), 
	.A(n73));
   AOI222_X1 U104 (.ZN(n75), 
	.C2(n74), 
	.C1(U_dsdc_n1953), 
	.B2(n74), 
	.B1(U_dsdc_bm_bank_age_0__3_), 
	.A2(U_dsdc_n1953), 
	.A1(U_dsdc_bm_bank_age_0__3_));
   AOI222_X1 U105 (.ZN(U_dsdc_n2080), 
	.C2(n75), 
	.C1(U_dsdc_n434), 
	.B2(n75), 
	.B1(U_dsdc_n1954), 
	.A2(U_dsdc_n434), 
	.A1(U_dsdc_n1954));
   OR2_X1 U106 (.ZN(n76), 
	.A2(U_dsdc_n1359), 
	.A1(U_dsdc_n1805));
   NAND4_X1 U107 (.ZN(n89), 
	.A4(n76), 
	.A3(U_dsdc_n1368), 
	.A2(U_dsdc_n1978), 
	.A1(U_dsdc_n1342));
   NAND3_X1 U108 (.ZN(n77), 
	.A3(FE_PHN3309_U_dsdc_cas_latency_cnt_2_), 
	.A2(U_dsdc_n1087), 
	.A1(U_dsdc_n1393));
   NAND2_X1 U110 (.ZN(n79), 
	.A2(n67), 
	.A1(U_dsdc_cas_latency_2_));
   OAI211_X1 U111 (.ZN(U_dsdc_N4128), 
	.C2(U_dsdc_n1090), 
	.C1(FE_PHN1585_U_dsdc_n1094), 
	.B(n79), 
	.A(n77));
   OAI21_X1 U112 (.ZN(n80), 
	.B2(U_dmc_n61), 
	.B1(U_dmc_n5), 
	.A(U_dmc_n60));
   NOR2_X1 U113 (.ZN(n81), 
	.A2(n80), 
	.A1(ctl_burst_done));
   OAI211_X1 U114 (.ZN(miu_burst_done), 
	.C2(U_cr_n502), 
	.C1(U_cr_n503), 
	.B(n81), 
	.A(FE_PHN1400_U_cr_n197));
   OAI21_X2 U115 (.ZN(U_dsdc_n1025), 
	.B2(U_dsdc_n1023), 
	.B1(U_dsdc_n1024), 
	.A(U_dsdc_bm_num_open_bank_4_));
   AOI21_X2 U116 (.ZN(U_dsdc_n561), 
	.B2(U_dsdc_bm_row_addr_2__0_), 
	.B1(U_dsdc_n159), 
	.A(U_dsdc_n560));
   OAI211_X2 U117 (.ZN(debug_ad_bank_addr[0]), 
	.C2(FE_PHN1645_U_cr_n65), 
	.C1(U_addrdec_n73), 
	.B(U_addrdec_n70), 
	.A(U_addrdec_n71));
   NAND2_X1 U118 (.ZN(U_dsdc_n913), 
	.A2(U_dsdc_n979), 
	.A1(U_dsdc_n981));
   NAND2_X1 U119 (.ZN(U_dsdc_n987), 
	.A2(debug_ad_bank_addr[0]), 
	.A1(debug_ad_bank_addr[1]));
   AOI22_X1 U120 (.ZN(U_addrdec_n96), 
	.B2(U_addrdec_n39), 
	.B1(hiu_addr[1]), 
	.A2(hiu_addr[2]), 
	.A1(U_addrdec_n220));
   AOI22_X1 U121 (.ZN(U_addrdec_n97), 
	.B2(U_addrdec_n39), 
	.B1(hiu_addr[4]), 
	.A2(hiu_addr[5]), 
	.A1(U_addrdec_n220));
   AOI22_X1 U122 (.ZN(U_addrdec_n99), 
	.B2(U_addrdec_n39), 
	.B1(hiu_addr[6]), 
	.A2(hiu_addr[7]), 
	.A1(U_addrdec_n220));
   AOI22_X1 U123 (.ZN(U_addrdec_n98), 
	.B2(U_addrdec_n39), 
	.B1(hiu_addr[5]), 
	.A2(hiu_addr[6]), 
	.A1(U_addrdec_n220));
   NOR2_X2 U124 (.ZN(U_dsdc_n538), 
	.A2(U_dsdc_n333), 
	.A1(U_dsdc_n537));
   OAI211_X2 U125 (.ZN(U_addrdec_n85), 
	.C2(U_addrdec_n84), 
	.C1(n[24]), 
	.B(U_addrdec_n82), 
	.A(U_addrdec_n83));
   INV_X4 U126 (.ZN(debug_ad_bank_addr[1]), 
	.A(n14));
   INV_X4 U128 (.ZN(U_addrdec_n40), 
	.A(big_endian));
   NAND2_X4 U129 (.ZN(n83), 
	.A2(U_dsdc_n998), 
	.A1(U_dsdc_n1166));
   INV_X4 U130 (.ZN(U_dsdc_DP_OP_1642_126_2028_n85), 
	.A(U_dsdc_n601));
   AND2_X4 U131 (.ZN(n86), 
	.A2(U_dsdc_n604), 
	.A1(U_dsdc_bm_row_addr_1__8_));
endmodule

module DW_memctl (
	hready_resp, 
	hresp, 
	hrdata, 
	s_ras_n, 
	s_cas_n, 
	s_cke, 
	s_wr_data, 
	s_addr, 
	s_bank_addr, 
	s_dout_valid, 
	s_sel_n, 
	s_dqm, 
	s_we_n, 
	s_dqs, 
	s_sa, 
	s_scl, 
	s_rd_ready, 
	s_rd_start, 
	s_rd_pop, 
	s_rd_end, 
	s_rd_dqs_mask, 
	s_cas_latency, 
	s_read_pipe, 
	s_sda_out, 
	s_sda_oe_n, 
	gpo, 
	debug_ad_bank_addr, 
	debug_ad_row_addr, 
	debug_ad_col_addr, 
	debug_ad_sf_bank_addr, 
	debug_ad_sf_row_addr, 
	debug_ad_sf_col_addr, 
	debug_hiu_addr, 
	debug_sm_burst_done, 
	debug_sm_pop_n, 
	debug_sm_push_n, 
	debug_smc_cs, 
	debug_ref_req, 
	hclk, 
	hclk_2x, 
	hresetn, 
	scan_mode, 
	haddr, 
	hsel_mem, 
	hsel_reg, 
	hwrite, 
	htrans, 
	hsize, 
	hburst, 
	hready, 
	hwdata, 
	s_rd_data, 
	s_sda_in, 
	gpi, 
	remap, 
	power_down, 
	clear_sr_dp, 
	big_endian, 
	FE_OFN28_HRESETn, 
	FE_OFN29_HRESETn, 
	FE_OFN30_HRESETn, 
	FE_OFN34_HRESETn, 
	FE_OFN42_HRESETn, 
	FE_OFN43_HRESETn, 
	FE_OFN55_HRESETn, 
	HCLK__L5_N11, 
	HCLK__L5_N12, 
	HCLK__L5_N13, 
	HCLK__L5_N14, 
	HCLK__L5_N15, 
	HCLK__L5_N16, 
	HCLK__L5_N17, 
	HCLK__L5_N18, 
	HCLK__L5_N27, 
	HCLK__L5_N28, 
	HCLK__L5_N29, 
	HCLK__L5_N30, 
	HCLK__L5_N31, 
	HCLK__L5_N32, 
	HCLK__L5_N33, 
	HCLK__L5_N34, 
	HCLK__L5_N35, 
	HCLK__L5_N36, 
	HCLK__L5_N37, 
	HCLK__L5_N38, 
	HCLK__L5_N39, 
	HCLK__L5_N4, 
	HCLK__L5_N5, 
	HCLK__L5_N6);
   output hready_resp;
   output [1:0] hresp;
   output [31:0] hrdata;
   output s_ras_n;
   output s_cas_n;
   output s_cke;
   output [15:0] s_wr_data;
   output [15:0] s_addr;
   output [1:0] s_bank_addr;
   output [1:0] s_dout_valid;
   output [0:0] s_sel_n;
   output [1:0] s_dqm;
   output s_we_n;
   output [1:0] s_dqs;
   output [2:0] s_sa;
   output s_scl;
   input s_rd_ready;
   output s_rd_start;
   output s_rd_pop;
   output s_rd_end;
   output s_rd_dqs_mask;
   output [2:0] s_cas_latency;
   output [2:0] s_read_pipe;
   output s_sda_out;
   output s_sda_oe_n;
   output [7:0] gpo;
   output [1:0] debug_ad_bank_addr;
   output [15:0] debug_ad_row_addr;
   output [15:0] debug_ad_col_addr;
   output [1:0] debug_ad_sf_bank_addr;
   output [15:0] debug_ad_sf_row_addr;
   output [15:0] debug_ad_sf_col_addr;
   output [31:0] debug_hiu_addr;
   output debug_sm_burst_done;
   output debug_sm_pop_n;
   output debug_sm_push_n;
   output [3:0] debug_smc_cs;
   output debug_ref_req;
   input hclk;
   input hclk_2x;
   input hresetn;
   input scan_mode;
   input [31:0] haddr;
   input hsel_mem;
   input hsel_reg;
   input hwrite;
   input [1:0] htrans;
   input [2:0] hsize;
   input [2:0] hburst;
   input hready;
   input [31:0] hwdata;
   input [31:0] s_rd_data;
   input s_sda_in;
   input [7:0] gpi;
   input remap;
   input power_down;
   input clear_sr_dp;
   input big_endian;
   input FE_OFN28_HRESETn;
   input FE_OFN29_HRESETn;
   input FE_OFN30_HRESETn;
   input FE_OFN34_HRESETn;
   input FE_OFN42_HRESETn;
   input FE_OFN43_HRESETn;
   input FE_OFN55_HRESETn;
   input HCLK__L5_N11;
   input HCLK__L5_N12;
   input HCLK__L5_N13;
   input HCLK__L5_N14;
   input HCLK__L5_N15;
   input HCLK__L5_N16;
   input HCLK__L5_N17;
   input HCLK__L5_N18;
   input HCLK__L5_N27;
   input HCLK__L5_N28;
   input HCLK__L5_N29;
   input HCLK__L5_N30;
   input HCLK__L5_N31;
   input HCLK__L5_N32;
   input HCLK__L5_N33;
   input HCLK__L5_N34;
   input HCLK__L5_N35;
   input HCLK__L5_N36;
   input HCLK__L5_N37;
   input HCLK__L5_N38;
   input HCLK__L5_N39;
   input HCLK__L5_N4;
   input HCLK__L5_N5;
   input HCLK__L5_N6;

   // Internal wires
   wire FE_PHN5173_big_endian;
   wire FE_PHN4651_miu_data_25_;
   wire FE_PHN4648_miu_data_16_;
   wire FE_PHN4622_big_endian;
   wire FE_PHN3010_miu_data_21_;
   wire FE_PHN3009_miu_data_6_;
   wire FE_PHN2962_miu_data_26_;
   wire FE_PHN2961_miu_data_0_;
   wire FE_PHN2960_miu_data_22_;
   wire FE_PHN2959_miu_data_18_;
   wire FE_PHN2958_miu_data_19_;
   wire FE_PHN2956_miu_data_23_;
   wire FE_PHN2950_miu_data_12_;
   wire FE_PHN2932_miu_data_10_;
   wire FE_PHN2931_miu_data_3_;
   wire FE_PHN2925_miu_data_5_;
   wire FE_PHN2919_miu_data_9_;
   wire FE_PHN2907_big_endian;
   wire FE_PHN976_miu_data_25_;
   wire FE_PHN974_miu_data_28_;
   wire FE_PHN973_miu_data_31_;
   wire FE_PHN879_miu_data_9_;
   wire FE_PHN878_miu_data_1_;
   wire FE_PHN877_miu_data_6_;
   wire FE_PHN874_miu_data_0_;
   wire FE_PHN873_miu_data_3_;
   wire FE_PHN871_miu_data_7_;
   wire FE_PHN805_miu_data_22_;
   wire FE_PHN794_miu_data_23_;
   wire FE_PHN766_miu_data_18_;
   wire FE_PHN754_miu_data_16_;
   wire FE_PHN746_miu_data_26_;
   wire FE_PHN724_miu_data_21_;
   wire FE_PHN718_miu_data_12_;
   wire FE_PHN709_miu_data_19_;
   wire FE_PHN689_miu_data_20_;
   wire FE_PHN686_miu_data_5_;
   wire FE_PHN684_miu_data_17_;
   wire FE_PHN680_miu_data_24_;
   wire FE_PHN677_miu_data_10_;
   wire FE_PHN669_big_endian;
   wire FE_OFN191_HRESETn;
   wire FE_OFN160_HRESETn;
   wire FE_OFN151_HRESETn;
   wire FE_OFN57_HRESETn;
   wire FE_OFN53_HRESETn;
   wire FE_OFN51_HRESETn;
   wire FE_OFN46_HRESETn;
   wire FE_OFN35_HRESETn;
   wire FE_OFN31_HRESETn;
   wire hiu_wrap_burst;
   wire hiu_rw;
   wire hiu_terminate;
   wire miu_burst_done;
   wire miu_pop_n;
   wire miu_push_n;
   wire n2;
   wire SYNOPSYS_UNCONNECTED_1;
   wire SYNOPSYS_UNCONNECTED_2;
   wire SYNOPSYS_UNCONNECTED_3;
   wire SYNOPSYS_UNCONNECTED_4;
   wire SYNOPSYS_UNCONNECTED_5;
   wire SYNOPSYS_UNCONNECTED_6;
   wire SYNOPSYS_UNCONNECTED_7;
   wire SYNOPSYS_UNCONNECTED_8;
   wire SYNOPSYS_UNCONNECTED_9;
   wire SYNOPSYS_UNCONNECTED_10;
   wire SYNOPSYS_UNCONNECTED_11;
   wire SYNOPSYS_UNCONNECTED_12;
   wire SYNOPSYS_UNCONNECTED_13;
   wire SYNOPSYS_UNCONNECTED_14;
   wire SYNOPSYS_UNCONNECTED_15;
   wire SYNOPSYS_UNCONNECTED_16;
   wire SYNOPSYS_UNCONNECTED_17;
   wire SYNOPSYS_UNCONNECTED_18;
   wire SYNOPSYS_UNCONNECTED_19;
   wire SYNOPSYS_UNCONNECTED_20;
   wire SYNOPSYS_UNCONNECTED_21;
   wire SYNOPSYS_UNCONNECTED_22;
   wire SYNOPSYS_UNCONNECTED_23;
   wire SYNOPSYS_UNCONNECTED_24;
   wire SYNOPSYS_UNCONNECTED_25;
   wire SYNOPSYS_UNCONNECTED_26;
   wire SYNOPSYS_UNCONNECTED_27;
   wire SYNOPSYS_UNCONNECTED_28;
   wire SYNOPSYS_UNCONNECTED_29;
   wire SYNOPSYS_UNCONNECTED_30;
   wire SYNOPSYS_UNCONNECTED_31;
   wire SYNOPSYS_UNCONNECTED_32;
   wire SYNOPSYS_UNCONNECTED_33;
   wire SYNOPSYS_UNCONNECTED_34;
   wire SYNOPSYS_UNCONNECTED_35;
   wire SYNOPSYS_UNCONNECTED_36;
   wire SYNOPSYS_UNCONNECTED_37;
   wire SYNOPSYS_UNCONNECTED_38;
   wire SYNOPSYS_UNCONNECTED_39;
   wire SYNOPSYS_UNCONNECTED_40;
   wire SYNOPSYS_UNCONNECTED_41;
   wire SYNOPSYS_UNCONNECTED_42;
   wire SYNOPSYS_UNCONNECTED_43;
   wire SYNOPSYS_UNCONNECTED_44;
   wire SYNOPSYS_UNCONNECTED_45;
   wire SYNOPSYS_UNCONNECTED_46;
   wire SYNOPSYS_UNCONNECTED_47;
   wire SYNOPSYS_UNCONNECTED_48;
   wire SYNOPSYS_UNCONNECTED_49;
   wire SYNOPSYS_UNCONNECTED_50;
   wire SYNOPSYS_UNCONNECTED_51;
   wire SYNOPSYS_UNCONNECTED_52;
   wire SYNOPSYS_UNCONNECTED_53;
   wire SYNOPSYS_UNCONNECTED_54;
   wire SYNOPSYS_UNCONNECTED_55;
   wire SYNOPSYS_UNCONNECTED_56;
   wire SYNOPSYS_UNCONNECTED_57;
   wire SYNOPSYS_UNCONNECTED_58;
   wire SYNOPSYS_UNCONNECTED_59;
   wire SYNOPSYS_UNCONNECTED_60;
   wire SYNOPSYS_UNCONNECTED_61;
   wire SYNOPSYS_UNCONNECTED_62;
   wire SYNOPSYS_UNCONNECTED_63;
   wire SYNOPSYS_UNCONNECTED_64;
   wire SYNOPSYS_UNCONNECTED_65;
   wire SYNOPSYS_UNCONNECTED_66;
   wire SYNOPSYS_UNCONNECTED_67;
   wire SYNOPSYS_UNCONNECTED_68;
   wire SYNOPSYS_UNCONNECTED_69;
   wire SYNOPSYS_UNCONNECTED_70;
   wire SYNOPSYS_UNCONNECTED_71;
   wire SYNOPSYS_UNCONNECTED_72;
   wire SYNOPSYS_UNCONNECTED_73;
   wire SYNOPSYS_UNCONNECTED_74;
   wire SYNOPSYS_UNCONNECTED_75;
   wire SYNOPSYS_UNCONNECTED_76;
   wire SYNOPSYS_UNCONNECTED_77;
   wire SYNOPSYS_UNCONNECTED_78;
   wire SYNOPSYS_UNCONNECTED_79;
   wire SYNOPSYS_UNCONNECTED_80;
   wire SYNOPSYS_UNCONNECTED_81;
   wire SYNOPSYS_UNCONNECTED_82;
   wire SYNOPSYS_UNCONNECTED_83;
   wire SYNOPSYS_UNCONNECTED_84;
   wire SYNOPSYS_UNCONNECTED_85;
   wire SYNOPSYS_UNCONNECTED_86;
   wire SYNOPSYS_UNCONNECTED_87;
   wire SYNOPSYS_UNCONNECTED_88;
   wire SYNOPSYS_UNCONNECTED_89;
   wire SYNOPSYS_UNCONNECTED_90;
   wire SYNOPSYS_UNCONNECTED_91;
   wire SYNOPSYS_UNCONNECTED_92;
   wire SYNOPSYS_UNCONNECTED_93;
   wire SYNOPSYS_UNCONNECTED_94;
   wire SYNOPSYS_UNCONNECTED_95;
   wire SYNOPSYS_UNCONNECTED_96;
   wire SYNOPSYS_UNCONNECTED_97;
   wire SYNOPSYS_UNCONNECTED_98;
   wire SYNOPSYS_UNCONNECTED_99;
   wire SYNOPSYS_UNCONNECTED_100;
   wire SYNOPSYS_UNCONNECTED_101;
   wire SYNOPSYS_UNCONNECTED_102;
   wire SYNOPSYS_UNCONNECTED_103;
   wire SYNOPSYS_UNCONNECTED_104;
   wire SYNOPSYS_UNCONNECTED_105;
   wire SYNOPSYS_UNCONNECTED_106;
   wire SYNOPSYS_UNCONNECTED_107;
   wire SYNOPSYS_UNCONNECTED_108;
   wire SYNOPSYS_UNCONNECTED_109;
   wire SYNOPSYS_UNCONNECTED_110;
   wire SYNOPSYS_UNCONNECTED_111;
   wire SYNOPSYS_UNCONNECTED_112;
   wire SYNOPSYS_UNCONNECTED_113;
   wire SYNOPSYS_UNCONNECTED_114;
   wire SYNOPSYS_UNCONNECTED_115;
   wire SYNOPSYS_UNCONNECTED_116;
   wire SYNOPSYS_UNCONNECTED_117;
   wire SYNOPSYS_UNCONNECTED_118;
   wire SYNOPSYS_UNCONNECTED_119;
   wire SYNOPSYS_UNCONNECTED_120;
   wire SYNOPSYS_UNCONNECTED_121;
   wire SYNOPSYS_UNCONNECTED_122;
   wire SYNOPSYS_UNCONNECTED_123;
   wire SYNOPSYS_UNCONNECTED_124;
   wire SYNOPSYS_UNCONNECTED_125;
   wire SYNOPSYS_UNCONNECTED_126;
   wire SYNOPSYS_UNCONNECTED_127;
   wire SYNOPSYS_UNCONNECTED_128;
   wire SYNOPSYS_UNCONNECTED_129;
   wire SYNOPSYS_UNCONNECTED_130;
   wire SYNOPSYS_UNCONNECTED_131;
   wire SYNOPSYS_UNCONNECTED_132;
   wire SYNOPSYS_UNCONNECTED_133;
   wire SYNOPSYS_UNCONNECTED_134;
   wire SYNOPSYS_UNCONNECTED_135;
   wire SYNOPSYS_UNCONNECTED_136;
   wire SYNOPSYS_UNCONNECTED_137;
   wire SYNOPSYS_UNCONNECTED_138;
   wire SYNOPSYS_UNCONNECTED_139;
   wire SYNOPSYS_UNCONNECTED_140;
   wire SYNOPSYS_UNCONNECTED_141;
   wire SYNOPSYS_UNCONNECTED_142;
   wire SYNOPSYS_UNCONNECTED_143;
   wire SYNOPSYS_UNCONNECTED_144;
   wire SYNOPSYS_UNCONNECTED_145;
   wire SYNOPSYS_UNCONNECTED_146;
   wire SYNOPSYS_UNCONNECTED_147;
   wire SYNOPSYS_UNCONNECTED_148;
   wire SYNOPSYS_UNCONNECTED_149;
   wire SYNOPSYS_UNCONNECTED_150;
   wire [1:0] hiu_req;
   wire [5:0] hiu_burst_size;
   wire [31:0] hiu_data;
   wire [3:0] hiu_haddr;
   wire [2:0] hiu_hsize;
   wire [31:0] miu_data;

   assign debug_smc_cs[0] = 1'b0 ;
   assign debug_smc_cs[1] = 1'b0 ;
   assign debug_smc_cs[2] = 1'b0 ;
   assign debug_smc_cs[3] = 1'b0 ;
   assign debug_sm_push_n = 1'b0 ;
   assign debug_sm_pop_n = 1'b0 ;
   assign debug_sm_burst_done = 1'b0 ;
   assign debug_hiu_addr[0] = 1'b0 ;
   assign debug_ad_sf_col_addr[0] = 1'b0 ;
   assign debug_ad_sf_col_addr[1] = 1'b0 ;
   assign debug_ad_sf_col_addr[2] = 1'b0 ;
   assign debug_ad_sf_col_addr[3] = 1'b0 ;
   assign debug_ad_sf_col_addr[4] = 1'b0 ;
   assign debug_ad_sf_col_addr[5] = 1'b0 ;
   assign debug_ad_sf_col_addr[6] = 1'b0 ;
   assign debug_ad_sf_col_addr[7] = 1'b0 ;
   assign debug_ad_sf_col_addr[8] = 1'b0 ;
   assign debug_ad_sf_col_addr[9] = 1'b0 ;
   assign debug_ad_sf_col_addr[10] = 1'b0 ;
   assign debug_ad_sf_col_addr[11] = 1'b0 ;
   assign debug_ad_sf_col_addr[12] = 1'b0 ;
   assign debug_ad_sf_col_addr[13] = 1'b0 ;
   assign debug_ad_sf_col_addr[14] = 1'b0 ;
   assign debug_ad_sf_col_addr[15] = 1'b0 ;
   assign debug_ad_sf_row_addr[0] = 1'b0 ;
   assign debug_ad_sf_row_addr[1] = 1'b0 ;
   assign debug_ad_sf_row_addr[2] = 1'b0 ;
   assign debug_ad_sf_row_addr[3] = 1'b0 ;
   assign debug_ad_sf_row_addr[4] = 1'b0 ;
   assign debug_ad_sf_row_addr[5] = 1'b0 ;
   assign debug_ad_sf_row_addr[6] = 1'b0 ;
   assign debug_ad_sf_row_addr[7] = 1'b0 ;
   assign debug_ad_sf_row_addr[8] = 1'b0 ;
   assign debug_ad_sf_row_addr[9] = 1'b0 ;
   assign debug_ad_sf_row_addr[10] = 1'b0 ;
   assign debug_ad_sf_row_addr[11] = 1'b0 ;
   assign debug_ad_sf_row_addr[12] = 1'b0 ;
   assign debug_ad_sf_row_addr[13] = 1'b0 ;
   assign debug_ad_sf_row_addr[14] = 1'b0 ;
   assign debug_ad_sf_row_addr[15] = 1'b0 ;
   assign debug_ad_sf_bank_addr[0] = 1'b0 ;
   assign debug_ad_sf_bank_addr[1] = 1'b0 ;
   assign hresp[0] = 1'b0 ;
   assign hresp[1] = 1'b0 ;

   CLKBUF_X3 FE_PHC5173_big_endian (.Z(FE_PHN5173_big_endian), 
	.A(FE_PHN4622_big_endian));
   BUF_X8 FE_PHC4651_miu_data_25_ (.Z(FE_PHN4651_miu_data_25_), 
	.A(miu_data[25]));
   BUF_X16 FE_PHC4648_miu_data_16_ (.Z(FE_PHN4648_miu_data_16_), 
	.A(miu_data[16]));
   BUF_X32 FE_PHC4622_big_endian (.Z(FE_PHN4622_big_endian), 
	.A(FE_PHN2907_big_endian));
   BUF_X32 FE_PHC3010_miu_data_21_ (.Z(FE_PHN3010_miu_data_21_), 
	.A(miu_data[21]));
   BUF_X32 FE_PHC3009_miu_data_6_ (.Z(FE_PHN3009_miu_data_6_), 
	.A(miu_data[6]));
   BUF_X32 FE_PHC2962_miu_data_26_ (.Z(FE_PHN2962_miu_data_26_), 
	.A(miu_data[26]));
   BUF_X32 FE_PHC2961_miu_data_0_ (.Z(FE_PHN2961_miu_data_0_), 
	.A(miu_data[0]));
   BUF_X32 FE_PHC2960_miu_data_22_ (.Z(FE_PHN2960_miu_data_22_), 
	.A(miu_data[22]));
   BUF_X32 FE_PHC2959_miu_data_18_ (.Z(FE_PHN2959_miu_data_18_), 
	.A(miu_data[18]));
   BUF_X32 FE_PHC2958_miu_data_19_ (.Z(FE_PHN2958_miu_data_19_), 
	.A(miu_data[19]));
   BUF_X32 FE_PHC2956_miu_data_23_ (.Z(FE_PHN2956_miu_data_23_), 
	.A(miu_data[23]));
   BUF_X32 FE_PHC2950_miu_data_12_ (.Z(FE_PHN2950_miu_data_12_), 
	.A(miu_data[12]));
   BUF_X32 FE_PHC2932_miu_data_10_ (.Z(FE_PHN2932_miu_data_10_), 
	.A(miu_data[10]));
   BUF_X32 FE_PHC2931_miu_data_3_ (.Z(FE_PHN2931_miu_data_3_), 
	.A(miu_data[3]));
   BUF_X32 FE_PHC2925_miu_data_5_ (.Z(FE_PHN2925_miu_data_5_), 
	.A(miu_data[5]));
   BUF_X32 FE_PHC2919_miu_data_9_ (.Z(FE_PHN2919_miu_data_9_), 
	.A(miu_data[9]));
   CLKBUF_X3 FE_PHC2907_big_endian (.Z(FE_PHN2907_big_endian), 
	.A(FE_PHN669_big_endian));
   BUF_X32 FE_PHC976_miu_data_25_ (.Z(FE_PHN976_miu_data_25_), 
	.A(FE_PHN4651_miu_data_25_));
   BUF_X32 FE_PHC974_miu_data_28_ (.Z(FE_PHN974_miu_data_28_), 
	.A(miu_data[28]));
   BUF_X32 FE_PHC973_miu_data_31_ (.Z(FE_PHN973_miu_data_31_), 
	.A(miu_data[31]));
   BUF_X32 FE_PHC879_miu_data_9_ (.Z(FE_PHN879_miu_data_9_), 
	.A(FE_PHN2919_miu_data_9_));
   BUF_X32 FE_PHC878_miu_data_1_ (.Z(FE_PHN878_miu_data_1_), 
	.A(miu_data[1]));
   BUF_X32 FE_PHC877_miu_data_6_ (.Z(FE_PHN877_miu_data_6_), 
	.A(FE_PHN3009_miu_data_6_));
   BUF_X32 FE_PHC874_miu_data_0_ (.Z(FE_PHN874_miu_data_0_), 
	.A(FE_PHN2961_miu_data_0_));
   BUF_X32 FE_PHC873_miu_data_3_ (.Z(FE_PHN873_miu_data_3_), 
	.A(FE_PHN2931_miu_data_3_));
   BUF_X32 FE_PHC871_miu_data_7_ (.Z(FE_PHN871_miu_data_7_), 
	.A(miu_data[7]));
   BUF_X32 FE_PHC805_miu_data_22_ (.Z(FE_PHN805_miu_data_22_), 
	.A(FE_PHN2960_miu_data_22_));
   BUF_X32 FE_PHC794_miu_data_23_ (.Z(FE_PHN794_miu_data_23_), 
	.A(FE_PHN2956_miu_data_23_));
   BUF_X32 FE_PHC766_miu_data_18_ (.Z(FE_PHN766_miu_data_18_), 
	.A(FE_PHN2959_miu_data_18_));
   BUF_X32 FE_PHC754_miu_data_16_ (.Z(FE_PHN754_miu_data_16_), 
	.A(FE_PHN4648_miu_data_16_));
   BUF_X32 FE_PHC746_miu_data_26_ (.Z(FE_PHN746_miu_data_26_), 
	.A(FE_PHN2962_miu_data_26_));
   BUF_X32 FE_PHC724_miu_data_21_ (.Z(FE_PHN724_miu_data_21_), 
	.A(FE_PHN3010_miu_data_21_));
   BUF_X32 FE_PHC718_miu_data_12_ (.Z(FE_PHN718_miu_data_12_), 
	.A(FE_PHN2950_miu_data_12_));
   BUF_X32 FE_PHC709_miu_data_19_ (.Z(FE_PHN709_miu_data_19_), 
	.A(FE_PHN2958_miu_data_19_));
   BUF_X32 FE_PHC689_miu_data_20_ (.Z(FE_PHN689_miu_data_20_), 
	.A(miu_data[20]));
   BUF_X32 FE_PHC686_miu_data_5_ (.Z(FE_PHN686_miu_data_5_), 
	.A(FE_PHN2925_miu_data_5_));
   BUF_X32 FE_PHC684_miu_data_17_ (.Z(FE_PHN684_miu_data_17_), 
	.A(miu_data[17]));
   BUF_X32 FE_PHC680_miu_data_24_ (.Z(FE_PHN680_miu_data_24_), 
	.A(miu_data[24]));
   BUF_X32 FE_PHC677_miu_data_10_ (.Z(FE_PHN677_miu_data_10_), 
	.A(FE_PHN2932_miu_data_10_));
   CLKBUF_X3 FE_PHC669_big_endian (.Z(FE_PHN669_big_endian), 
	.A(big_endian));
   BUF_X4 FE_OFC191_HRESETn (.Z(FE_OFN191_HRESETn), 
	.A(FE_OFN31_HRESETn));
   BUF_X4 FE_OFC160_HRESETn (.Z(FE_OFN160_HRESETn), 
	.A(FE_OFN51_HRESETn));
   BUF_X4 FE_OFC151_HRESETn (.Z(FE_OFN151_HRESETn), 
	.A(FE_OFN57_HRESETn));
   BUF_X8 FE_OFC57_HRESETn (.Z(FE_OFN57_HRESETn), 
	.A(FE_OFN35_HRESETn));
   BUF_X8 FE_OFC53_HRESETn (.Z(FE_OFN53_HRESETn), 
	.A(FE_OFN28_HRESETn));
   BUF_X8 FE_OFC51_HRESETn (.Z(FE_OFN51_HRESETn), 
	.A(FE_OFN30_HRESETn));
   BUF_X8 FE_OFC46_HRESETn (.Z(FE_OFN46_HRESETn), 
	.A(FE_OFN31_HRESETn));
   INV_X8 FE_OFC35_HRESETn (.ZN(FE_OFN35_HRESETn), 
	.A(hresetn));
   INV_X8 FE_OFC31_HRESETn (.ZN(FE_OFN31_HRESETn), 
	.A(hresetn));
   DW_memctl_hiu U_hiu (.hclk(HCLK__L5_N13), 
	.hresetn(hresetn), 
	.hsel_mem(hsel_mem), 
	.hsel_reg(hsel_reg), 
	.htrans(htrans), 
	.hwrite(hwrite), 
	.hsize(hsize), 
	.hburst(hburst), 
	.hready(hready), 
	.hready_resp(hready_resp), 
	.hresp({ SYNOPSYS_UNCONNECTED_1,
		SYNOPSYS_UNCONNECTED_2 }), 
	.haddr(haddr), 
	.hwdata(hwdata), 
	.hrdata(hrdata), 
	.hiu_req(hiu_req), 
	.hiu_burst_size(hiu_burst_size), 
	.hiu_wrap_burst(hiu_wrap_burst), 
	.hiu_rw(hiu_rw), 
	.hiu_terminate(hiu_terminate), 
	.hiu_addr({ debug_hiu_addr[31],
		debug_hiu_addr[30],
		debug_hiu_addr[29],
		debug_hiu_addr[28],
		debug_hiu_addr[27],
		debug_hiu_addr[26],
		debug_hiu_addr[25],
		debug_hiu_addr[24],
		debug_hiu_addr[23],
		debug_hiu_addr[22],
		debug_hiu_addr[21],
		debug_hiu_addr[20],
		debug_hiu_addr[19],
		debug_hiu_addr[18],
		debug_hiu_addr[17],
		debug_hiu_addr[16],
		debug_hiu_addr[15],
		debug_hiu_addr[14],
		debug_hiu_addr[13],
		debug_hiu_addr[12],
		debug_hiu_addr[11],
		debug_hiu_addr[10],
		debug_hiu_addr[9],
		debug_hiu_addr[8],
		debug_hiu_addr[7],
		debug_hiu_addr[6],
		debug_hiu_addr[5],
		debug_hiu_addr[4],
		debug_hiu_addr[3],
		debug_hiu_addr[2],
		debug_hiu_addr[1],
		SYNOPSYS_UNCONNECTED_3 }), 
	.hiu_data(hiu_data), 
	.hiu_haddr(hiu_haddr), 
	.hiu_hsize(hiu_hsize), 
	.miu_burst_done(miu_burst_done), 
	.miu_push_n(miu_push_n), 
	.miu_pop_n(miu_pop_n), 
	.miu_data({ FE_PHN973_miu_data_31_,
		miu_data[30],
		miu_data[29],
		FE_PHN974_miu_data_28_,
		miu_data[27],
		FE_PHN746_miu_data_26_,
		FE_PHN976_miu_data_25_,
		FE_PHN680_miu_data_24_,
		FE_PHN794_miu_data_23_,
		FE_PHN805_miu_data_22_,
		FE_PHN724_miu_data_21_,
		FE_PHN689_miu_data_20_,
		FE_PHN709_miu_data_19_,
		FE_PHN766_miu_data_18_,
		FE_PHN684_miu_data_17_,
		FE_PHN754_miu_data_16_,
		miu_data[15],
		miu_data[14],
		n2,
		FE_PHN718_miu_data_12_,
		miu_data[11],
		FE_PHN677_miu_data_10_,
		FE_PHN879_miu_data_9_,
		miu_data[8],
		FE_PHN871_miu_data_7_,
		FE_PHN877_miu_data_6_,
		FE_PHN686_miu_data_5_,
		miu_data[4],
		FE_PHN873_miu_data_3_,
		miu_data[2],
		FE_PHN878_miu_data_1_,
		FE_PHN874_miu_data_0_ }), 
	.miu_data_width({ 1'b0,
		1'b0 }), 
	.miu_col_width({ 1'b0,
		1'b0,
		1'b0,
		1'b0 }), 
	.big_endian(FE_PHN5173_big_endian), 
	.FE_OFN28_HRESETn(FE_OFN28_HRESETn), 
	.FE_OFN29_HRESETn(FE_OFN29_HRESETn), 
	.FE_OFN30_HRESETn(FE_OFN30_HRESETn), 
	.FE_OFN34_HRESETn(FE_OFN34_HRESETn), 
	.FE_OFN42_HRESETn(FE_OFN42_HRESETn), 
	.FE_OFN43_HRESETn(FE_OFN43_HRESETn), 
	.FE_OFN55_HRESETn(FE_OFN55_HRESETn), 
	.FE_OFN31_HRESETn(FE_OFN31_HRESETn), 
	.FE_OFN35_HRESETn(FE_OFN35_HRESETn), 
	.FE_OFN46_HRESETn(FE_OFN46_HRESETn), 
	.FE_OFN51_HRESETn(FE_OFN51_HRESETn), 
	.FE_OFN53_HRESETn(FE_OFN53_HRESETn), 
	.FE_OFN57_HRESETn(FE_OFN57_HRESETn), 
	.HCLK__L5_N14(HCLK__L5_N14), 
	.HCLK__L5_N15(HCLK__L5_N15), 
	.HCLK__L5_N16(HCLK__L5_N16), 
	.HCLK__L5_N17(HCLK__L5_N17), 
	.HCLK__L5_N18(HCLK__L5_N18), 
	.HCLK__L5_N27(HCLK__L5_N27), 
	.HCLK__L5_N32(HCLK__L5_N32), 
	.HCLK__L5_N33(HCLK__L5_N33), 
	.HCLK__L5_N34(HCLK__L5_N34), 
	.HCLK__L5_N35(HCLK__L5_N35), 
	.HCLK__L5_N36(HCLK__L5_N36), 
	.HCLK__L5_N37(HCLK__L5_N37), 
	.HCLK__L5_N38(HCLK__L5_N38), 
	.HCLK__L5_N39(HCLK__L5_N39), 
	.HCLK__L5_N4(HCLK__L5_N4), 
	.HCLK__L5_N5(HCLK__L5_N5), 
	.HCLK__L5_N6(HCLK__L5_N6), 
	.FE_OFN151_HRESETn(FE_OFN151_HRESETn), 
	.FE_OFN160_HRESETn(FE_OFN160_HRESETn), 
	.FE_OFN191_HRESETn(FE_OFN191_HRESETn), 
	.FE_OFN214_hiu_burst_size_4_(hiu_burst_size[4]), 
	.FE_OFN217_hiu_burst_size_2_(hiu_burst_size[2]), 
	.FE_OFN220_hiu_burst_size_0_(hiu_burst_size[0]));
   DW_memctl_miu U_miu (.hclk(hclk), 
	.hclk_2x(hclk_2x), 
	.hresetn(hresetn), 
	.scan_mode(scan_mode), 
	.hiu_mem_req(hiu_req[1]), 
	.hiu_reg_req(hiu_req[0]), 
	.hiu_rw(hiu_rw), 
	.hiu_burst_size(hiu_burst_size), 
	.hiu_wrapped_burst(hiu_wrap_burst), 
	.hiu_terminate(hiu_terminate), 
	.hiu_addr({ debug_hiu_addr[31],
		debug_hiu_addr[30],
		debug_hiu_addr[29],
		debug_hiu_addr[28],
		debug_hiu_addr[27],
		debug_hiu_addr[26],
		debug_hiu_addr[25],
		debug_hiu_addr[24],
		debug_hiu_addr[23],
		debug_hiu_addr[22],
		debug_hiu_addr[21],
		debug_hiu_addr[20],
		debug_hiu_addr[19],
		debug_hiu_addr[18],
		debug_hiu_addr[17],
		debug_hiu_addr[16],
		debug_hiu_addr[15],
		debug_hiu_addr[14],
		debug_hiu_addr[13],
		debug_hiu_addr[12],
		debug_hiu_addr[11],
		debug_hiu_addr[10],
		debug_hiu_addr[9],
		debug_hiu_addr[8],
		debug_hiu_addr[7],
		debug_hiu_addr[6],
		debug_hiu_addr[5],
		debug_hiu_addr[4],
		debug_hiu_addr[3],
		debug_hiu_addr[2],
		debug_hiu_addr[1],
		1'b0 }), 
	.hiu_haddr(hiu_haddr), 
	.hiu_hsize(hiu_hsize), 
	.hiu_wr_data(hiu_data), 
	.s_rd_data(s_rd_data), 
	.miu_burst_done(miu_burst_done), 
	.miu_pop_n(miu_pop_n), 
	.miu_push_n(miu_push_n), 
	.miu_col_addr_width({ SYNOPSYS_UNCONNECTED_4,
		SYNOPSYS_UNCONNECTED_5,
		SYNOPSYS_UNCONNECTED_6,
		SYNOPSYS_UNCONNECTED_7 }), 
	.miu_data_width({ SYNOPSYS_UNCONNECTED_8,
		SYNOPSYS_UNCONNECTED_9 }), 
	.m_addr({ SYNOPSYS_UNCONNECTED_10,
		SYNOPSYS_UNCONNECTED_11,
		SYNOPSYS_UNCONNECTED_12,
		SYNOPSYS_UNCONNECTED_13,
		SYNOPSYS_UNCONNECTED_14,
		SYNOPSYS_UNCONNECTED_15,
		SYNOPSYS_UNCONNECTED_16,
		SYNOPSYS_UNCONNECTED_17,
		SYNOPSYS_UNCONNECTED_18,
		SYNOPSYS_UNCONNECTED_19,
		SYNOPSYS_UNCONNECTED_20,
		SYNOPSYS_UNCONNECTED_21,
		SYNOPSYS_UNCONNECTED_22,
		SYNOPSYS_UNCONNECTED_23,
		SYNOPSYS_UNCONNECTED_24,
		SYNOPSYS_UNCONNECTED_25 }), 
	.s_addr(s_addr), 
	.s_bank_addr(s_bank_addr), 
	.s_ras_n(s_ras_n), 
	.s_cas_n(s_cas_n), 
	.s_sel_n(s_sel_n), 
	.s_cke(s_cke), 
	.s_we_n(s_we_n), 
	.s_wr_data(s_wr_data), 
	.s_dqm(s_dqm), 
	.s_dout_valid(s_dout_valid), 
	.s_rd_ready(s_rd_ready), 
	.s_rd_start(s_rd_start), 
	.s_rd_pop(s_rd_pop), 
	.s_rd_end(s_rd_end), 
	.s_rd_dqs_mask(s_rd_dqs_mask), 
	.s_cas_latency(s_cas_latency), 
	.s_read_pipe(s_read_pipe), 
	.sf_cas_latency({ SYNOPSYS_UNCONNECTED_26,
		SYNOPSYS_UNCONNECTED_27,
		SYNOPSYS_UNCONNECTED_28 }), 
	.s_sa(s_sa), 
	.s_scl(s_scl), 
	.s_dqs(s_dqs), 
	.s_sda_out(s_sda_out), 
	.s_sda_in(s_sda_in), 
	.s_sda_oe_n(s_sda_oe_n), 
	.sm_addr({ SYNOPSYS_UNCONNECTED_29,
		SYNOPSYS_UNCONNECTED_30,
		SYNOPSYS_UNCONNECTED_31,
		SYNOPSYS_UNCONNECTED_32,
		SYNOPSYS_UNCONNECTED_33,
		SYNOPSYS_UNCONNECTED_34,
		SYNOPSYS_UNCONNECTED_35,
		SYNOPSYS_UNCONNECTED_36,
		SYNOPSYS_UNCONNECTED_37,
		SYNOPSYS_UNCONNECTED_38,
		SYNOPSYS_UNCONNECTED_39,
		SYNOPSYS_UNCONNECTED_40,
		SYNOPSYS_UNCONNECTED_41,
		SYNOPSYS_UNCONNECTED_42,
		SYNOPSYS_UNCONNECTED_43,
		SYNOPSYS_UNCONNECTED_44,
		SYNOPSYS_UNCONNECTED_45,
		SYNOPSYS_UNCONNECTED_46,
		SYNOPSYS_UNCONNECTED_47,
		SYNOPSYS_UNCONNECTED_48,
		SYNOPSYS_UNCONNECTED_49,
		SYNOPSYS_UNCONNECTED_50,
		SYNOPSYS_UNCONNECTED_51 }), 
	.sm_bs_n({ SYNOPSYS_UNCONNECTED_52,
		SYNOPSYS_UNCONNECTED_53,
		SYNOPSYS_UNCONNECTED_54,
		SYNOPSYS_UNCONNECTED_55 }), 
	.sm_dout_valid({ SYNOPSYS_UNCONNECTED_56,
		SYNOPSYS_UNCONNECTED_57,
		SYNOPSYS_UNCONNECTED_58,
		SYNOPSYS_UNCONNECTED_59 }), 
	.sm_wp_n({ SYNOPSYS_UNCONNECTED_60,
		SYNOPSYS_UNCONNECTED_61,
		SYNOPSYS_UNCONNECTED_62 }), 
	.sm_rd_data({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }), 
	.sm_wr_data({ SYNOPSYS_UNCONNECTED_63,
		SYNOPSYS_UNCONNECTED_64,
		SYNOPSYS_UNCONNECTED_65,
		SYNOPSYS_UNCONNECTED_66,
		SYNOPSYS_UNCONNECTED_67,
		SYNOPSYS_UNCONNECTED_68,
		SYNOPSYS_UNCONNECTED_69,
		SYNOPSYS_UNCONNECTED_70,
		SYNOPSYS_UNCONNECTED_71,
		SYNOPSYS_UNCONNECTED_72,
		SYNOPSYS_UNCONNECTED_73,
		SYNOPSYS_UNCONNECTED_74,
		SYNOPSYS_UNCONNECTED_75,
		SYNOPSYS_UNCONNECTED_76,
		SYNOPSYS_UNCONNECTED_77,
		SYNOPSYS_UNCONNECTED_78,
		SYNOPSYS_UNCONNECTED_79,
		SYNOPSYS_UNCONNECTED_80,
		SYNOPSYS_UNCONNECTED_81,
		SYNOPSYS_UNCONNECTED_82,
		SYNOPSYS_UNCONNECTED_83,
		SYNOPSYS_UNCONNECTED_84,
		SYNOPSYS_UNCONNECTED_85,
		SYNOPSYS_UNCONNECTED_86,
		SYNOPSYS_UNCONNECTED_87,
		SYNOPSYS_UNCONNECTED_88,
		SYNOPSYS_UNCONNECTED_89,
		SYNOPSYS_UNCONNECTED_90,
		SYNOPSYS_UNCONNECTED_91,
		SYNOPSYS_UNCONNECTED_92,
		SYNOPSYS_UNCONNECTED_93,
		SYNOPSYS_UNCONNECTED_94 }), 
	.remap(1'b0), 
	.sm_clken(1'b0), 
	.sm_ready(1'b0), 
	.sm_data_width_set0({ 1'b0,
		1'b0,
		1'b0 }), 
	.m_wr_data({ SYNOPSYS_UNCONNECTED_95,
		SYNOPSYS_UNCONNECTED_96,
		SYNOPSYS_UNCONNECTED_97,
		SYNOPSYS_UNCONNECTED_98,
		SYNOPSYS_UNCONNECTED_99,
		SYNOPSYS_UNCONNECTED_100,
		SYNOPSYS_UNCONNECTED_101,
		SYNOPSYS_UNCONNECTED_102,
		SYNOPSYS_UNCONNECTED_103,
		SYNOPSYS_UNCONNECTED_104,
		SYNOPSYS_UNCONNECTED_105,
		SYNOPSYS_UNCONNECTED_106,
		SYNOPSYS_UNCONNECTED_107,
		SYNOPSYS_UNCONNECTED_108,
		SYNOPSYS_UNCONNECTED_109,
		SYNOPSYS_UNCONNECTED_110 }), 
	.m_dout_valid({ SYNOPSYS_UNCONNECTED_111,
		SYNOPSYS_UNCONNECTED_112 }), 
	.s_ebi_gnt(1'b0), 
	.sm_ebi_gnt(1'b0), 
	.power_down(power_down), 
	.sf_power_down(1'b0), 
	.sm_power_down(1'b0), 
	.clear_sr_dp(clear_sr_dp), 
	.sf_clear_dp(1'b0), 
	.big_endian(FE_PHN5173_big_endian), 
	.miu_rd_data_out({ miu_data[31],
		miu_data[30],
		miu_data[29],
		miu_data[28],
		miu_data[27],
		miu_data[26],
		miu_data[25],
		miu_data[24],
		miu_data[23],
		miu_data[22],
		miu_data[21],
		miu_data[20],
		miu_data[19],
		miu_data[18],
		miu_data[17],
		miu_data[16],
		miu_data[15],
		miu_data[14],
		n2,
		miu_data[12],
		miu_data[11],
		miu_data[10],
		miu_data[9],
		miu_data[8],
		miu_data[7],
		miu_data[6],
		miu_data[5],
		miu_data[4],
		miu_data[3],
		miu_data[2],
		miu_data[1],
		miu_data[0] }), 
	.gpi(gpi), 
	.gpo(gpo), 
	.debug_ad_bank_addr(debug_ad_bank_addr), 
	.debug_ad_row_addr(debug_ad_row_addr), 
	.debug_ad_sf_bank_addr({ SYNOPSYS_UNCONNECTED_113,
		SYNOPSYS_UNCONNECTED_114 }), 
	.debug_ad_sf_row_addr({ SYNOPSYS_UNCONNECTED_115,
		SYNOPSYS_UNCONNECTED_116,
		SYNOPSYS_UNCONNECTED_117,
		SYNOPSYS_UNCONNECTED_118,
		SYNOPSYS_UNCONNECTED_119,
		SYNOPSYS_UNCONNECTED_120,
		SYNOPSYS_UNCONNECTED_121,
		SYNOPSYS_UNCONNECTED_122,
		SYNOPSYS_UNCONNECTED_123,
		SYNOPSYS_UNCONNECTED_124,
		SYNOPSYS_UNCONNECTED_125,
		SYNOPSYS_UNCONNECTED_126,
		SYNOPSYS_UNCONNECTED_127,
		SYNOPSYS_UNCONNECTED_128,
		SYNOPSYS_UNCONNECTED_129,
		SYNOPSYS_UNCONNECTED_130 }), 
	.debug_ad_sf_col_addr({ SYNOPSYS_UNCONNECTED_131,
		SYNOPSYS_UNCONNECTED_132,
		SYNOPSYS_UNCONNECTED_133,
		SYNOPSYS_UNCONNECTED_134,
		SYNOPSYS_UNCONNECTED_135,
		SYNOPSYS_UNCONNECTED_136,
		SYNOPSYS_UNCONNECTED_137,
		SYNOPSYS_UNCONNECTED_138,
		SYNOPSYS_UNCONNECTED_139,
		SYNOPSYS_UNCONNECTED_140,
		SYNOPSYS_UNCONNECTED_141,
		SYNOPSYS_UNCONNECTED_142,
		SYNOPSYS_UNCONNECTED_143,
		SYNOPSYS_UNCONNECTED_144,
		SYNOPSYS_UNCONNECTED_145,
		SYNOPSYS_UNCONNECTED_146 }), 
	.debug_smc_cs({ SYNOPSYS_UNCONNECTED_147,
		SYNOPSYS_UNCONNECTED_148,
		SYNOPSYS_UNCONNECTED_149,
		SYNOPSYS_UNCONNECTED_150 }), 
	.debug_ref_req(debug_ref_req), 
	.debug_ad_col_addr_15_(debug_ad_col_addr[15]), 
	.debug_ad_col_addr_14_(debug_ad_col_addr[14]), 
	.debug_ad_col_addr_11_(debug_ad_col_addr[11]), 
	.debug_ad_col_addr_10_(debug_ad_col_addr[10]), 
	.debug_ad_col_addr_9_(debug_ad_col_addr[9]), 
	.debug_ad_col_addr_8_(debug_ad_col_addr[8]), 
	.debug_ad_col_addr_7_(debug_ad_col_addr[7]), 
	.debug_ad_col_addr_6_(debug_ad_col_addr[6]), 
	.debug_ad_col_addr_5_(debug_ad_col_addr[5]), 
	.debug_ad_col_addr_4_(debug_ad_col_addr[4]), 
	.debug_ad_col_addr_3_(debug_ad_col_addr[3]), 
	.debug_ad_col_addr_2_(debug_ad_col_addr[2]), 
	.debug_ad_col_addr_1_(debug_ad_col_addr[1]), 
	.debug_ad_col_addr_0_(debug_ad_col_addr[0]), 
	.debug_ad_col_addr_13__BAR_BAR(debug_ad_col_addr[13]), 
	.debug_ad_col_addr_12__BAR_BAR(debug_ad_col_addr[12]), 
	.FE_OFN28_HRESETn(FE_OFN28_HRESETn), 
	.FE_OFN31_HRESETn(FE_OFN31_HRESETn), 
	.FE_OFN35_HRESETn(FE_OFN35_HRESETn), 
	.FE_OFN46_HRESETn(FE_OFN46_HRESETn), 
	.FE_OFN51_HRESETn(FE_OFN51_HRESETn), 
	.FE_OFN53_HRESETn(FE_OFN53_HRESETn), 
	.FE_OFN57_HRESETn(FE_OFN57_HRESETn), 
	.HCLK__L5_N11(HCLK__L5_N11), 
	.HCLK__L5_N12(HCLK__L5_N12), 
	.HCLK__L5_N17(HCLK__L5_N17), 
	.HCLK__L5_N28(HCLK__L5_N28), 
	.HCLK__L5_N29(HCLK__L5_N29), 
	.HCLK__L5_N30(HCLK__L5_N30), 
	.HCLK__L5_N31(HCLK__L5_N31), 
	.HCLK__L5_N32(HCLK__L5_N32), 
	.HCLK__L5_N33(HCLK__L5_N33), 
	.HCLK__L5_N34(HCLK__L5_N34), 
	.HCLK__L5_N35(HCLK__L5_N35), 
	.HCLK__L5_N36(HCLK__L5_N36), 
	.HCLK__L5_N6(HCLK__L5_N6), 
	.FE_OFN151_HRESETn(FE_OFN151_HRESETn), 
	.FE_OFN160_HRESETn(FE_OFN160_HRESETn), 
	.FE_OFN191_HRESETn(FE_OFN191_HRESETn), 
	.FE_OFN214_hiu_burst_size_4_(hiu_burst_size[4]), 
	.FE_OFN217_hiu_burst_size_2_(hiu_burst_size[2]), 
	.FE_OFN220_hiu_burst_size_0_(hiu_burst_size[0]));
endmodule

module cortexm0ds_logic (
	hclk, 
	hreset_n, 
	haddr_o, 
	hburst_o, 
	hmastlock_o, 
	hprot_o, 
	hsize_o, 
	htrans_o, 
	hwdata_o, 
	hwrite_o, 
	hrdata_i, 
	hready_i, 
	hresp_i, 
	nmi_i, 
	irq_i, 
	txev_o, 
	rxev_i, 
	lockup_o, 
	sys_reset_req_o, 
	sleeping_o, 
	vis_r0_o, 
	vis_r1_o, 
	vis_r2_o, 
	vis_r3_o, 
	vis_r4_o, 
	vis_r5_o, 
	vis_r6_o, 
	vis_r7_o, 
	vis_r8_o, 
	vis_r9_o, 
	vis_r10_o, 
	vis_r11_o, 
	vis_r12_o, 
	vis_r14_o, 
	vis_msp_o, 
	vis_psp_o, 
	vis_pc_o, 
	vis_apsr_o, 
	vis_tbit_o, 
	vis_ipsr_o, 
	vis_control_o, 
	vis_primask_o, 
	FE_OFN28_HRESETn, 
	FE_OFN29_HRESETn, 
	FE_OFN30_HRESETn, 
	FE_OFN34_HRESETn, 
	FE_OFN42_HRESETn, 
	FE_OFN43_HRESETn, 
	FE_OFN55_HRESETn, 
	SPCPT1_HADDR_29_, 
	HCLK__L5_N1, 
	HCLK__L5_N13, 
	HCLK__L5_N19, 
	HCLK__L5_N2, 
	HCLK__L5_N20, 
	HCLK__L5_N21, 
	HCLK__L5_N22, 
	HCLK__L5_N23, 
	HCLK__L5_N24, 
	HCLK__L5_N25, 
	HCLK__L5_N26, 
	HCLK__L5_N27, 
	HCLK__L5_N3, 
	HCLK__L5_N39, 
	HCLK__L5_N4, 
	HCLK__L5_N5, 
	HCLK__L5_N7, 
	HCLK__L5_N8, 
	HCLK__L5_N9);
   input hclk;
   input hreset_n;
   output [31:0] haddr_o;
   output [2:0] hburst_o;
   output hmastlock_o;
   output [3:0] hprot_o;
   output [2:0] hsize_o;
   output [1:0] htrans_o;
   output [31:0] hwdata_o;
   output hwrite_o;
   input [31:0] hrdata_i;
   input hready_i;
   input hresp_i;
   input nmi_i;
   input [15:0] irq_i;
   output txev_o;
   input rxev_i;
   output lockup_o;
   output sys_reset_req_o;
   output sleeping_o;
   output [31:0] vis_r0_o;
   output [31:0] vis_r1_o;
   output [31:0] vis_r2_o;
   output [31:0] vis_r3_o;
   output [31:0] vis_r4_o;
   output [31:0] vis_r5_o;
   output [31:0] vis_r6_o;
   output [31:0] vis_r7_o;
   output [31:0] vis_r8_o;
   output [31:0] vis_r9_o;
   output [31:0] vis_r10_o;
   output [31:0] vis_r11_o;
   output [31:0] vis_r12_o;
   output [31:0] vis_r14_o;
   output [29:0] vis_msp_o;
   output [29:0] vis_psp_o;
   output [30:0] vis_pc_o;
   output [3:0] vis_apsr_o;
   output vis_tbit_o;
   output [5:0] vis_ipsr_o;
   output vis_control_o;
   output vis_primask_o;
   input FE_OFN28_HRESETn;
   input FE_OFN29_HRESETn;
   input FE_OFN30_HRESETn;
   input FE_OFN34_HRESETn;
   input FE_OFN42_HRESETn;
   input FE_OFN43_HRESETn;
   input FE_OFN55_HRESETn;
   input SPCPT1_HADDR_29_;
   input HCLK__L5_N1;
   input HCLK__L5_N13;
   input HCLK__L5_N19;
   input HCLK__L5_N2;
   input HCLK__L5_N20;
   input HCLK__L5_N21;
   input HCLK__L5_N22;
   input HCLK__L5_N23;
   input HCLK__L5_N24;
   input HCLK__L5_N25;
   input HCLK__L5_N26;
   input HCLK__L5_N27;
   input HCLK__L5_N3;
   input HCLK__L5_N39;
   input HCLK__L5_N4;
   input HCLK__L5_N5;
   input HCLK__L5_N7;
   input HCLK__L5_N8;
   input HCLK__L5_N9;

   // Internal wires
   wire FE_PSN5239_n2057;
   wire FE_PSN5238_n3097;
   wire FE_PSN5237_n2184;
   wire FE_PSN5236_n16960;
   wire FE_PHN5254_n1134;
   wire FE_PHN5252_n389;
   wire FE_PHN5251_n5743;
   wire FE_PHN5250_n5747;
   wire FE_PHN5249_n5740;
   wire FE_PHN5248_n395;
   wire FE_PHN5247_n14432;
   wire FE_PHN5246_n1137;
   wire FE_PHN5245_n1134;
   wire FE_PHN5244_n4915;
   wire FE_PHN5243_n5745;
   wire FE_PHN5242_n5749;
   wire FE_PHN5238_n5748;
   wire FE_PHN5236_n5742;
   wire FE_PHN5233_n5760;
   wire FE_PHN5232_n385;
   wire FE_PHN5231_n1136;
   wire FE_PHN5230_n419;
   wire FE_PHN5229_n1135;
   wire FE_PHN5228_n1141;
   wire FE_PHN5227_n1138;
   wire FE_PHN5226_U227_Z_0;
   wire FE_PHN5225_n5746;
   wire FE_PHN5224_n5751;
   wire FE_PHN5223_n5752;
   wire FE_PHN5222_n5750;
   wire FE_PHN5221_n5763;
   wire FE_PHN5220_n5754;
   wire FE_PHN5219_n5756;
   wire FE_PHN5217_n380;
   wire FE_PHN5216_n1146;
   wire FE_PHN5215_n387;
   wire FE_PHN5214_n1133;
   wire FE_PHN5213_n1132;
   wire FE_PHN5212_n1130;
   wire FE_PHN5211_n1139;
   wire FE_PHN5210_n395;
   wire FE_PHN5209_n14432;
   wire FE_PHN5208_n389;
   wire FE_PHN5207_n1134;
   wire FE_PHN5206_n1137;
   wire FE_PHN5205_n5761;
   wire FE_PHN5204_n4915;
   wire FE_PHN5202_n5741;
   wire FE_PHN5201_n5744;
   wire FE_PHN5200_n5753;
   wire FE_PHN5199_n5766;
   wire FE_PHN5198_n5739;
   wire FE_PHN5197_n5765;
   wire FE_PHN5196_n5745;
   wire FE_PHN5195_n5749;
   wire FE_PHN5194_n5742;
   wire FE_PHN5193_n4389;
   wire FE_PHN5192_n17126;
   wire FE_PHN5188_n5768;
   wire FE_PHN5187_n5767;
   wire FE_PHN5186_n5769;
   wire FE_PHN5185_n5743;
   wire FE_PHN5184_n5748;
   wire FE_PHN5183_n5747;
   wire FE_PHN5182_n5740;
   wire FE_PHN5178_IRQ_15_;
   wire FE_PHN5177_IRQ_11_;
   wire FE_PHN5170_U591_Z_0;
   wire FE_PHN5169_n5349;
   wire FE_PHN5168_n5352;
   wire FE_PHN5167_n5081;
   wire FE_PHN5166_U503_Z_0;
   wire FE_PHN5163_n5262;
   wire FE_PHN5161_n4874;
   wire FE_PHN5160_n5362;
   wire FE_PHN5158_n4979;
   wire FE_PHN5156_n5361;
   wire FE_PHN5155_n5483;
   wire FE_PHN5151_n5128;
   wire FE_PHN5150_n5378;
   wire FE_PHN5149_n5347;
   wire FE_PHN5146_n5159;
   wire FE_PHN5145_U769_Z_0;
   wire FE_PHN5141_n4875;
   wire FE_PHN5139_n5319;
   wire FE_PHN5137_n5610;
   wire FE_PHN5136_n5360;
   wire FE_PHN5135_n5391;
   wire FE_PHN5134_n5413;
   wire FE_PHN5131_U247_Z_0;
   wire FE_PHN5130_n5369;
   wire FE_PHN5129_n5491;
   wire FE_PHN5127_n5018;
   wire FE_PHN5126_n5280;
   wire FE_PHN5125_n5443;
   wire FE_PHN5124_n5308;
   wire FE_PHN5123_n4848;
   wire FE_PHN5122_n5052;
   wire FE_PHN5121_n5089;
   wire FE_PHN5120_n5617;
   wire FE_PHN5119_U528_Z_0;
   wire FE_PHN5114_n5279;
   wire FE_PHN5113_U761_Z_0;
   wire FE_PHN5108_n5133;
   wire FE_PHN5107_n5538;
   wire FE_PHN5106_n5364;
   wire FE_PHN5105_n5204;
   wire FE_PHN5104_U583_Z_0;
   wire FE_PHN5099_n5611;
   wire FE_PHN5097_U646_Z_0;
   wire FE_PHN5096_U428_Z_0;
   wire FE_PHN5094_n5142;
   wire FE_PHN5093_n5220;
   wire FE_PHN5091_U359_Z_0;
   wire FE_PHN5090_n5201;
   wire FE_PHN5089_U644_Z_0;
   wire FE_PHN5088_n5355;
   wire FE_PHN5086_n5202;
   wire FE_PHN5085_n5337;
   wire FE_PHN5084_U275_Z_0;
   wire FE_PHN5080_U711_Z_0;
   wire FE_PHN5077_U589_Z_0;
   wire FE_PHN5076_U595_Z_0;
   wire FE_PHN5074_n5260;
   wire FE_PHN5066_n5653;
   wire FE_PHN5065_n5223;
   wire FE_PHN5061_n5042;
   wire FE_PHN5060_n5136;
   wire FE_PHN5059_n5367;
   wire FE_PHN5055_n5209;
   wire FE_PHN5053_n5271;
   wire FE_PHN5052_n5383;
   wire FE_PHN5050_n5511;
   wire FE_PHN5049_U677_Z_0;
   wire FE_PHN5046_n4963;
   wire FE_PHN5045_n5200;
   wire FE_PHN5044_n5339;
   wire FE_PHN5043_n4878;
   wire FE_PHN5039_U441_Z_0;
   wire FE_PHN5035_n5602;
   wire FE_PHN5034_n5104;
   wire FE_PHN5031_U784_Z_0;
   wire FE_PHN5029_n5084;
   wire FE_PHN5028_n4995;
   wire FE_PHN5027_n5384;
   wire FE_PHN5026_U363_Z_0;
   wire FE_PHN5025_U309_Z_0;
   wire FE_PHN5023_n5381;
   wire FE_PHN5019_n5492;
   wire FE_PHN5018_n5493;
   wire FE_PHN5017_n5221;
   wire FE_PHN5015_n5489;
   wire FE_PHN5014_n5294;
   wire FE_PHN5013_n5307;
   wire FE_PHN5010_n4924;
   wire FE_PHN5008_n5019;
   wire FE_PHN5006_n5640;
   wire FE_PHN5002_n5643;
   wire FE_PHN5001_n5376;
   wire FE_PHN5000_n5508;
   wire FE_PHN4999_U320_Z_0;
   wire FE_PHN4997_n5490;
   wire FE_PHN4995_n5109;
   wire FE_PHN4994_n5336;
   wire FE_PHN4991_U234_Z_0;
   wire FE_PHN4990_n5092;
   wire FE_PHN4989_n5496;
   wire FE_PHN4988_n5218;
   wire FE_PHN4986_U800_Z_0;
   wire FE_PHN4985_n5792;
   wire FE_PHN4984_U305_Z_0;
   wire FE_PHN4983_U557_Z_0;
   wire FE_PHN4982_U606_Z_0;
   wire FE_PHN4980_n5283;
   wire FE_PHN4977_n5353;
   wire FE_PHN4976_n5599;
   wire FE_PHN4974_n5634;
   wire FE_PHN4972_n5261;
   wire FE_PHN4971_n5380;
   wire FE_PHN4970_n5365;
   wire FE_PHN4969_n5198;
   wire FE_PHN4967_n5394;
   wire FE_PHN4963_n5356;
   wire FE_PHN4960_U324_Z_0;
   wire FE_PHN4959_n5350;
   wire FE_PHN4958_U411_Z_0;
   wire FE_PHN4956_n5073;
   wire FE_PHN4955_n5214;
   wire FE_PHN4954_U471_Z_0;
   wire FE_PHN4953_n5066;
   wire FE_PHN4950_n5403;
   wire FE_PHN4949_n5515;
   wire FE_PHN4947_n5357;
   wire FE_PHN4946_n5372;
   wire FE_PHN4944_U323_Z_0;
   wire FE_PHN4943_U566_Z_0;
   wire FE_PHN4941_n5275;
   wire FE_PHN4940_n5379;
   wire FE_PHN4937_n5788;
   wire FE_PHN4935_n5390;
   wire FE_PHN4933_n5226;
   wire FE_PHN4932_U506_Z_0;
   wire FE_PHN4931_n5273;
   wire FE_PHN4930_U563_Z_0;
   wire FE_PHN4927_U395_Z_0;
   wire FE_PHN4924_n5286;
   wire FE_PHN4923_U318_Z_0;
   wire FE_PHN4921_U673_Z_0;
   wire FE_PHN4920_U726_Z_0;
   wire FE_PHN4919_n5494;
   wire FE_PHN4916_n5738;
   wire FE_PHN4912_n5335;
   wire FE_PHN4911_n5210;
   wire FE_PHN4910_n5497;
   wire FE_PHN4909_n5277;
   wire FE_PHN4907_U619_Z_0;
   wire FE_PHN4906_n5541;
   wire FE_PHN4905_U692_Z_0;
   wire FE_PHN4904_n5374;
   wire FE_PHN4902_n5479;
   wire FE_PHN4900_U263_Z_0;
   wire FE_PHN4898_n5495;
   wire FE_PHN4897_U513_Z_0;
   wire FE_PHN4896_n5134;
   wire FE_PHN4895_U745_Z_0;
   wire FE_PHN4891_U663_Z_0;
   wire FE_PHN4890_U481_Z_0;
   wire FE_PHN4888_n4998;
   wire FE_PHN4887_n5341;
   wire FE_PHN4886_n5216;
   wire FE_PHN4885_n5559;
   wire FE_PHN4884_U504_Z_0;
   wire FE_PHN4883_n5354;
   wire FE_PHN4882_U660_Z_0;
   wire FE_PHN4876_n5480;
   wire FE_PHN4874_n5630;
   wire FE_PHN4873_n5566;
   wire FE_PHN4870_n5334;
   wire FE_PHN4869_U475_Z_0;
   wire FE_PHN4868_n5608;
   wire FE_PHN4867_n5506;
   wire FE_PHN4866_n5037;
   wire FE_PHN4865_U500_Z_0;
   wire FE_PHN4864_U585_Z_0;
   wire FE_PHN4863_U466_Z_0;
   wire FE_PHN4862_U291_Z_0;
   wire FE_PHN4861_n5278;
   wire FE_PHN4860_U779_Z_0;
   wire FE_PHN4859_n5563;
   wire FE_PHN4857_U667_Z_0;
   wire FE_PHN4854_n5276;
   wire FE_PHN4853_n5063;
   wire FE_PHN4850_n5168;
   wire FE_PHN4847_n5382;
   wire FE_PHN4844_U712_Z_0;
   wire FE_PHN4840_n5577;
   wire FE_PHN4839_n5569;
   wire FE_PHN4838_n5131;
   wire FE_PHN4835_U454_Z_0;
   wire FE_PHN4834_U743_Z_0;
   wire FE_PHN4833_n5343;
   wire FE_PHN4831_n4982;
   wire FE_PHN4830_U748_Z_0;
   wire FE_PHN4829_n5791;
   wire FE_PHN4828_n5574;
   wire FE_PHN4827_n5087;
   wire FE_PHN4823_n5631;
   wire FE_PHN4822_n5389;
   wire FE_PHN4821_n5607;
   wire FE_PHN4820_U242_Z_0;
   wire FE_PHN4815_U651_Z_0;
   wire FE_PHN4814_U445_Z_0;
   wire FE_PHN4813_n5683;
   wire FE_PHN4810_U708_Z_0;
   wire FE_PHN4809_n5264;
   wire FE_PHN4808_n5345;
   wire FE_PHN4807_n5340;
   wire FE_PHN4804_n14928;
   wire FE_PHN4802_n5263;
   wire FE_PHN4801_n5543;
   wire FE_PHN4797_U325_Z_0;
   wire FE_PHN4796_n5122;
   wire FE_PHN4795_n5368;
   wire FE_PHN4794_n5215;
   wire FE_PHN4790_n5125;
   wire FE_PHN4788_U496_Z_0;
   wire FE_PHN4784_n5627;
   wire FE_PHN4783_n4938;
   wire FE_PHN4782_n5548;
   wire FE_PHN4781_U728_Z_0;
   wire FE_PHN4779_n4937;
   wire FE_PHN4778_n5614;
   wire FE_PHN4774_U683_Z_0;
   wire FE_PHN4772_U628_Z_0;
   wire FE_PHN4767_n5265;
   wire FE_PHN4761_U634_Z_0;
   wire FE_PHN4756_n5056;
   wire FE_PHN4750_n5565;
   wire FE_PHN4749_n4925;
   wire FE_PHN4748_n276;
   wire FE_PHN4743_U656_Z_0;
   wire FE_PHN4739_n5586;
   wire FE_PHN4737_n5712;
   wire FE_PHN4735_n4939;
   wire FE_PHN4734_n5555;
   wire FE_PHN4733_n4935;
   wire FE_PHN4732_n5561;
   wire FE_PHN4731_n4936;
   wire FE_PHN4730_n4926;
   wire FE_PHN4729_n4942;
   wire FE_PHN4726_n5760;
   wire FE_PHN4725_n385;
   wire FE_PHN4724_n1136;
   wire FE_PHN4723_n419;
   wire FE_PHN4722_n1135;
   wire FE_PHN4721_n1141;
   wire FE_PHN4720_n1138;
   wire FE_PHN4712_n4923;
   wire FE_PHN4711_U227_Z_0;
   wire FE_PHN4710_n5751;
   wire FE_PHN4709_n5752;
   wire FE_PHN4708_n5746;
   wire FE_PHN4707_n5750;
   wire FE_PHN4706_n5763;
   wire FE_PHN4704_n5754;
   wire FE_PHN4703_n5756;
   wire FE_PHN4702_n1146;
   wire FE_PHN4701_n380;
   wire FE_PHN4700_n387;
   wire FE_PHN4699_n1132;
   wire FE_PHN4698_n1133;
   wire FE_PHN4697_n1130;
   wire FE_PHN4696_n1139;
   wire FE_PHN4695_n395;
   wire FE_PHN4694_n14432;
   wire FE_PHN4693_n389;
   wire FE_PHN4692_n4917;
   wire FE_PHN4691_n4919;
   wire FE_PHN4690_n4918;
   wire FE_PHN4689_n5761;
   wire FE_PHN4688_n4915;
   wire FE_PHN4687_n5741;
   wire FE_PHN4686_n5744;
   wire FE_PHN4685_n5753;
   wire FE_PHN4684_n5766;
   wire FE_PHN4683_n5739;
   wire FE_PHN4682_n5765;
   wire FE_PHN4681_n5745;
   wire FE_PHN4680_n5749;
   wire FE_PHN4679_n5742;
   wire FE_PHN4675_n4902;
   wire FE_PHN4674_n4394;
   wire FE_PHN4673_n4389;
   wire FE_PHN4672_n4300;
   wire FE_PHN4671_n4903;
   wire FE_PHN4670_n4193;
   wire FE_PHN4669_n4324;
   wire FE_PHN4668_n4391;
   wire FE_PHN4667_n4397;
   wire FE_PHN4666_n4190;
   wire FE_PHN4662_n5768;
   wire FE_PHN4661_n5767;
   wire FE_PHN4660_n5769;
   wire FE_PHN4659_n5743;
   wire FE_PHN4658_n5747;
   wire FE_PHN4657_n5748;
   wire FE_PHN4656_n5740;
   wire FE_PHN4655_n4909;
   wire FE_PHN4654_n4912;
   wire FE_PHN4653_n3273;
   wire FE_PHN4652_n4920;
   wire FE_PHN4641_IRQ_14_;
   wire FE_PHN4639_n5692;
   wire FE_PHN4638_IRQ_11_;
   wire FE_PHN4637_IRQ_9_;
   wire FE_PHN4634_IRQ_1_;
   wire FE_PHN4631_NMI;
   wire FE_PHN4630_IRQ_15_;
   wire FE_PHN4629_n17127;
   wire FE_PHN4624_n17126;
   wire FE_PHN4615_U762_Z_0;
   wire FE_PHN4611_n5710;
   wire FE_PHN4608_U802_Z_0;
   wire FE_PHN4607_n5652;
   wire FE_PHN4602_n4890;
   wire FE_PHN4601_U317_Z_0;
   wire FE_PHN4597_U789_Z_0;
   wire FE_PHN4596_U781_Z_0;
   wire FE_PHN4595_U791_Z_0;
   wire FE_PHN4590_U518_Z_0;
   wire FE_PHN4588_n5704;
   wire FE_PHN4586_n5097;
   wire FE_PHN4585_n5706;
   wire FE_PHN4584_n5737;
   wire FE_PHN4583_n5651;
   wire FE_PHN4580_U763_Z_0;
   wire FE_PHN4579_n5705;
   wire FE_PHN4577_n5612;
   wire FE_PHN4576_U782_Z_0;
   wire FE_PHN4575_n4862;
   wire FE_PHN4573_n5130;
   wire FE_PHN4572_U783_Z_0;
   wire FE_PHN4571_U144_Z_0;
   wire FE_PHN4570_n5568;
   wire FE_PHN4569_n5103;
   wire FE_PHN4567_n5172;
   wire FE_PHN4566_U771_Z_0;
   wire FE_PHN4565_n5015;
   wire FE_PHN4564_n5012;
   wire FE_PHN4563_n5450;
   wire FE_PHN4562_n5702;
   wire FE_PHN4561_n4857;
   wire FE_PHN4560_n5267;
   wire FE_PHN4559_n5457;
   wire FE_PHN4557_n5299;
   wire FE_PHN4556_n5396;
   wire FE_PHN4555_U772_Z_0;
   wire FE_PHN4554_n5178;
   wire FE_PHN4553_n5604;
   wire FE_PHN4552_n4885;
   wire FE_PHN4550_n4856;
   wire FE_PHN4549_n5284;
   wire FE_PHN4548_n5449;
   wire FE_PHN4545_n5420;
   wire FE_PHN4544_n5770;
   wire FE_PHN4541_n5772;
   wire FE_PHN4540_n5297;
   wire FE_PHN4539_n5428;
   wire FE_PHN4538_n5187;
   wire FE_PHN4536_n5603;
   wire FE_PHN4535_n5641;
   wire FE_PHN4534_n5072;
   wire FE_PHN4533_n5062;
   wire FE_PHN4532_n5135;
   wire FE_PHN4531_n5174;
   wire FE_PHN4529_n5300;
   wire FE_PHN4526_U788_Z_0;
   wire FE_PHN4525_n5433;
   wire FE_PHN4524_U691_Z_0;
   wire FE_PHN4523_n5487;
   wire FE_PHN4518_n5141;
   wire FE_PHN4517_n5115;
   wire FE_PHN4516_n5288;
   wire FE_PHN4515_n5083;
   wire FE_PHN4514_n5468;
   wire FE_PHN4512_U770_Z_0;
   wire FE_PHN4511_n5170;
   wire FE_PHN4510_n5040;
   wire FE_PHN4509_n5622;
   wire FE_PHN4508_n5463;
   wire FE_PHN4506_n5470;
   wire FE_PHN4505_n5169;
   wire FE_PHN4504_n5181;
   wire FE_PHN4500_n5039;
   wire FE_PHN4499_n5138;
   wire FE_PHN4496_n5461;
   wire FE_PHN4495_n5075;
   wire FE_PHN4494_n5472;
   wire FE_PHN4493_n5557;
   wire FE_PHN4492_n5186;
   wire FE_PHN4490_n5453;
   wire FE_PHN4488_n4884;
   wire FE_PHN4487_n5478;
   wire FE_PHN4486_n4969;
   wire FE_PHN4485_n5196;
   wire FE_PHN4484_n4985;
   wire FE_PHN4482_n5455;
   wire FE_PHN4481_n5459;
   wire FE_PHN4479_U787_Z_0;
   wire FE_PHN4478_U775_Z_0;
   wire FE_PHN4477_n5173;
   wire FE_PHN4476_n5633;
   wire FE_PHN4475_n5597;
   wire FE_PHN4474_n5427;
   wire FE_PHN4472_n4869;
   wire FE_PHN4471_n5190;
   wire FE_PHN4468_n5426;
   wire FE_PHN4467_n5553;
   wire FE_PHN4466_n5312;
   wire FE_PHN4463_n5161;
   wire FE_PHN4462_n5564;
   wire FE_PHN4460_n5469;
   wire FE_PHN4459_n5401;
   wire FE_PHN4458_n5437;
   wire FE_PHN4457_n5121;
   wire FE_PHN4456_n5197;
   wire FE_PHN4454_U786_Z_0;
   wire FE_PHN4453_U459_Z_0;
   wire FE_PHN4452_n5296;
   wire FE_PHN4451_n5598;
   wire FE_PHN4450_n5486;
   wire FE_PHN4449_n5021;
   wire FE_PHN4448_n5576;
   wire FE_PHN4447_n5567;
   wire FE_PHN4446_n5093;
   wire FE_PHN4444_n5447;
   wire FE_PHN4441_U764_Z_0;
   wire FE_PHN4440_n5616;
   wire FE_PHN4439_n5600;
   wire FE_PHN4438_n5636;
   wire FE_PHN4437_n5046;
   wire FE_PHN4436_n5464;
   wire FE_PHN4433_n5579;
   wire FE_PHN4432_n5086;
   wire FE_PHN4431_n4865;
   wire FE_PHN4430_n5485;
   wire FE_PHN4427_n5020;
   wire FE_PHN4426_n5366;
   wire FE_PHN4425_n5558;
   wire FE_PHN4422_n5392;
   wire FE_PHN4421_n5477;
   wire FE_PHN4420_n5539;
   wire FE_PHN4419_n5444;
   wire FE_PHN4418_n5022;
   wire FE_PHN4417_n5398;
   wire FE_PHN4416_n5067;
   wire FE_PHN4413_n5430;
   wire FE_PHN4412_n5442;
   wire FE_PHN4411_n5434;
   wire FE_PHN4407_n4870;
   wire FE_PHN4406_n5432;
   wire FE_PHN4405_n5476;
   wire FE_PHN4404_n5171;
   wire FE_PHN4403_n5438;
   wire FE_PHN4402_n5033;
   wire FE_PHN4401_n5287;
   wire FE_PHN4400_n5397;
   wire FE_PHN4399_n5606;
   wire FE_PHN4396_n5452;
   wire FE_PHN4394_U774_Z_0;
   wire FE_PHN4393_n5462;
   wire FE_PHN4392_n5575;
   wire FE_PHN4387_n5069;
   wire FE_PHN4386_n5439;
   wire FE_PHN4385_n5182;
   wire FE_PHN4383_n4891;
   wire FE_PHN4382_n5424;
   wire FE_PHN4380_n5550;
   wire FE_PHN4379_n5412;
   wire FE_PHN4378_n5448;
   wire FE_PHN4377_n5421;
   wire FE_PHN4376_n5184;
   wire FE_PHN4375_n5466;
   wire FE_PHN4374_n5298;
   wire FE_PHN4373_n5030;
   wire FE_PHN4372_n5010;
   wire FE_PHN4371_n5175;
   wire FE_PHN4369_n5041;
   wire FE_PHN4368_n5123;
   wire FE_PHN4367_n5411;
   wire FE_PHN4366_n5414;
   wire FE_PHN4364_n5074;
   wire FE_PHN4363_n5108;
   wire FE_PHN4362_n5043;
   wire FE_PHN4361_n4987;
   wire FE_PHN4358_n4872;
   wire FE_PHN4357_n5192;
   wire FE_PHN4356_n5191;
   wire FE_PHN4355_n5441;
   wire FE_PHN4352_n5473;
   wire FE_PHN4351_n5051;
   wire FE_PHN4350_n5091;
   wire FE_PHN4348_n5410;
   wire FE_PHN4346_n5316;
   wire FE_PHN4343_n5419;
   wire FE_PHN4340_n5106;
   wire FE_PHN4338_n5132;
   wire FE_PHN4337_n5509;
   wire FE_PHN4336_n5304;
   wire FE_PHN4335_n5386;
   wire FE_PHN4334_n5393;
   wire FE_PHN4333_n5395;
   wire FE_PHN4332_n5180;
   wire FE_PHN4331_n5399;
   wire FE_PHN4330_n5435;
   wire FE_PHN4329_n5205;
   wire FE_PHN4327_n5183;
   wire FE_PHN4326_U279_Z_0;
   wire FE_PHN4325_n4986;
   wire FE_PHN4324_U105_Z_0;
   wire FE_PHN4322_U780_Z_0;
   wire FE_PHN4320_n5451;
   wire FE_PHN4319_n5189;
   wire FE_PHN4318_n5521;
   wire FE_PHN4317_n5289;
   wire FE_PHN4316_n5799;
   wire FE_PHN4314_n5629;
   wire FE_PHN4313_n5596;
   wire FE_PHN4312_n5199;
   wire FE_PHN4311_n5195;
   wire FE_PHN4305_n5422;
   wire FE_PHN4303_U766_Z_0;
   wire FE_PHN4302_n5440;
   wire FE_PHN4301_n5409;
   wire FE_PHN4298_U785_Z_0;
   wire FE_PHN4297_U261_Z_0;
   wire FE_PHN4295_n5436;
   wire FE_PHN4291_n5207;
   wire FE_PHN4289_n4854;
   wire FE_PHN4288_n1319;
   wire FE_PHN4287_n5415;
   wire FE_PHN4283_n5309;
   wire FE_PHN4282_n5418;
   wire FE_PHN4280_n5624;
   wire FE_PHN4279_n5301;
   wire FE_PHN4274_n5176;
   wire FE_PHN4273_n5225;
   wire FE_PHN4272_U479_Z_0;
   wire FE_PHN4271_n5159;
   wire FE_PHN4270_U509_Z_0;
   wire FE_PHN4269_U429_Z_0;
   wire FE_PHN4267_n5363;
   wire FE_PHN4266_n5483;
   wire FE_PHN4264_U777_Z_0;
   wire FE_PHN4263_n5028;
   wire FE_PHN4262_n5013;
   wire FE_PHN4261_n5481;
   wire FE_PHN4260_n5045;
   wire FE_PHN4259_n5049;
   wire FE_PHN4258_n5081;
   wire FE_PHN4257_n5318;
   wire FE_PHN4249_n5308;
   wire FE_PHN4248_n5203;
   wire FE_PHN4247_n5270;
   wire FE_PHN4240_n5364;
   wire FE_PHN4237_n5076;
   wire FE_PHN4235_n5413;
   wire FE_PHN4234_n5224;
   wire FE_PHN4233_n5542;
   wire FE_PHN4232_U359_Z_0;
   wire FE_PHN4231_n5443;
   wire FE_PHN4230_n5268;
   wire FE_PHN4229_U761_Z_0;
   wire FE_PHN4227_n5317;
   wire FE_PHN4221_n5360;
   wire FE_PHN4220_n5361;
   wire FE_PHN4219_n4979;
   wire FE_PHN4218_n5202;
   wire FE_PHN4217_n5079;
   wire FE_PHN4216_n5514;
   wire FE_PHN4215_n5638;
   wire FE_PHN4214_n5621;
   wire FE_PHN4213_n5391;
   wire FE_PHN4212_U590_Z_0;
   wire FE_PHN4205_n5538;
   wire FE_PHN4202_U784_Z_0;
   wire FE_PHN4201_n5643;
   wire FE_PHN4200_n5112;
   wire FE_PHN4199_n5369;
   wire FE_PHN4198_n5209;
   wire FE_PHN4196_U275_Z_0;
   wire FE_PHN4193_n5266;
   wire FE_PHN4192_n5384;
   wire FE_PHN4191_n5018;
   wire FE_PHN4187_n4995;
   wire FE_PHN4185_n5511;
   wire FE_PHN4182_n5348;
   wire FE_PHN4181_n5554;
   wire FE_PHN4180_n5610;
   wire FE_PHN4178_n5070;
   wire FE_PHN4177_n5273;
   wire FE_PHN4176_n5394;
   wire FE_PHN4175_n5200;
   wire FE_PHN4174_U243_Z_0;
   wire FE_PHN4172_n5367;
   wire FE_PHN4171_n5019;
   wire FE_PHN4170_n5319;
   wire FE_PHN4169_n5261;
   wire FE_PHN4168_n5136;
   wire FE_PHN4167_n5139;
   wire FE_PHN4166_n5133;
   wire FE_PHN4165_n5280;
   wire FE_PHN4161_n5107;
   wire FE_PHN4160_n5218;
   wire FE_PHN4154_n5213;
   wire FE_PHN4150_n5362;
   wire FE_PHN4149_n5560;
   wire FE_PHN4148_n5383;
   wire FE_PHN4147_n5279;
   wire FE_PHN4146_n5357;
   wire FE_PHN4145_n5405;
   wire FE_PHN4142_n5365;
   wire FE_PHN4141_n5376;
   wire FE_PHN4140_n5217;
   wire FE_PHN4139_n5611;
   wire FE_PHN4138_U295_Z_0;
   wire FE_PHN4136_n5640;
   wire FE_PHN4135_n5339;
   wire FE_PHN4133_n4874;
   wire FE_PHN4132_n5517;
   wire FE_PHN4129_n5201;
   wire FE_PHN4126_n5776;
   wire FE_PHN4124_n5356;
   wire FE_PHN4123_n5124;
   wire FE_PHN4122_n5489;
   wire FE_PHN4120_n5403;
   wire FE_PHN4119_n5294;
   wire FE_PHN4118_n5277;
   wire FE_PHN4117_n5084;
   wire FE_PHN4115_n5335;
   wire FE_PHN4109_n5219;
   wire FE_PHN4108_n5599;
   wire FE_PHN4104_n4878;
   wire FE_PHN4102_n5109;
   wire FE_PHN4101_n5562;
   wire FE_PHN4096_U506_Z_0;
   wire FE_PHN4094_n5492;
   wire FE_PHN4093_n5493;
   wire FE_PHN4090_n5349;
   wire FE_PHN4089_n5352;
   wire FE_PHN4088_n5496;
   wire FE_PHN4085_n5374;
   wire FE_PHN4084_n5479;
   wire FE_PHN4083_n5347;
   wire FE_PHN4082_n5334;
   wire FE_PHN4078_n5508;
   wire FE_PHN4077_n5480;
   wire FE_PHN4076_n5044;
   wire FE_PHN4072_n5221;
   wire FE_PHN4067_n5292;
   wire FE_PHN4061_n5630;
   wire FE_PHN4060_n5278;
   wire FE_PHN4059_n5491;
   wire FE_PHN4058_n5089;
   wire FE_PHN4057_n5378;
   wire FE_PHN4054_U475_Z_0;
   wire FE_PHN4053_U660_Z_0;
   wire FE_PHN4052_n5355;
   wire FE_PHN4051_n5286;
   wire FE_PHN4050_n5635;
   wire FE_PHN4048_U726_Z_0;
   wire FE_PHN4047_U257_Z_0;
   wire FE_PHN4044_n5271;
   wire FE_PHN4043_n5336;
   wire FE_PHN4042_n5372;
   wire FE_PHN4041_n5214;
   wire FE_PHN4040_n5052;
   wire FE_PHN4039_U441_Z_0;
   wire FE_PHN4035_U779_Z_0;
   wire FE_PHN4034_U606_Z_0;
   wire FE_PHN4032_n5128;
   wire FE_PHN4031_n5220;
   wire FE_PHN4027_n5343;
   wire FE_PHN4026_n5337;
   wire FE_PHN4024_U411_Z_0;
   wire FE_PHN4023_U673_Z_0;
   wire FE_PHN4022_n5350;
   wire FE_PHN4021_n5617;
   wire FE_PHN4020_n5541;
   wire FE_PHN4018_n5566;
   wire FE_PHN4017_n5379;
   wire FE_PHN4012_n5602;
   wire FE_PHN4005_n4998;
   wire FE_PHN4004_n5211;
   wire FE_PHN4003_n5063;
   wire FE_PHN4002_n5104;
   wire FE_PHN4001_n5087;
   wire FE_PHN4000_n4984;
   wire FE_PHN3989_U448_Z_0;
   wire FE_PHN3987_n5216;
   wire FE_PHN3986_n5497;
   wire FE_PHN3985_n5577;
   wire FE_PHN3983_n5263;
   wire FE_PHN3982_n5260;
   wire FE_PHN3981_n5559;
   wire FE_PHN3977_n5495;
   wire FE_PHN3976_U395_Z_0;
   wire FE_PHN3975_n5385;
   wire FE_PHN3974_n5381;
   wire FE_PHN3973_n5042;
   wire FE_PHN3972_n5490;
   wire FE_PHN3971_U291_Z_0;
   wire FE_PHN3970_n5037;
   wire FE_PHN3969_n5092;
   wire FE_PHN3963_n5125;
   wire FE_PHN3962_n5634;
   wire FE_PHN3961_n5283;
   wire FE_PHN3960_n5631;
   wire FE_PHN3959_n5608;
   wire FE_PHN3958_n5353;
   wire FE_PHN3954_n5569;
   wire FE_PHN3950_U325_Z_0;
   wire FE_PHN3949_n5382;
   wire FE_PHN3948_n5198;
   wire FE_PHN3943_n5307;
   wire FE_PHN3942_n5563;
   wire FE_PHN3941_n5548;
   wire FE_PHN3937_n5131;
   wire FE_PHN3934_n4875;
   wire FE_PHN3931_n5368;
   wire FE_PHN3930_n5275;
   wire FE_PHN3928_n5515;
   wire FE_PHN3927_n5116;
   wire FE_PHN3926_n5574;
   wire FE_PHN3925_U329_Z_0;
   wire FE_PHN3924_n5607;
   wire FE_PHN3923_n5351;
   wire FE_PHN3922_n5627;
   wire FE_PHN3921_n5204;
   wire FE_PHN3919_n5122;
   wire FE_PHN3918_n5264;
   wire FE_PHN3917_n5226;
   wire FE_PHN3916_n5073;
   wire FE_PHN3915_n5380;
   wire FE_PHN3912_n5212;
   wire FE_PHN3911_n5276;
   wire FE_PHN3910_n5370;
   wire FE_PHN3909_n5215;
   wire FE_PHN3908_n5543;
   wire FE_PHN3907_n5494;
   wire FE_PHN3906_n5016;
   wire FE_PHN3904_U624_Z_0;
   wire FE_PHN3903_U644_Z_0;
   wire FE_PHN3902_n5650;
   wire FE_PHN3900_U386_Z_0;
   wire FE_PHN3898_n5389;
   wire FE_PHN3896_n5345;
   wire FE_PHN3893_n5341;
   wire FE_PHN3892_n5210;
   wire FE_PHN3888_n5614;
   wire FE_PHN3887_U712_Z_0;
   wire FE_PHN3886_n5262;
   wire FE_PHN3885_U239_Z_0;
   wire FE_PHN3884_n5354;
   wire FE_PHN3883_n4963;
   wire FE_PHN3882_U466_Z_0;
   wire FE_PHN3880_n5738;
   wire FE_PHN3879_n5340;
   wire FE_PHN3878_U353_Z_0;
   wire FE_PHN3877_U234_Z_0;
   wire FE_PHN3875_n5390;
   wire FE_PHN3874_n5142;
   wire FE_PHN3872_n5066;
   wire FE_PHN3871_n5506;
   wire FE_PHN3869_U769_Z_0;
   wire FE_PHN3868_U503_Z_0;
   wire FE_PHN3866_n5265;
   wire FE_PHN3865_U345_Z_0;
   wire FE_PHN3864_U428_Z_0;
   wire FE_PHN3863_U646_Z_0;
   wire FE_PHN3862_U711_Z_0;
   wire FE_PHN3857_U363_Z_0;
   wire FE_PHN3856_U677_Z_0;
   wire FE_PHN3853_U628_Z_0;
   wire FE_PHN3851_U504_Z_0;
   wire FE_PHN3847_U471_Z_0;
   wire FE_PHN3845_U800_Z_0;
   wire FE_PHN3843_U619_Z_0;
   wire FE_PHN3842_U263_Z_0;
   wire FE_PHN3839_U745_Z_0;
   wire FE_PHN3836_U612_Z_0;
   wire FE_PHN3828_n5168;
   wire FE_PHN3823_U585_Z_0;
   wire FE_PHN3821_U481_Z_0;
   wire FE_PHN3814_U425_Z_0;
   wire FE_PHN3811_U513_Z_0;
   wire FE_PHN3808_n270;
   wire FE_PHN3806_U663_Z_0;
   wire FE_PHN3803_U748_Z_0;
   wire FE_PHN3802_U490_Z_0;
   wire FE_PHN3799_U335_Z_0;
   wire FE_PHN3798_U454_Z_0;
   wire FE_PHN3797_U391_Z_0;
   wire FE_PHN3796_U754_Z_0;
   wire FE_PHN3793_n4982;
   wire FE_PHN3787_U242_Z_0;
   wire FE_PHN3785_U667_Z_0;
   wire FE_PHN3784_U651_Z_0;
   wire FE_PHN3782_U728_Z_0;
   wire FE_PHN3780_n5134;
   wire FE_PHN3779_n286;
   wire FE_PHN3778_U743_Z_0;
   wire FE_PHN3775_U500_Z_0;
   wire FE_PHN3774_U708_Z_0;
   wire FE_PHN3769_U407_Z_0;
   wire FE_PHN3765_U683_Z_0;
   wire FE_PHN3764_n5004;
   wire FE_PHN3763_U233_Z_0;
   wire FE_PHN3762_U496_Z_0;
   wire FE_PHN3755_n8706;
   wire FE_PHN3753_U445_Z_0;
   wire FE_PHN3744_U610_Z_0;
   wire FE_PHN3735_n284;
   wire FE_PHN3733_U463_Z_0;
   wire FE_PHN3730_U497_Z_0;
   wire FE_PHN3726_n5193;
   wire FE_PHN3725_U594_Z_0;
   wire FE_PHN3718_U680_Z_0;
   wire FE_PHN3717_n278;
   wire FE_PHN3699_n5056;
   wire FE_PHN3690_n8698;
   wire FE_PHN3682_U634_Z_0;
   wire FE_PHN3681_n5302;
   wire FE_PHN3663_U656_Z_0;
   wire FE_PHN3662_n276;
   wire FE_PHN3661_n4852;
   wire FE_PHN3654_n5733;
   wire FE_PHN3648_n5594;
   wire FE_PHN3647_U493_Z_0;
   wire FE_PHN3642_n5179;
   wire FE_PHN3641_n282;
   wire FE_PHN3639_n5735;
   wire FE_PHN3637_n5429;
   wire FE_PHN3636_U341_Z_0;
   wire FE_PHN3635_n5645;
   wire FE_PHN3634_n5475;
   wire FE_PHN3633_n4989;
   wire FE_PHN3631_n294;
   wire FE_PHN3630_n5194;
   wire FE_PHN3629_n5400;
   wire FE_PHN3627_n5147;
   wire FE_PHN3626_n5446;
   wire FE_PHN3625_n5732;
   wire FE_PHN3624_n4992;
   wire FE_PHN3623_n5058;
   wire FE_PHN3622_n5416;
   wire FE_PHN3621_n5499;
   wire FE_PHN3620_n4848;
   wire FE_PHN3617_n5586;
   wire FE_PHN3616_n4853;
   wire FE_PHN3615_n4746;
   wire FE_PHN3612_n5731;
   wire FE_PHN3611_n288;
   wire FE_PHN3610_n5725;
   wire FE_PHN3609_n5327;
   wire FE_PHN3608_n5784;
   wire FE_PHN3606_U98_Z_0;
   wire FE_PHN3605_n5402;
   wire FE_PHN3604_n5730;
   wire FE_PHN3603_n5583;
   wire FE_PHN3602_n4829;
   wire FE_PHN3601_n5094;
   wire FE_PHN3599_n5377;
   wire FE_PHN3598_n5500;
   wire FE_PHN3597_U721_Z_0;
   wire FE_PHN3596_n5145;
   wire FE_PHN3595_n5720;
   wire FE_PHN3594_n5330;
   wire FE_PHN3593_n5269;
   wire FE_PHN3592_n5714;
   wire FE_PHN3591_n5726;
   wire FE_PHN3590_n5588;
   wire FE_PHN3589_n5059;
   wire FE_PHN3587_n5359;
   wire FE_PHN3586_n5293;
   wire FE_PHN3585_n5734;
   wire FE_PHN3584_n4990;
   wire FE_PHN3583_n4980;
   wire FE_PHN3582_U453_Z_0;
   wire FE_PHN3581_n5032;
   wire FE_PHN3580_n5148;
   wire FE_PHN3578_n5406;
   wire FE_PHN3577_n5295;
   wire FE_PHN3576_U97_Z_0;
   wire FE_PHN3574_n5587;
   wire FE_PHN3573_U320_Z_0;
   wire FE_PHN3572_n5590;
   wire FE_PHN3571_n5223;
   wire FE_PHN3570_n5222;
   wire FE_PHN3569_n5282;
   wire FE_PHN3568_n5556;
   wire FE_PHN3567_n5342;
   wire FE_PHN3566_n5031;
   wire FE_PHN3565_n5404;
   wire FE_PHN3564_n5375;
   wire FE_PHN3563_n5482;
   wire FE_PHN3562_n5371;
   wire FE_PHN3561_U630_Z_0;
   wire FE_PHN3560_n5303;
   wire FE_PHN3559_n5373;
   wire FE_PHN3558_n5591;
   wire FE_PHN3557_n5274;
   wire FE_PHN3556_n5206;
   wire FE_PHN3555_n5281;
   wire FE_PHN3554_n5060;
   wire FE_PHN3553_n5647;
   wire FE_PHN3552_U246_Z_0;
   wire FE_PHN3551_n5593;
   wire FE_PHN3550_n5417;
   wire FE_PHN3548_U627_Z_0;
   wire FE_PHN3547_n5728;
   wire FE_PHN3546_U319_Z_0;
   wire FE_PHN3545_U586_Z_0;
   wire FE_PHN3544_n5716;
   wire FE_PHN3542_U597_Z_0;
   wire FE_PHN3541_U519_Z_0;
   wire FE_PHN3540_U235_Z_0;
   wire FE_PHN3539_U321_Z_0;
   wire FE_PHN3538_U632_Z_0;
   wire FE_PHN3537_U591_Z_0;
   wire FE_PHN3536_n4938;
   wire FE_PHN3535_U247_Z_0;
   wire FE_PHN3534_n4924;
   wire FE_PHN3533_U583_Z_0;
   wire FE_PHN3532_U528_Z_0;
   wire FE_PHN3531_U595_Z_0;
   wire FE_PHN3530_U589_Z_0;
   wire FE_PHN3529_U309_Z_0;
   wire FE_PHN3528_U557_Z_0;
   wire FE_PHN3527_U305_Z_0;
   wire FE_PHN3526_U566_Z_0;
   wire FE_PHN3525_U324_Z_0;
   wire FE_PHN3524_U563_Z_0;
   wire FE_PHN3523_U318_Z_0;
   wire FE_PHN3522_U323_Z_0;
   wire FE_PHN3521_n4937;
   wire FE_PHN3520_n4925;
   wire FE_PHN3519_n4935;
   wire FE_PHN3518_n4936;
   wire FE_PHN3517_n4926;
   wire FE_PHN3516_n4942;
   wire FE_PHN3512_n5510;
   wire FE_PHN3506_U795_Z_0;
   wire FE_PHN3502_U755_Z_0;
   wire FE_PHN3501_n5516;
   wire FE_PHN3500_n5099;
   wire FE_PHN3497_n5792;
   wire FE_PHN3496_n262;
   wire FE_PHN3482_n5711;
   wire FE_PHN3478_n5793;
   wire FE_PHN3477_n5790;
   wire FE_PHN3474_n5689;
   wire FE_PHN3472_n5826;
   wire FE_PHN3470_n5795;
   wire FE_PHN3466_n214;
   wire FE_PHN3437_n5783;
   wire FE_PHN3421_n5684;
   wire FE_PHN3414_n5679;
   wire FE_PHN3411_n222;
   wire FE_PHN3405_n5677;
   wire FE_PHN3391_n5673;
   wire FE_PHN3387_n5655;
   wire FE_PHN3377_n5682;
   wire FE_PHN3375_n5676;
   wire FE_PHN3353_n5675;
   wire FE_PHN3290_n4923;
   wire FE_PHN3282_n5685;
   wire FE_PHN3278_n4934;
   wire FE_PHN3277_n4939;
   wire FE_PHN3276_n4930;
   wire FE_PHN3275_n4928;
   wire FE_PHN3274_n4933;
   wire FE_PHN3273_n5800;
   wire FE_PHN3217_n5736;
   wire FE_PHN3211_U229_Z_0;
   wire FE_PHN3209_n5791;
   wire FE_PHN3206_n5712;
   wire FE_PHN3205_n5827;
   wire FE_PHN3204_n13813;
   wire FE_PHN3202_n13951;
   wire FE_PHN3201_n13870;
   wire FE_PHN3200_n5763;
   wire FE_PHN3199_n5756;
   wire FE_PHN3198_n5767;
   wire FE_PHN3190_n4931;
   wire FE_PHN3153_n5668;
   wire FE_PHN3143_U227_Z_0;
   wire FE_PHN3142_n5765;
   wire FE_PHN3140_n4921;
   wire FE_PHN3139_n5755;
   wire FE_PHN3138_n5758;
   wire FE_PHN3137_n4910;
   wire FE_PHN3136_n4907;
   wire FE_PHN3135_n4914;
   wire FE_PHN3134_n5762;
   wire FE_PHN3133_n14432;
   wire FE_PHN3103_n4847;
   wire FE_PHN3102_n5237;
   wire FE_PHN3101_n5235;
   wire FE_PHN3100_n5573;
   wire FE_PHN3099_n5601;
   wire FE_PHN3098_n5238;
   wire FE_PHN3097_n5236;
   wire FE_PHN3094_n5761;
   wire FE_PHN3093_n4918;
   wire FE_PHN3092_n14001;
   wire FE_PHN3091_n5768;
   wire FE_PHN3090_n5751;
   wire FE_PHN3089_n5754;
   wire FE_PHN3088_n5744;
   wire FE_PHN3084_n5658;
   wire FE_PHN3078_n5729;
   wire FE_PHN3076_U692_Z_0;
   wire FE_PHN3074_n5798;
   wire FE_PHN3073_n5782;
   wire FE_PHN3072_n5788;
   wire FE_PHN3071_n5717;
   wire FE_PHN3070_n4879;
   wire FE_PHN3069_n4945;
   wire FE_PHN3068_n13795;
   wire FE_PHN3067_n13989;
   wire FE_PHN3066_n13963;
   wire FE_PHN3065_n13932;
   wire FE_PHN3064_n13835;
   wire FE_PHN3063_n13919;
   wire FE_PHN3061_n13894;
   wire FE_PHN3060_n14956;
   wire FE_PHN3059_n13907;
   wire FE_PHN3058_n13758;
   wire FE_PHN3057_n5769;
   wire FE_PHN3056_n5748;
   wire FE_PHN3055_n166;
   wire FE_PHN3050_n5713;
   wire FE_PHN3048_n11928;
   wire FE_PHN3018_IRQ_14_;
   wire FE_PHN3001_n4895;
   wire FE_PHN3000_n419;
   wire FE_PHN2995_IRQ_8_;
   wire FE_PHN2994_IRQ_11_;
   wire FE_PHN2993_IRQ_13_;
   wire FE_PHN2992_IRQ_2_;
   wire FE_PHN2991_IRQ_3_;
   wire FE_PHN2990_IRQ_7_;
   wire FE_PHN2989_IRQ_10_;
   wire FE_PHN2988_IRQ_9_;
   wire FE_PHN2987_IRQ_6_;
   wire FE_PHN2986_IRQ_4_;
   wire FE_PHN2985_IRQ_0_;
   wire FE_PHN2984_IRQ_5_;
   wire FE_PHN2983_IRQ_1_;
   wire FE_PHN2982_NMI;
   wire FE_PHN2981_n5760;
   wire FE_PHN2980_IRQ_15_;
   wire FE_PHN2976_n5656;
   wire FE_PHN2974_n5757;
   wire FE_PHN2973_n4908;
   wire FE_PHN2972_n5759;
   wire FE_PHN2970_n1444;
   wire FE_PHN2969_n4917;
   wire FE_PHN2968_n4919;
   wire FE_PHN2967_n4920;
   wire FE_PHN2966_n5766;
   wire FE_PHN2965_n5750;
   wire FE_PHN2955_n5741;
   wire FE_PHN2954_n5753;
   wire FE_PHN2953_n5739;
   wire FE_PHN2952_n5740;
   wire FE_PHN2951_n4916;
   wire FE_PHN2948_n5752;
   wire FE_PHN2947_n4911;
   wire FE_PHN2946_n4913;
   wire FE_PHN2945_n4906;
   wire FE_PHN2944_n4909;
   wire FE_PHN2943_n4912;
   wire FE_PHN2939_n4915;
   wire FE_PHN2936_n5746;
   wire FE_PHN2935_n5745;
   wire FE_PHN2928_n1145;
   wire FE_PHN2927_n5692;
   wire FE_PHN2926_n5683;
   wire FE_PHN2922_n5747;
   wire FE_PHN2921_n5749;
   wire FE_PHN2920_n5743;
   wire FE_PHN2918_n5742;
   wire FE_PHN2916_n171;
   wire FE_PHN2912_n17127;
   wire FE_PHN2911_n17126;
   wire FE_PHN2903_n5707;
   wire FE_PHN2902_n5703;
   wire FE_PHN2901_n5706;
   wire FE_PHN2900_n5702;
   wire FE_PHN2899_n5799;
   wire FE_PHN2898_n5710;
   wire FE_PHN2897_U763_Z_0;
   wire FE_PHN2896_U762_Z_0;
   wire FE_PHN2895_U774_Z_0;
   wire FE_PHN2894_U781_Z_0;
   wire FE_PHN2893_U789_Z_0;
   wire FE_PHN2892_n5704;
   wire FE_PHN2891_n5651;
   wire FE_PHN2890_U791_Z_0;
   wire FE_PHN2889_n4862;
   wire FE_PHN2888_n5705;
   wire FE_PHN2887_U771_Z_0;
   wire FE_PHN2886_U782_Z_0;
   wire FE_PHN2885_U783_Z_0;
   wire FE_PHN2884_U772_Z_0;
   wire FE_PHN2883_U353_Z_0;
   wire FE_PHN2882_U775_Z_0;
   wire FE_PHN2881_U788_Z_0;
   wire FE_PHN2879_U441_Z_0;
   wire FE_PHN2878_U787_Z_0;
   wire FE_PHN2877_U786_Z_0;
   wire FE_PHN2875_U770_Z_0;
   wire FE_PHN2874_U764_Z_0;
   wire FE_PHN2873_U459_Z_0;
   wire FE_PHN2872_U261_Z_0;
   wire FE_PHN2871_U363_Z_0;
   wire FE_PHN2870_U780_Z_0;
   wire FE_PHN2869_U279_Z_0;
   wire FE_PHN2868_U425_Z_0;
   wire FE_PHN2867_U800_Z_0;
   wire FE_PHN2866_U479_Z_0;
   wire FE_PHN2865_n4854;
   wire FE_PHN2864_U429_Z_0;
   wire FE_PHN2863_U606_Z_0;
   wire FE_PHN2862_U513_Z_0;
   wire FE_PHN2861_U275_Z_0;
   wire FE_PHN2860_U667_Z_0;
   wire FE_PHN2859_U726_Z_0;
   wire FE_PHN2858_U359_Z_0;
   wire FE_PHN2857_U766_Z_0;
   wire FE_PHN2856_U395_Z_0;
   wire FE_PHN2855_U497_Z_0;
   wire FE_PHN2854_U509_Z_0;
   wire FE_PHN2853_U506_Z_0;
   wire FE_PHN2852_U660_Z_0;
   wire FE_PHN2851_U448_Z_0;
   wire FE_PHN2849_U761_Z_0;
   wire FE_PHN2848_U411_Z_0;
   wire FE_PHN2847_U475_Z_0;
   wire FE_PHN2846_U407_Z_0;
   wire FE_PHN2845_U673_Z_0;
   wire FE_PHN2844_U610_Z_0;
   wire FE_PHN2843_U291_Z_0;
   wire FE_PHN2842_U463_Z_0;
   wire FE_PHN2841_U777_Z_0;
   wire FE_PHN2839_U801_Z_0;
   wire FE_PHN2838_U493_Z_0;
   wire FE_PHN2837_U785_Z_0;
   wire FE_PHN2836_U257_Z_0;
   wire FE_PHN2835_U466_Z_0;
   wire FE_PHN2834_U712_Z_0;
   wire FE_PHN2833_U727_Z_0;
   wire FE_PHN2832_U784_Z_0;
   wire FE_PHN2831_U644_Z_0;
   wire FE_PHN2830_U711_Z_0;
   wire FE_PHN2829_U295_Z_0;
   wire FE_PHN2828_U386_Z_0;
   wire FE_PHN2827_U503_Z_0;
   wire FE_PHN2826_n5097;
   wire FE_PHN2824_U428_Z_0;
   wire FE_PHN2823_U263_Z_0;
   wire FE_PHN2822_U504_Z_0;
   wire FE_PHN2821_U677_Z_0;
   wire FE_PHN2820_U646_Z_0;
   wire FE_PHN2819_U471_Z_0;
   wire FE_PHN2818_n5650;
   wire FE_PHN2817_U779_Z_0;
   wire FE_PHN2816_U721_Z_0;
   wire FE_PHN2815_U490_Z_0;
   wire FE_PHN2814_U612_Z_0;
   wire FE_PHN2813_U391_Z_0;
   wire FE_PHN2812_U683_Z_0;
   wire FE_PHN2811_U728_Z_0;
   wire FE_PHN2810_U663_Z_0;
   wire FE_PHN2809_U445_Z_0;
   wire FE_PHN2808_U651_Z_0;
   wire FE_PHN2807_U745_Z_0;
   wire FE_PHN2806_U680_Z_0;
   wire FE_PHN2805_U454_Z_0;
   wire FE_PHN2804_U743_Z_0;
   wire FE_PHN2803_U769_Z_0;
   wire FE_PHN2802_U496_Z_0;
   wire FE_PHN2801_n5457;
   wire FE_PHN2800_U453_Z_0;
   wire FE_PHN2799_U708_Z_0;
   wire FE_PHN2798_U748_Z_0;
   wire FE_PHN2796_n5267;
   wire FE_PHN2795_U481_Z_0;
   wire FE_PHN2794_U500_Z_0;
   wire FE_PHN2793_U656_Z_0;
   wire FE_PHN2792_U634_Z_0;
   wire FE_PHN2791_n5297;
   wire FE_PHN2790_n5284;
   wire FE_PHN2789_n5130;
   wire FE_PHN2788_n5062;
   wire FE_PHN2787_n5603;
   wire FE_PHN2786_n5072;
   wire FE_PHN2785_n5288;
   wire FE_PHN2784_n5568;
   wire FE_PHN2783_n5622;
   wire FE_PHN2782_n5487;
   wire FE_PHN2781_n5169;
   wire FE_PHN2780_n5612;
   wire FE_PHN2779_n5604;
   wire FE_PHN2778_n5075;
   wire FE_PHN2777_n5557;
   wire FE_PHN2776_n5141;
   wire FE_PHN2775_n5470;
   wire FE_PHN2774_n5083;
   wire FE_PHN2773_n5170;
   wire FE_PHN2772_n5172;
   wire FE_PHN2771_n5468;
   wire FE_PHN2770_n5178;
   wire FE_PHN2769_n5299;
   wire FE_PHN2768_n5478;
   wire FE_PHN2767_n5450;
   wire FE_PHN2766_n5186;
   wire FE_PHN2765_n5039;
   wire FE_PHN2764_n5173;
   wire FE_PHN2763_n5196;
   wire FE_PHN2762_n5174;
   wire FE_PHN2761_n5472;
   wire FE_PHN2760_n5455;
   wire FE_PHN2759_n5396;
   wire FE_PHN2758_n5296;
   wire FE_PHN2757_n5641;
   wire FE_PHN2756_n4985;
   wire FE_PHN2755_n5461;
   wire FE_PHN2754_n5633;
   wire FE_PHN2753_n5553;
   wire FE_PHN2752_n5187;
   wire FE_PHN2751_n4969;
   wire FE_PHN2750_n5015;
   wire FE_PHN2749_n5598;
   wire FE_PHN2748_n5312;
   wire FE_PHN2747_n5437;
   wire FE_PHN2746_n5428;
   wire FE_PHN2745_n5426;
   wire FE_PHN2744_n5486;
   wire FE_PHN2743_n5597;
   wire FE_PHN2742_n5121;
   wire FE_PHN2741_n5040;
   wire FE_PHN2740_n5420;
   wire FE_PHN2739_n5161;
   wire FE_PHN2738_n5469;
   wire FE_PHN2737_n5135;
   wire FE_PHN2736_n5103;
   wire FE_PHN2735_n5021;
   wire FE_PHN2734_n5464;
   wire FE_PHN2733_n5616;
   wire FE_PHN2732_n5636;
   wire FE_PHN2731_n5138;
   wire FE_PHN2730_n5046;
   wire FE_PHN2729_n5463;
   wire FE_PHN2728_n5115;
   wire FE_PHN2727_n5086;
   wire FE_PHN2726_n5022;
   wire FE_PHN2725_n5392;
   wire FE_PHN2724_n5477;
   wire FE_PHN2723_n5485;
   wire FE_PHN2722_n5012;
   wire FE_PHN2721_n5433;
   wire FE_PHN2720_n5020;
   wire FE_PHN2719_n5181;
   wire FE_PHN2718_n5300;
   wire FE_PHN2717_n5438;
   wire FE_PHN2716_n5366;
   wire FE_PHN2715_n5397;
   wire FE_PHN2714_n5442;
   wire FE_PHN2713_n5171;
   wire FE_PHN2712_n5287;
   wire FE_PHN2711_n5453;
   wire FE_PHN2710_n5427;
   wire FE_PHN2709_n5564;
   wire FE_PHN2708_n5452;
   wire FE_PHN2707_n5459;
   wire FE_PHN2706_n5575;
   wire FE_PHN2705_n5432;
   wire FE_PHN2703_n5197;
   wire FE_PHN2702_n5449;
   wire FE_PHN2701_n5430;
   wire FE_PHN2700_n5069;
   wire FE_PHN2699_n5462;
   wire FE_PHN2698_n5439;
   wire FE_PHN2697_n5184;
   wire FE_PHN2696_n5424;
   wire FE_PHN2695_n5401;
   wire FE_PHN2694_n5466;
   wire FE_PHN2693_n5190;
   wire FE_PHN2692_n5398;
   wire FE_PHN2691_n5550;
   wire FE_PHN2690_n5051;
   wire FE_PHN2689_n5043;
   wire FE_PHN2688_n5421;
   wire FE_PHN2687_n5175;
   wire FE_PHN2686_n5576;
   wire FE_PHN2685_n5030;
   wire FE_PHN2684_n5010;
   wire FE_PHN2683_n5191;
   wire FE_PHN2682_n5447;
   wire FE_PHN2681_n5108;
   wire FE_PHN2680_n5041;
   wire FE_PHN2679_n5123;
   wire FE_PHN2678_n5606;
   wire FE_PHN2676_n4987;
   wire FE_PHN2675_n5539;
   wire FE_PHN2674_n5476;
   wire FE_PHN2673_n5091;
   wire FE_PHN2672_n5538;
   wire FE_PHN2671_n5473;
   wire FE_PHN2670_n5192;
   wire FE_PHN2669_n5434;
   wire FE_PHN2668_n5444;
   wire FE_PHN2667_n5183;
   wire FE_PHN2666_n5106;
   wire FE_PHN2665_n5410;
   wire FE_PHN2664_n5093;
   wire FE_PHN2663_n5195;
   wire FE_PHN2662_n5132;
   wire FE_PHN2661_n5304;
   wire FE_PHN2660_n5567;
   wire FE_PHN2659_n5435;
   wire FE_PHN2658_n5448;
   wire FE_PHN2657_n5399;
   wire FE_PHN2655_n5393;
   wire FE_PHN2654_n5411;
   wire FE_PHN2653_n5451;
   wire FE_PHN2652_n5298;
   wire FE_PHN2651_n5412;
   wire FE_PHN2650_n5289;
   wire FE_PHN2649_n5182;
   wire FE_PHN2648_n4986;
   wire FE_PHN2647_n5189;
   wire FE_PHN2646_n5440;
   wire FE_PHN2645_n5301;
   wire FE_PHN2644_n5558;
   wire FE_PHN2643_n5180;
   wire FE_PHN2642_n5414;
   wire FE_PHN2641_n5441;
   wire FE_PHN2640_n5418;
   wire FE_PHN2639_n5643;
   wire FE_PHN2637_n5395;
   wire FE_PHN2636_n5363;
   wire FE_PHN2635_n5207;
   wire FE_PHN2634_n5028;
   wire FE_PHN2633_n5176;
   wire FE_PHN2632_n5419;
   wire FE_PHN2631_n5203;
   wire FE_PHN2630_n5629;
   wire FE_PHN2629_n5409;
   wire FE_PHN2628_n5348;
   wire FE_PHN2627_n5013;
   wire FE_PHN2626_n5360;
   wire FE_PHN2625_n5266;
   wire FE_PHN2624_n5415;
   wire FE_PHN2623_n5159;
   wire FE_PHN2622_n5483;
   wire FE_PHN2621_n5521;
   wire FE_PHN2620_n5367;
   wire FE_PHN2619_n5273;
   wire FE_PHN2618_n5596;
   wire FE_PHN2617_n5481;
   wire FE_PHN2616_n5205;
   wire FE_PHN2615_n5045;
   wire FE_PHN2614_n4979;
   wire FE_PHN2613_n5270;
   wire FE_PHN2612_n5199;
   wire FE_PHN2611_n5436;
   wire FE_PHN2610_n5308;
   wire FE_PHN2609_n5112;
   wire FE_PHN2608_n5624;
   wire FE_PHN2607_n5076;
   wire FE_PHN2606_n5364;
   wire FE_PHN2605_n5384;
   wire FE_PHN2604_n5309;
   wire FE_PHN2603_n5343;
   wire FE_PHN2602_n5386;
   wire FE_PHN2601_n5413;
   wire FE_PHN2600_n5362;
   wire FE_PHN2599_n5361;
   wire FE_PHN2598_n5224;
   wire FE_PHN2597_n5422;
   wire FE_PHN2596_n5261;
   wire FE_PHN2595_n5357;
   wire FE_PHN2594_n5443;
   wire FE_PHN2593_n5638;
   wire FE_PHN2592_n5219;
   wire FE_PHN2591_n5394;
   wire FE_PHN2590_n5554;
   wire FE_PHN2589_n5081;
   wire FE_PHN2588_n5225;
   wire FE_PHN2587_n5374;
   wire FE_PHN2586_n5049;
   wire FE_PHN2585_n4995;
   wire FE_PHN2584_n5202;
   wire FE_PHN2583_n5070;
   wire FE_PHN2582_n5403;
   wire FE_PHN2581_n5107;
   wire FE_PHN2580_n5271;
   wire FE_PHN2579_n5128;
   wire FE_PHN2578_n5125;
   wire FE_PHN2577_n5079;
   wire FE_PHN2576_n5201;
   wire FE_PHN2574_n5019;
   wire FE_PHN2573_n5405;
   wire FE_PHN2572_n5365;
   wire FE_PHN2571_n5355;
   wire FE_PHN2570_n5479;
   wire FE_PHN2569_n5136;
   wire FE_PHN2568_n5200;
   wire FE_PHN2566_n5336;
   wire FE_PHN2564_n5319;
   wire FE_PHN2563_n5372;
   wire FE_PHN2562_n5278;
   wire FE_PHN2561_n5139;
   wire FE_PHN2560_n5560;
   wire FE_PHN2559_n5368;
   wire FE_PHN2557_n5369;
   wire FE_PHN2556_n5640;
   wire FE_PHN2555_n5335;
   wire FE_PHN2554_n5316;
   wire FE_PHN2553_n5218;
   wire FE_PHN2552_n5562;
   wire FE_PHN2551_n5268;
   wire FE_PHN2550_n5131;
   wire FE_PHN2549_n5334;
   wire FE_PHN2548_n5213;
   wire FE_PHN2547_n5383;
   wire FE_PHN2546_n5018;
   wire FE_PHN2545_n5317;
   wire FE_PHN2544_n5621;
   wire FE_PHN2543_n5217;
   wire FE_PHN2542_n5491;
   wire FE_PHN2541_n5356;
   wire FE_PHN2540_n5063;
   wire FE_PHN2539_n5347;
   wire FE_PHN2538_n5109;
   wire FE_PHN2537_n5211;
   wire FE_PHN2536_n5209;
   wire FE_PHN2535_n5339;
   wire FE_PHN2534_n5630;
   wire FE_PHN2533_n5349;
   wire FE_PHN2532_n5376;
   wire FE_PHN2531_n5566;
   wire FE_PHN2530_n5133;
   wire FE_PHN2529_n5634;
   wire FE_PHN2528_n5283;
   wire FE_PHN2527_n5279;
   wire FE_PHN2526_n5044;
   wire FE_PHN2525_n5381;
   wire FE_PHN2524_n5292;
   wire FE_PHN2523_n5563;
   wire FE_PHN2522_n5378;
   wire FE_PHN2521_n5263;
   wire FE_PHN2520_n5212;
   wire FE_PHN2519_n5221;
   wire FE_PHN2518_n5543;
   wire FE_PHN2517_n5220;
   wire FE_PHN2516_n5542;
   wire FE_PHN2515_n5617;
   wire FE_PHN2514_n5610;
   wire FE_PHN2513_n5280;
   wire FE_PHN2512_n5391;
   wire FE_PHN2511_n5104;
   wire FE_PHN2510_n5599;
   wire FE_PHN2509_n5124;
   wire FE_PHN2508_n5264;
   wire FE_PHN2507_n5084;
   wire FE_PHN2506_n5480;
   wire FE_PHN2505_n5385;
   wire FE_PHN2504_n5337;
   wire FE_PHN2503_n5497;
   wire FE_PHN2502_n5037;
   wire FE_PHN2501_n4984;
   wire FE_PHN2500_n5216;
   wire FE_PHN2499_n5142;
   wire FE_PHN2498_n5350;
   wire FE_PHN2497_n5602;
   wire FE_PHN2496_n5052;
   wire FE_PHN2495_n5042;
   wire FE_PHN2494_n5489;
   wire FE_PHN2493_n5198;
   wire FE_PHN2492_n5611;
   wire FE_PHN2491_n5066;
   wire FE_PHN2490_n5294;
   wire FE_PHN2489_n5087;
   wire FE_PHN2488_n4998;
   wire FE_PHN2487_n5607;
   wire FE_PHN2486_n5276;
   wire FE_PHN2485_n5379;
   wire FE_PHN2484_n5574;
   wire FE_PHN2483_n5226;
   wire FE_PHN2482_n5352;
   wire FE_PHN2481_n5277;
   wire FE_PHN2480_n5494;
   wire FE_PHN2479_n5116;
   wire FE_PHN2478_n5631;
   wire FE_PHN2477_n5380;
   wire FE_PHN2476_n5548;
   wire FE_PHN2475_n5215;
   wire FE_PHN2474_n5214;
   wire FE_PHN2473_n5092;
   wire FE_PHN2472_n5122;
   wire FE_PHN2471_n5089;
   wire FE_PHN2470_n5382;
   wire FE_PHN2469_n5351;
   wire FE_PHN2468_n5260;
   wire FE_PHN2467_n5492;
   wire FE_PHN2466_n5493;
   wire FE_PHN2465_n5559;
   wire FE_PHN2464_n5318;
   wire FE_PHN2463_n5354;
   wire FE_PHN2462_n5627;
   wire FE_PHN2461_n5490;
   wire FE_PHN2460_n5286;
   wire FE_PHN2459_n5608;
   wire FE_PHN2458_n5353;
   wire FE_PHN2457_n5635;
   wire FE_PHN2456_n5496;
   wire FE_PHN2454_n5345;
   wire FE_PHN2453_n5541;
   wire FE_PHN2452_n5569;
   wire FE_PHN2451_n4963;
   wire FE_PHN2450_n5341;
   wire FE_PHN2449_n5370;
   wire FE_PHN2448_n5614;
   wire FE_PHN2447_n5275;
   wire FE_PHN2446_n5262;
   wire FE_PHN2445_n5016;
   wire FE_PHN2444_n5390;
   wire FE_PHN2443_n5389;
   wire FE_PHN2442_n5495;
   wire FE_PHN2441_n5210;
   wire FE_PHN2440_n5307;
   wire FE_PHN2439_n5340;
   wire FE_PHN2438_n5073;
   wire FE_PHN2437_n5204;
   wire FE_PHN2436_n5577;
   wire FE_PHN2435_n5265;
   wire FE_PHN2430_n5520;
   wire FE_PHN2429_n5505;
   wire FE_PHN2428_n5507;
   wire FE_PHN2426_n5581;
   wire FE_PHN2420_n5652;
   wire FE_PHN2415_n5792;
   wire FE_PHN2412_n5512;
   wire FE_PHN2403_n5711;
   wire FE_PHN2385_n5625;
   wire FE_PHN2379_n5793;
   wire FE_PHN2378_n5618;
   wire FE_PHN2376_n5571;
   wire FE_PHN2364_n5639;
   wire FE_PHN2355_U594_Z_0;
   wire FE_PHN2348_n5790;
   wire FE_PHN2347_n5513;
   wire FE_PHN2346_U243_Z_0;
   wire FE_PHN2333_n5600;
   wire FE_PHN2330_n5579;
   wire FE_PHN2302_n5509;
   wire FE_PHN2300_U239_Z_0;
   wire FE_PHN2294_U325_Z_0;
   wire FE_PHN2286_U329_Z_0;
   wire FE_PHN2270_n5067;
   wire FE_PHN2254_n5074;
   wire FE_PHN2245_n5033;
   wire FE_PHN2241_U234_Z_0;
   wire FE_PHN2240_n5514;
   wire FE_PHN2233_U624_Z_0;
   wire FE_PHN2232_n5511;
   wire FE_PHN2225_U619_Z_0;
   wire FE_PHN2224_U628_Z_0;
   wire FE_PHN2223_n5508;
   wire FE_PHN2219_U585_Z_0;
   wire FE_PHN2215_U242_Z_0;
   wire FE_PHN2212_U233_Z_0;
   wire FE_PHN2210_U320_Z_0;
   wire FE_PHN2200_U593_Z_0;
   wire FE_PHN2196_U245_Z_0;
   wire FE_PHN2189_U620_Z_0;
   wire FE_PHN2187_U618_Z_0;
   wire FE_PHN2181_U584_Z_0;
   wire FE_PHN2180_n5517;
   wire FE_PHN2179_U627_Z_0;
   wire FE_PHN2166_U596_Z_0;
   wire FE_PHN2164_n4863;
   wire FE_PHN2163_U332_Z_0;
   wire FE_PHN2157_U328_Z_0;
   wire FE_PHN2156_U311_Z_0;
   wire FE_PHN2154_U302_Z_0;
   wire FE_PHN2150_U310_Z_0;
   wire FE_PHN2149_U621_Z_0;
   wire FE_PHN2148_U597_Z_0;
   wire FE_PHN2145_U303_Z_0;
   wire FE_PHN2143_U631_Z_0;
   wire FE_PHN2141_U301_Z_0;
   wire FE_PHN2140_n5515;
   wire FE_PHN2125_U236_Z_0;
   wire FE_PHN2120_U322_Z_0;
   wire FE_PHN2114_U586_Z_0;
   wire FE_PHN2109_U235_Z_0;
   wire FE_PHN2107_U300_Z_0;
   wire FE_PHN2106_n5506;
   wire FE_PHN2105_U519_Z_0;
   wire FE_PHN2104_U524_Z_0;
   wire FE_PHN2103_U314_Z_0;
   wire FE_PHN2102_U331_Z_0;
   wire FE_PHN2101_U246_Z_0;
   wire FE_PHN2100_U592_Z_0;
   wire FE_PHN2099_U321_Z_0;
   wire FE_PHN2098_U587_Z_0;
   wire FE_PHN2097_U626_Z_0;
   wire FE_PHN2096_U326_Z_0;
   wire FE_PHN2095_U629_Z_0;
   wire FE_PHN2094_U306_Z_0;
   wire FE_PHN2093_U632_Z_0;
   wire FE_PHN2092_U534_Z_0;
   wire FE_PHN2091_U232_Z_0;
   wire FE_PHN2090_U307_Z_0;
   wire FE_PHN2089_U565_Z_0;
   wire FE_PHN2088_U583_Z_0;
   wire FE_PHN2087_U617_Z_0;
   wire FE_PHN2086_n4882;
   wire FE_PHN2085_U591_Z_0;
   wire FE_PHN2084_U238_Z_0;
   wire FE_PHN2083_U327_Z_0;
   wire FE_PHN2082_U532_Z_0;
   wire FE_PHN2081_U623_Z_0;
   wire FE_PHN2080_U622_Z_0;
   wire FE_PHN2079_U523_Z_0;
   wire FE_PHN2078_U312_Z_0;
   wire FE_PHN2077_U555_Z_0;
   wire FE_PHN2076_U564_Z_0;
   wire FE_PHN2075_U333_Z_0;
   wire FE_PHN2074_U557_Z_0;
   wire FE_PHN2073_U240_Z_0;
   wire FE_PHN2072_U324_Z_0;
   wire FE_PHN2071_U237_Z_0;
   wire FE_PHN2070_U625_Z_0;
   wire FE_PHN2069_U589_Z_0;
   wire FE_PHN2068_U330_Z_0;
   wire FE_PHN2067_U588_Z_0;
   wire FE_PHN2066_U305_Z_0;
   wire FE_PHN2065_U556_Z_0;
   wire FE_PHN2064_U308_Z_0;
   wire FE_PHN2063_U598_Z_0;
   wire FE_PHN2062_U595_Z_0;
   wire FE_PHN2061_U304_Z_0;
   wire FE_PHN2060_U318_Z_0;
   wire FE_PHN2059_U563_Z_0;
   wire FE_PHN2058_U309_Z_0;
   wire FE_PHN2057_U528_Z_0;
   wire FE_PHN2056_U323_Z_0;
   wire FE_PHN2055_U241_Z_0;
   wire FE_PHN2054_U533_Z_0;
   wire FE_PHN2053_U315_Z_0;
   wire FE_PHN2052_U244_Z_0;
   wire FE_PHN2050_n5694;
   wire FE_PHN2049_n222;
   wire FE_PHN2048_n227;
   wire FE_PHN2047_n216;
   wire FE_PHN2046_n5699;
   wire FE_PHN2045_n1000;
   wire FE_PHN2043_n230;
   wire FE_PHN2042_n1051;
   wire FE_PHN2041_n220;
   wire FE_PHN2039_U144_Z_0;
   wire FE_PHN2035_n214;
   wire FE_PHN2028_n5776;
   wire FE_PHN1983_n4923;
   wire FE_PHN1978_n4938;
   wire FE_PHN1970_U754_Z_0;
   wire FE_PHN1967_U122_Z_0;
   wire FE_PHN1934_n4924;
   wire FE_PHN1920_n4935;
   wire FE_PHN1919_n5712;
   wire FE_PHN1915_n4936;
   wire FE_PHN1914_n4942;
   wire FE_PHN1912_n4926;
   wire FE_PHN1910_n4937;
   wire FE_PHN1909_n4931;
   wire FE_PHN1908_n4925;
   wire FE_PHN1906_n5800;
   wire FE_PHN1905_n5828;
   wire FE_PHN1903_n5795;
   wire FE_PHN1902_n4903;
   wire FE_PHN1901_n4902;
   wire FE_PHN1900_n4324;
   wire FE_PHN1899_n4326;
   wire FE_PHN1898_U317_Z_0;
   wire FE_PHN1894_n5149;
   wire FE_PHN1875_n5653;
   wire FE_PHN1846_U590_Z_0;
   wire FE_PHN1809_n4874;
   wire FE_PHN1759_U630_Z_0;
   wire FE_PHN1751_U319_Z_0;
   wire FE_PHN1748_n5510;
   wire FE_PHN1744_U531_Z_0;
   wire FE_PHN1743_U313_Z_0;
   wire FE_PHN1742_U566_Z_0;
   wire FE_PHN1741_U247_Z_0;
   wire FE_PHN1717_n5114;
   wire FE_PHN1682_n16735;
   wire FE_PHN1674_n13951;
   wire FE_PHN1673_n14956;
   wire FE_PHN1672_n13963;
   wire FE_PHN1671_n13870;
   wire FE_PHN1670_n13932;
   wire FE_PHN1669_n13894;
   wire FE_PHN1668_n4389;
   wire FE_PHN1667_n13989;
   wire FE_PHN1666_n13919;
   wire FE_PHN1665_n1127;
   wire FE_PHN1664_n13747;
   wire FE_PHN1657_n5779;
   wire FE_PHN1655_n4860;
   wire FE_PHN1654_U105_Z_0;
   wire FE_PHN1653_U802_Z_0;
   wire FE_PHN1652_U134_Z_0;
   wire FE_PHN1651_U121_Z_0;
   wire FE_PHN1649_U755_Z_0;
   wire FE_PHN1648_U811_Z_0;
   wire FE_PHN1646_U518_Z_0;
   wire FE_PHN1644_U795_Z_0;
   wire FE_PHN1636_n4878;
   wire FE_PHN1633_U98_Z_0;
   wire FE_PHN1632_U97_Z_0;
   wire FE_PHN1631_n4943;
   wire FE_PHN1629_n5784;
   wire FE_PHN1627_n5786;
   wire FE_PHN1626_n5736;
   wire FE_PHN1625_n4864;
   wire FE_PHN1624_n4881;
   wire FE_PHN1615_n5827;
   wire FE_PHN1614_U665_Z_0;
   wire FE_PHN1613_n5777;
   wire FE_PHN1612_n5781;
   wire FE_PHN1610_n4886;
   wire FE_PHN1606_n13795;
   wire FE_PHN1603_n13813;
   wire FE_PHN1602_n13835;
   wire FE_PHN1601_n13758;
   wire FE_PHN1600_n13907;
   wire FE_PHN1599_n1431;
   wire FE_PHN1598_n4328;
   wire FE_PHN1588_n5737;
   wire FE_PHN1586_n5256;
   wire FE_PHN1577_n5684;
   wire FE_PHN1571_n5771;
   wire FE_PHN1566_n8706;
   wire FE_PHN1565_n8698;
   wire FE_PHN1559_n5682;
   wire FE_PHN1551_n1319;
   wire FE_PHN1538_n5772;
   wire FE_PHN1512_n4331;
   wire FE_PHN1508_n10553;
   wire FE_PHN1503_IRQ_14_;
   wire FE_PHN1502_n11928;
   wire FE_PHN1501_n779;
   wire FE_PHN1500_n5785;
   wire FE_PHN1499_n5783;
   wire FE_PHN1490_n5787;
   wire FE_PHN1488_U691_Z_0;
   wire FE_PHN1472_n5738;
   wire FE_PHN1469_n4875;
   wire FE_PHN1468_n5662;
   wire FE_PHN1463_n5665;
   wire FE_PHN1462_n5660;
   wire FE_PHN1461_n4944;
   wire FE_PHN1457_n5654;
   wire FE_PHN1450_n5788;
   wire FE_PHN1448_n5782;
   wire FE_PHN1433_n5824;
   wire FE_PHN1431_n5775;
   wire FE_PHN1429_n4945;
   wire FE_PHN1428_n5789;
   wire FE_PHN1426_U227_Z_0;
   wire FE_PHN1425_n14001;
   wire FE_PHN1399_n5723;
   wire FE_PHN1398_n5727;
   wire FE_PHN1397_n5725;
   wire FE_PHN1396_n5730;
   wire FE_PHN1395_n5719;
   wire FE_PHN1394_n5721;
   wire FE_PHN1393_n5724;
   wire FE_PHN1392_n4932;
   wire FE_PHN1391_n4930;
   wire FE_PHN1390_n4876;
   wire FE_PHN1389_n4934;
   wire FE_PHN1385_n4928;
   wire FE_PHN1379_n5798;
   wire FE_PHN1377_n4879;
   wire FE_PHN1367_n4895;
   wire FE_PHN1366_IRQ_8_;
   wire FE_PHN1365_IRQ_10_;
   wire FE_PHN1364_n4896;
   wire FE_PHN1363_IRQ_4_;
   wire FE_PHN1362_n4397;
   wire FE_PHN1361_IRQ_7_;
   wire FE_PHN1360_IRQ_1_;
   wire FE_PHN1359_IRQ_13_;
   wire FE_PHN1358_n4394;
   wire FE_PHN1357_IRQ_5_;
   wire FE_PHN1356_n4336;
   wire FE_PHN1355_IRQ_0_;
   wire FE_PHN1354_n4190;
   wire FE_PHN1353_IRQ_6_;
   wire FE_PHN1352_n4391;
   wire FE_PHN1351_IRQ_11_;
   wire FE_PHN1350_IRQ_15_;
   wire FE_PHN1349_IRQ_2_;
   wire FE_PHN1348_n4300;
   wire FE_PHN1347_NMI;
   wire FE_PHN1346_IRQ_9_;
   wire FE_PHN1345_IRQ_3_;
   wire FE_PHN1344_n4193;
   wire FE_PHN1341_SYNOPSYS_UNCONNECTED_531;
   wire FE_PHN1339_SYNOPSYS_UNCONNECTED_540;
   wire FE_PHN1331_SYNOPSYS_UNCONNECTED_522;
   wire FE_PHN1320_SYNOPSYS_UNCONNECTED_518;
   wire FE_PHN1283_n5770;
   wire FE_PHN1255_n5735;
   wire FE_PHN1241_U229_Z_0;
   wire FE_PHN1237_U809_Z_0;
   wire FE_PHN1196_n5664;
   wire FE_PHN1195_n5663;
   wire FE_PHN1183_n5659;
   wire FE_PHN1177_n4929;
   wire FE_PHN1175_n4933;
   wire FE_PHN1174_n4939;
   wire FE_PHN1172_n5826;
   wire FE_PHN1164_n1444;
   wire FE_PHN1159_n5676;
   wire FE_PHN1157_n5823;
   wire FE_PHN1145_n5729;
   wire FE_PHN1142_n5733;
   wire FE_PHN1141_n5713;
   wire FE_PHN1139_n5734;
   wire FE_PHN1138_n5715;
   wire FE_PHN1137_n5732;
   wire FE_PHN1136_n5731;
   wire FE_PHN1135_n5722;
   wire FE_PHN1134_n5716;
   wire FE_PHN1133_n5728;
   wire FE_PHN1131_n5718;
   wire FE_PHN1130_n5726;
   wire FE_PHN1129_n5714;
   wire FE_PHN1128_n5717;
   wire FE_PHN1126_U692_Z_0;
   wire FE_PHN1086_n5661;
   wire FE_PHN1085_n5720;
   wire FE_PHN1078_n5668;
   wire FE_PHN1063_n5667;
   wire FE_PHN1038_n5761;
   wire FE_PHN1037_n5007;
   wire FE_PHN1025_n3063;
   wire FE_PHN1024_n5690;
   wire FE_PHN1010_n5766;
   wire FE_PHN1009_n5765;
   wire FE_PHN1008_n5767;
   wire FE_PHN1007_n5768;
   wire FE_PHN1006_n5769;
   wire FE_PHN1005_n5764;
   wire FE_PHN1004_n5673;
   wire FE_PHN1003_n5675;
   wire FE_PHN991_n5679;
   wire FE_PHN972_n5755;
   wire FE_PHN965_n5658;
   wire FE_PHN963_n5671;
   wire FE_PHN946_n5677;
   wire FE_PHN941_n5674;
   wire FE_PHN939_n5680;
   wire FE_PHN936_n5683;
   wire FE_PHN935_n2982;
   wire FE_PHN928_n14432;
   wire FE_PHN904_n393;
   wire FE_PHN892_n14928;
   wire FE_PHN875_n423;
   wire FE_PHN870_n420;
   wire FE_PHN869_n427;
   wire FE_PHN859_n2624;
   wire FE_PHN856_n5656;
   wire FE_PHN852_n5763;
   wire FE_PHN851_n4920;
   wire FE_PHN849_n4918;
   wire FE_PHN847_n4917;
   wire FE_PHN846_n4915;
   wire FE_PHN845_n4919;
   wire FE_PHN844_n425;
   wire FE_PHN839_n5678;
   wire FE_PHN830_n5760;
   wire FE_PHN829_n5756;
   wire FE_PHN826_n4921;
   wire FE_PHN825_n4913;
   wire FE_PHN824_n4908;
   wire FE_PHN823_n4914;
   wire FE_PHN822_n4910;
   wire FE_PHN821_n4911;
   wire FE_PHN820_n4916;
   wire FE_PHN819_n4909;
   wire FE_PHN818_n4912;
   wire FE_PHN813_n5670;
   wire FE_PHN806_n1143;
   wire FE_PHN804_n429;
   wire FE_PHN803_n5757;
   wire FE_PHN802_n5762;
   wire FE_PHN801_n5758;
   wire FE_PHN793_n4907;
   wire FE_PHN783_n152;
   wire FE_PHN780_n2892;
   wire FE_PHN779_n5669;
   wire FE_PHN778_n160;
   wire FE_PHN776_n1108;
   wire FE_PHN775_n5689;
   wire FE_PHN774_n14825;
   wire FE_PHN770_n140;
   wire FE_PHN769_n5685;
   wire FE_PHN768_n72;
   wire FE_PHN765_n1144;
   wire FE_PHN763_n1140;
   wire FE_PHN762_n4906;
   wire FE_PHN760_n5666;
   wire FE_PHN756_n1145;
   wire FE_PHN755_n1142;
   wire FE_PHN753_n5759;
   wire FE_PHN752_n1337;
   wire FE_PHN749_n5657;
   wire FE_PHN748_n2415;
   wire FE_PHN743_n3096;
   wire FE_PHN741_n5681;
   wire FE_PHN739_n5751;
   wire FE_PHN738_n5745;
   wire FE_PHN737_n5744;
   wire FE_PHN735_n100;
   wire FE_PHN733_n5748;
   wire FE_PHN732_n5692;
   wire FE_PHN731_n5691;
   wire FE_PHN730_n5750;
   wire FE_PHN729_n5746;
   wire FE_PHN728_n2421;
   wire FE_PHN727_n3344;
   wire FE_PHN723_n5741;
   wire FE_PHN722_n5740;
   wire FE_PHN721_n5749;
   wire FE_PHN720_n5739;
   wire FE_PHN719_n190;
   wire FE_PHN717_n5743;
   wire FE_PHN716_n5753;
   wire FE_PHN715_n5754;
   wire FE_PHN712_n5687;
   wire FE_PHN711_n28;
   wire FE_PHN707_n5747;
   wire FE_PHN705_n5655;
   wire FE_PHN704_n5752;
   wire FE_PHN703_n44;
   wire FE_PHN702_n171;
   wire FE_PHN701_n5742;
   wire FE_PHN693_n166;
   wire FE_PHN685_n2516;
   wire FE_PHN679_n2465;
   wire FE_PHN675_n17126;
   wire FE_PHN674_n17127;
   wire FE_OFN667_n17122;
   wire FE_OFN666_n17077;
   wire FE_OFN665_n17074;
   wire FE_OFN663_n17058;
   wire FE_OFN661_n17057;
   wire FE_OFN659_n17053;
   wire FE_OFN656_n17048;
   wire FE_OFN654_n17038;
   wire FE_OFN652_n17033;
   wire FE_OFN651_n17027;
   wire FE_OFN648_n17017;
   wire FE_OFN646_n16977;
   wire FE_OFN645_n16939;
   wire FE_OFN644_n16936;
   wire FE_OFN643_n16916;
   wire FE_OFN642_n16913;
   wire FE_OFN641_n16902;
   wire FE_OFN639_n16897;
   wire FE_OFN638_n16891;
   wire FE_OFN636_n16886;
   wire FE_OFN635_n16877;
   wire FE_OFN634_n16871;
   wire FE_OFN633_n16868;
   wire FE_OFN632_n16859;
   wire FE_OFN631_n16851;
   wire FE_OFN629_n16850;
   wire FE_OFN628_n16833;
   wire FE_OFN627_n16828;
   wire FE_OFN626_n16820;
   wire FE_OFN625_n16814;
   wire FE_OFN610_n16690;
   wire FE_OFN608_n16686;
   wire FE_OFN602_n16656;
   wire FE_OFN598_n5805;
   wire FE_OFN587_n5162;
   wire FE_OFN583_n5036;
   wire FE_OFN573_n4905;
   wire FE_OFN568_n4401;
   wire FE_OFN567_n4069;
   wire FE_OFN566_n4065;
   wire FE_OFN565_n4058;
   wire FE_OFN560_n3199;
   wire FE_OFN559_n3180;
   wire FE_OFN549_n2774;
   wire FE_OFN544_n2612;
   wire FE_OFN543_n2585;
   wire FE_OFN542_n2562;
   wire FE_OFN541_n2556;
   wire FE_OFN539_n2519;
   wire FE_OFN538_n2501;
   wire FE_OFN537_n2496;
   wire FE_OFN534_n2388;
   wire FE_OFN533_n2357;
   wire FE_OFN530_n2350;
   wire FE_OFN529_n2338;
   wire FE_OFN527_n2336;
   wire FE_OFN525_n2332;
   wire FE_OFN523_n2329;
   wire FE_OFN519_n2257;
   wire FE_OFN516_n2196;
   wire FE_OFN514_n2062;
   wire FE_OFN512_n2058;
   wire FE_OFN511_n2057;
   wire FE_OFN510_n2028;
   wire FE_OFN509_n2012;
   wire FE_OFN506_n1834;
   wire FE_OFN504_n1832;
   wire FE_OFN495_n1670;
   wire FE_OFN493_n1632;
   wire FE_OFN490_n1622;
   wire FE_OFN486_n1579;
   wire FE_OFN485_n1519;
   wire FE_OFN484_n1354;
   wire FE_OFN483_n1233;
   wire FE_OFN479_n1148;
   wire FE_OFN469_n1034;
   wire FE_OFN466_n998;
   wire FE_OFN465_n945;
   wire FE_OFN461_n890;
   wire FE_OFN458_n860;
   wire FE_OFN456_n822;
   wire FE_OFN450_n808;
   wire FE_OFN429_n673;
   wire FE_OFN426_n659;
   wire FE_OFN425_n650;
   wire FE_OFN422_n641;
   wire FE_OFN419_n628;
   wire FE_OFN414_n556;
   wire FE_OFN411_n499;
   wire FE_OFN384_n118;
   wire FE_OFN383_n71;
   wire FE_OFN382_n64;
   wire FE_OFN208_n2015;
   wire FE_OFN195_HRESETn;
   wire FE_OFN194_HRESETn;
   wire FE_OFN192_HRESETn;
   wire FE_OFN190_HRESETn;
   wire FE_OFN185_HRESETn;
   wire FE_OFN184_HRESETn;
   wire FE_OFN182_HRESETn;
   wire FE_OFN181_HRESETn;
   wire FE_OFN180_HRESETn;
   wire FE_OFN179_HRESETn;
   wire FE_OFN178_HRESETn;
   wire FE_OFN177_HRESETn;
   wire FE_OFN175_HRESETn;
   wire FE_OFN174_HRESETn;
   wire FE_OFN167_HRESETn;
   wire FE_OFN166_HRESETn;
   wire FE_OFN165_HRESETn;
   wire FE_OFN164_HRESETn;
   wire FE_OFN163_HRESETn;
   wire FE_OFN159_HRESETn;
   wire FE_OFN152_HRESETn;
   wire FE_OFN145_HRESETn;
   wire FE_OFN144_HRESETn;
   wire FE_OFN139_HRESETn;
   wire FE_OFN138_HRESETn;
   wire FE_OFN135_HRESETn;
   wire FE_OFN132_n2391;
   wire FE_OFN131_n2391;
   wire FE_OFN130_n1750;
   wire FE_OFN129_n1750;
   wire FE_OFN128_n1809;
   wire FE_OFN127_n1809;
   wire FE_OFN126_n2416;
   wire FE_OFN125_n2416;
   wire FE_OFN124_n2079;
   wire FE_OFN123_n2079;
   wire FE_OFN118_HADDR_31_;
   wire FE_OFN117_HADDR_31_;
   wire FE_OFN115_HADDR_29_;
   wire FE_OFN113_HADDR_29_;
   wire FE_OFN112_HADDR_30_;
   wire FE_OFN111_HADDR_30_;
   wire FE_OFN110_HADDR_30_;
   wire FE_OFN109_n16964;
   wire FE_OFN108_n16964;
   wire FE_OFN107_n585;
   wire FE_OFN106_n585;
   wire FE_OFN105_n585;
   wire FE_OFN104_n715;
   wire FE_OFN103_n715;
   wire FE_OFN102_n715;
   wire FE_OFN100_n1086;
   wire FE_OFN99_n1086;
   wire FE_OFN98_n1104;
   wire FE_OFN95_n16864;
   wire FE_OFN93_n16864;
   wire FE_OFN91_n16864;
   wire FE_OFN90_n16849;
   wire FE_OFN89_n16849;
   wire FE_OFN88_n16849;
   wire FE_OFN87_n16848;
   wire FE_OFN86_n16848;
   wire FE_OFN85_n16839;
   wire FE_OFN84_n16839;
   wire FE_OFN83_n16839;
   wire FE_OFN82_n16856;
   wire FE_OFN81_n16856;
   wire FE_OFN80_n16856;
   wire FE_OFN79_n16834;
   wire FE_OFN78_n16834;
   wire FE_OFN77_n16834;
   wire FE_OFN75_n16806;
   wire FE_OFN73_n16806;
   wire FE_OFN72_n16867;
   wire FE_OFN70_n16867;
   wire FE_OFN68_HRESETn;
   wire FE_OFN66_HRESETn;
   wire FE_OFN65_HRESETn;
   wire FE_OFN61_HRESETn;
   wire FE_OFN60_HRESETn;
   wire FE_OFN56_HRESETn;
   wire FE_OFN52_HRESETn;
   wire FE_OFN49_HRESETn;
   wire FE_OFN48_HRESETn;
   wire FE_OFN41_HRESETn;
   wire FE_OFN40_HRESETn;
   wire FE_OFN38_HRESETn;
   wire FE_OFN33_HRESETn;
   wire FE_OFN21_n503;
   wire FE_OFN19_n1063;
   wire FE_OFN17_n16805;
   wire FE_OFN15_n16671;
   wire FE_OFN10_n1697;
   wire FE_OFN2_n2015;
   wire n8698;
   wire n8706;
   wire n9796;
   wire n9972;
   wire n10055;
   wire n10553;
   wire n11746;
   wire n11928;
   wire n11929;
   wire n11939;
   wire n11945;
   wire n11957;
   wire n11971;
   wire n13747;
   wire n13758;
   wire n13795;
   wire n13813;
   wire n13835;
   wire n13846;
   wire n13870;
   wire n13894;
   wire n13907;
   wire n13919;
   wire n13932;
   wire n13951;
   wire n13963;
   wire n13989;
   wire n14001;
   wire n14432;
   wire n14825;
   wire n14928;
   wire n14934;
   wire n14956;
   wire U811_Z_0;
   wire U810_Z_0;
   wire U809_Z_0;
   wire U806_Z_0;
   wire U805_Z_0;
   wire U804_Z_0;
   wire U803_Z_0;
   wire U802_Z_0;
   wire U801_Z_0;
   wire U800_Z_0;
   wire U799_Z_0;
   wire U798_Z_0;
   wire U797_Z_0;
   wire U795_Z_0;
   wire U792_Z_0;
   wire U791_Z_0;
   wire U790_Z_0;
   wire U789_Z_0;
   wire U788_Z_0;
   wire U787_Z_0;
   wire U786_Z_0;
   wire U785_Z_0;
   wire U784_Z_0;
   wire U783_Z_0;
   wire U782_Z_0;
   wire U781_Z_0;
   wire U780_Z_0;
   wire U779_Z_0;
   wire U778_Z_0;
   wire U777_Z_0;
   wire U776_Z_0;
   wire U775_Z_0;
   wire U774_Z_0;
   wire U773_Z_0;
   wire U772_Z_0;
   wire U771_Z_0;
   wire U770_Z_0;
   wire U769_Z_0;
   wire U768_Z_0;
   wire U767_Z_0;
   wire U766_Z_0;
   wire U765_Z_0;
   wire U764_Z_0;
   wire U763_Z_0;
   wire U762_Z_0;
   wire U761_Z_0;
   wire U760_Z_0;
   wire U756_Z_0;
   wire U755_Z_0;
   wire U754_Z_0;
   wire U752_Z_0;
   wire U751_Z_0;
   wire U750_Z_0;
   wire U749_Z_0;
   wire U748_Z_0;
   wire U747_Z_0;
   wire U746_Z_0;
   wire U745_Z_0;
   wire U744_Z_0;
   wire U743_Z_0;
   wire U742_Z_0;
   wire U741_Z_0;
   wire U740_Z_0;
   wire U739_Z_0;
   wire U738_Z_0;
   wire U737_Z_0;
   wire U736_Z_0;
   wire U735_Z_0;
   wire U734_Z_0;
   wire U733_Z_0;
   wire U732_Z_0;
   wire U731_Z_0;
   wire U730_Z_0;
   wire U729_Z_0;
   wire U728_Z_0;
   wire U727_Z_0;
   wire U726_Z_0;
   wire U725_Z_0;
   wire U724_Z_0;
   wire U723_Z_0;
   wire U722_Z_0;
   wire U721_Z_0;
   wire U720_Z_0;
   wire U719_Z_0;
   wire U718_Z_0;
   wire U717_Z_0;
   wire U716_Z_0;
   wire U715_Z_0;
   wire U714_Z_0;
   wire U713_Z_0;
   wire U712_Z_0;
   wire U711_Z_0;
   wire U710_Z_0;
   wire U709_Z_0;
   wire U708_Z_0;
   wire U707_Z_0;
   wire U706_Z_0;
   wire U705_Z_0;
   wire U704_Z_0;
   wire U703_Z_0;
   wire U702_Z_0;
   wire U701_Z_0;
   wire U700_Z_0;
   wire U699_Z_0;
   wire U698_Z_0;
   wire U697_Z_0;
   wire U696_Z_0;
   wire U695_Z_0;
   wire U694_Z_0;
   wire U693_Z_0;
   wire U692_Z_0;
   wire U691_Z_0;
   wire U687_Z_0;
   wire U686_Z_0;
   wire U685_Z_0;
   wire U684_Z_0;
   wire U683_Z_0;
   wire U682_Z_0;
   wire U681_Z_0;
   wire U680_Z_0;
   wire U679_Z_0;
   wire U678_Z_0;
   wire U677_Z_0;
   wire U676_Z_0;
   wire U675_Z_0;
   wire U674_Z_0;
   wire U673_Z_0;
   wire U672_Z_0;
   wire U671_Z_0;
   wire U670_Z_0;
   wire U669_Z_0;
   wire U668_Z_0;
   wire U667_Z_0;
   wire U666_Z_0;
   wire U665_Z_0;
   wire U664_Z_0;
   wire U663_Z_0;
   wire U662_Z_0;
   wire U661_Z_0;
   wire U660_Z_0;
   wire U659_Z_0;
   wire U658_Z_0;
   wire U657_Z_0;
   wire U656_Z_0;
   wire U655_Z_0;
   wire U654_Z_0;
   wire U653_Z_0;
   wire U652_Z_0;
   wire U651_Z_0;
   wire U650_Z_0;
   wire U649_Z_0;
   wire U648_Z_0;
   wire U647_Z_0;
   wire U646_Z_0;
   wire U645_Z_0;
   wire U644_Z_0;
   wire U643_Z_0;
   wire U642_Z_0;
   wire U641_Z_0;
   wire U640_Z_0;
   wire U639_Z_0;
   wire U638_Z_0;
   wire U637_Z_0;
   wire U636_Z_0;
   wire U635_Z_0;
   wire U634_Z_0;
   wire U633_Z_0;
   wire U632_Z_0;
   wire U631_Z_0;
   wire U630_Z_0;
   wire U629_Z_0;
   wire U628_Z_0;
   wire U627_Z_0;
   wire U626_Z_0;
   wire U625_Z_0;
   wire U624_Z_0;
   wire U623_Z_0;
   wire U622_Z_0;
   wire U621_Z_0;
   wire U620_Z_0;
   wire U619_Z_0;
   wire U618_Z_0;
   wire U617_Z_0;
   wire U614_Z_0;
   wire U613_Z_0;
   wire U612_Z_0;
   wire U611_Z_0;
   wire U610_Z_0;
   wire U609_Z_0;
   wire U608_Z_0;
   wire U607_Z_0;
   wire U606_Z_0;
   wire U605_Z_0;
   wire U604_Z_0;
   wire U603_Z_0;
   wire U602_Z_0;
   wire U601_Z_0;
   wire U600_Z_0;
   wire U599_Z_0;
   wire U598_Z_0;
   wire U597_Z_0;
   wire U596_Z_0;
   wire U595_Z_0;
   wire U594_Z_0;
   wire U593_Z_0;
   wire U592_Z_0;
   wire U591_Z_0;
   wire U590_Z_0;
   wire U589_Z_0;
   wire U588_Z_0;
   wire U587_Z_0;
   wire U586_Z_0;
   wire U585_Z_0;
   wire U584_Z_0;
   wire U583_Z_0;
   wire U582_Z_0;
   wire U581_Z_0;
   wire U580_Z_0;
   wire U579_Z_0;
   wire U578_Z_0;
   wire U577_Z_0;
   wire U576_Z_0;
   wire U575_Z_0;
   wire U574_Z_0;
   wire U573_Z_0;
   wire U572_Z_0;
   wire U571_Z_0;
   wire U570_Z_0;
   wire U569_Z_0;
   wire U568_Z_0;
   wire U567_Z_0;
   wire U566_Z_0;
   wire U565_Z_0;
   wire U564_Z_0;
   wire U563_Z_0;
   wire U562_Z_0;
   wire U561_Z_0;
   wire U560_Z_0;
   wire U559_Z_0;
   wire U558_Z_0;
   wire U557_Z_0;
   wire U556_Z_0;
   wire U555_Z_0;
   wire U554_Z_0;
   wire U553_Z_0;
   wire U552_Z_0;
   wire U551_Z_0;
   wire U550_Z_0;
   wire U549_Z_0;
   wire U548_Z_0;
   wire U547_Z_0;
   wire U546_Z_0;
   wire U545_Z_0;
   wire U544_Z_0;
   wire U543_Z_0;
   wire U542_Z_0;
   wire U541_Z_0;
   wire U540_Z_0;
   wire U539_Z_0;
   wire U538_Z_0;
   wire U537_Z_0;
   wire U536_Z_0;
   wire U535_Z_0;
   wire U534_Z_0;
   wire U533_Z_0;
   wire U532_Z_0;
   wire U531_Z_0;
   wire U530_Z_0;
   wire U529_Z_0;
   wire U528_Z_0;
   wire U527_Z_0;
   wire U526_Z_0;
   wire U525_Z_0;
   wire U524_Z_0;
   wire U523_Z_0;
   wire U522_Z_0;
   wire U521_Z_0;
   wire U520_Z_0;
   wire U519_Z_0;
   wire U518_Z_0;
   wire U517_Z_0;
   wire U516_Z_0;
   wire U515_Z_0;
   wire U514_Z_0;
   wire U513_Z_0;
   wire U512_Z_0;
   wire U511_Z_0;
   wire U510_Z_0;
   wire U509_Z_0;
   wire U508_Z_0;
   wire U507_Z_0;
   wire U506_Z_0;
   wire U505_Z_0;
   wire U504_Z_0;
   wire U503_Z_0;
   wire U502_Z_0;
   wire U501_Z_0;
   wire U500_Z_0;
   wire U499_Z_0;
   wire U498_Z_0;
   wire U497_Z_0;
   wire U496_Z_0;
   wire U495_Z_0;
   wire U494_Z_0;
   wire U493_Z_0;
   wire U492_Z_0;
   wire U491_Z_0;
   wire U490_Z_0;
   wire U489_Z_0;
   wire U488_Z_0;
   wire U487_Z_0;
   wire U486_Z_0;
   wire U483_Z_0;
   wire U482_Z_0;
   wire U481_Z_0;
   wire U480_Z_0;
   wire U479_Z_0;
   wire U478_Z_0;
   wire U477_Z_0;
   wire U476_Z_0;
   wire U475_Z_0;
   wire U474_Z_0;
   wire U473_Z_0;
   wire U472_Z_0;
   wire U471_Z_0;
   wire U470_Z_0;
   wire U469_Z_0;
   wire U468_Z_0;
   wire U467_Z_0;
   wire U466_Z_0;
   wire U465_Z_0;
   wire U464_Z_0;
   wire U463_Z_0;
   wire U462_Z_0;
   wire U461_Z_0;
   wire U460_Z_0;
   wire U459_Z_0;
   wire U458_Z_0;
   wire U457_Z_0;
   wire U456_Z_0;
   wire U455_Z_0;
   wire U454_Z_0;
   wire U453_Z_0;
   wire U452_Z_0;
   wire U449_Z_0;
   wire U448_Z_0;
   wire U447_Z_0;
   wire U446_Z_0;
   wire U445_Z_0;
   wire U444_Z_0;
   wire U443_Z_0;
   wire U442_Z_0;
   wire U441_Z_0;
   wire U440_Z_0;
   wire U439_Z_0;
   wire U438_Z_0;
   wire U437_Z_0;
   wire U436_Z_0;
   wire U435_Z_0;
   wire U434_Z_0;
   wire U433_Z_0;
   wire U432_Z_0;
   wire U431_Z_0;
   wire U430_Z_0;
   wire U429_Z_0;
   wire U428_Z_0;
   wire U427_Z_0;
   wire U426_Z_0;
   wire U425_Z_0;
   wire U424_Z_0;
   wire U423_Z_0;
   wire U422_Z_0;
   wire U421_Z_0;
   wire U420_Z_0;
   wire U419_Z_0;
   wire U418_Z_0;
   wire U415_Z_0;
   wire U414_Z_0;
   wire U413_Z_0;
   wire U412_Z_0;
   wire U411_Z_0;
   wire U410_Z_0;
   wire U409_Z_0;
   wire U408_Z_0;
   wire U407_Z_0;
   wire U406_Z_0;
   wire U405_Z_0;
   wire U404_Z_0;
   wire U403_Z_0;
   wire U402_Z_0;
   wire U401_Z_0;
   wire U400_Z_0;
   wire U399_Z_0;
   wire U398_Z_0;
   wire U397_Z_0;
   wire U396_Z_0;
   wire U395_Z_0;
   wire U394_Z_0;
   wire U393_Z_0;
   wire U392_Z_0;
   wire U391_Z_0;
   wire U390_Z_0;
   wire U389_Z_0;
   wire U388_Z_0;
   wire U387_Z_0;
   wire U386_Z_0;
   wire U385_Z_0;
   wire U384_Z_0;
   wire U383_Z_0;
   wire U382_Z_0;
   wire U381_Z_0;
   wire U380_Z_0;
   wire U379_Z_0;
   wire U378_Z_0;
   wire U377_Z_0;
   wire U376_Z_0;
   wire U375_Z_0;
   wire U374_Z_0;
   wire U373_Z_0;
   wire U372_Z_0;
   wire U371_Z_0;
   wire U370_Z_0;
   wire U369_Z_0;
   wire U368_Z_0;
   wire U367_Z_0;
   wire U366_Z_0;
   wire U365_Z_0;
   wire U364_Z_0;
   wire U363_Z_0;
   wire U362_Z_0;
   wire U361_Z_0;
   wire U360_Z_0;
   wire U359_Z_0;
   wire U358_Z_0;
   wire U357_Z_0;
   wire U356_Z_0;
   wire U355_Z_0;
   wire U354_Z_0;
   wire U353_Z_0;
   wire U352_Z_0;
   wire U349_Z_0;
   wire U348_Z_0;
   wire U347_Z_0;
   wire U346_Z_0;
   wire U345_Z_0;
   wire U344_Z_0;
   wire U343_Z_0;
   wire U342_Z_0;
   wire U341_Z_0;
   wire U340_Z_0;
   wire U339_Z_0;
   wire U338_Z_0;
   wire U337_Z_0;
   wire U336_Z_0;
   wire U335_Z_0;
   wire U334_Z_0;
   wire U333_Z_0;
   wire U332_Z_0;
   wire U331_Z_0;
   wire U330_Z_0;
   wire U329_Z_0;
   wire U328_Z_0;
   wire U327_Z_0;
   wire U326_Z_0;
   wire U325_Z_0;
   wire U324_Z_0;
   wire U323_Z_0;
   wire U322_Z_0;
   wire U321_Z_0;
   wire U320_Z_0;
   wire U319_Z_0;
   wire U318_Z_0;
   wire U317_Z_0;
   wire U315_Z_0;
   wire U314_Z_0;
   wire U313_Z_0;
   wire U312_Z_0;
   wire U311_Z_0;
   wire U310_Z_0;
   wire U309_Z_0;
   wire U308_Z_0;
   wire U307_Z_0;
   wire U306_Z_0;
   wire U305_Z_0;
   wire U304_Z_0;
   wire U303_Z_0;
   wire U302_Z_0;
   wire U301_Z_0;
   wire U300_Z_0;
   wire U299_Z_0;
   wire U298_Z_0;
   wire U297_Z_0;
   wire U296_Z_0;
   wire U295_Z_0;
   wire U294_Z_0;
   wire U293_Z_0;
   wire U292_Z_0;
   wire U291_Z_0;
   wire U290_Z_0;
   wire U289_Z_0;
   wire U288_Z_0;
   wire U287_Z_0;
   wire U286_Z_0;
   wire U285_Z_0;
   wire U284_Z_0;
   wire U283_Z_0;
   wire U282_Z_0;
   wire U281_Z_0;
   wire U280_Z_0;
   wire U279_Z_0;
   wire U278_Z_0;
   wire U277_Z_0;
   wire U276_Z_0;
   wire U275_Z_0;
   wire U274_Z_0;
   wire U273_Z_0;
   wire U272_Z_0;
   wire U271_Z_0;
   wire U270_Z_0;
   wire U269_Z_0;
   wire U268_Z_0;
   wire U265_Z_0;
   wire U264_Z_0;
   wire U263_Z_0;
   wire U262_Z_0;
   wire U261_Z_0;
   wire U260_Z_0;
   wire U259_Z_0;
   wire U258_Z_0;
   wire U257_Z_0;
   wire U256_Z_0;
   wire U255_Z_0;
   wire U254_Z_0;
   wire U253_Z_0;
   wire U252_Z_0;
   wire U251_Z_0;
   wire U250_Z_0;
   wire U247_Z_0;
   wire U246_Z_0;
   wire U245_Z_0;
   wire U244_Z_0;
   wire U243_Z_0;
   wire U242_Z_0;
   wire U241_Z_0;
   wire U240_Z_0;
   wire U239_Z_0;
   wire U238_Z_0;
   wire U237_Z_0;
   wire U236_Z_0;
   wire U235_Z_0;
   wire U234_Z_0;
   wire U233_Z_0;
   wire U232_Z_0;
   wire U229_Z_0;
   wire U227_Z_0;
   wire U189_Z_0;
   wire U186_Z_0;
   wire U180_Z_0;
   wire U175_Z_0;
   wire U163_Z_0;
   wire U158_Z_0;
   wire U144_Z_0;
   wire U134_Z_0;
   wire U122_Z_0;
   wire U121_Z_0;
   wire U105_Z_0;
   wire U98_Z_0;
   wire U97_Z_0;
   wire U4_DATA1_0;
   wire add_2073_SUM_1_;
   wire add_2073_SUM_7_;
   wire add_2073_SUM_31_;
   wire add_2073_B_1_;
   wire add_2073_A_2_;
   wire add_2073_A_3_;
   wire add_2073_A_4_;
   wire add_2073_A_5_;
   wire add_2073_A_6_;
   wire add_2073_A_7_;
   wire add_2073_A_8_;
   wire add_2073_A_9_;
   wire add_2073_A_10_;
   wire add_2073_A_11_;
   wire add_2073_A_12_;
   wire add_2073_A_13_;
   wire add_2073_A_14_;
   wire add_2073_A_15_;
   wire add_2073_A_16_;
   wire add_2073_A_17_;
   wire add_2073_A_18_;
   wire add_2073_A_19_;
   wire add_2073_A_20_;
   wire add_2073_A_21_;
   wire add_2073_A_22_;
   wire add_2073_A_23_;
   wire add_2073_A_24_;
   wire add_2073_A_25_;
   wire add_2073_A_26_;
   wire add_2073_A_27_;
   wire add_2073_A_28_;
   wire add_2073_A_29_;
   wire add_2073_A_30_;
   wire add_2073_A_31_;
   wire add_2073_A_32_;
   wire add_2082_B_1_;
   wire add_2082_B_4_;
   wire add_2082_A_1_;
   wire add_2082_A_2_;
   wire add_2082_A_3_;
   wire add_2082_A_4_;
   wire add_2082_A_5_;
   wire add_2082_A_6_;
   wire add_2082_A_7_;
   wire add_2082_A_8_;
   wire add_2082_A_9_;
   wire add_2082_A_10_;
   wire add_2082_A_11_;
   wire add_2082_A_12_;
   wire add_2082_A_13_;
   wire add_2082_A_14_;
   wire add_2082_A_15_;
   wire add_2082_A_16_;
   wire add_2082_A_17_;
   wire add_2082_A_18_;
   wire add_2082_A_19_;
   wire add_2082_A_20_;
   wire add_2082_A_21_;
   wire add_2082_A_22_;
   wire add_2082_A_23_;
   wire add_2082_A_24_;
   wire add_2082_A_25_;
   wire add_2082_A_26_;
   wire add_2082_A_27_;
   wire add_2082_A_28_;
   wire add_2082_A_29_;
   wire add_2082_A_30_;
   wire add_2082_A_31_;
   wire add_2072_SUM_1_;
   wire add_2072_SUM_2_;
   wire add_2072_SUM_3_;
   wire add_2072_SUM_4_;
   wire add_2072_SUM_5_;
   wire add_2072_SUM_6_;
   wire add_2072_SUM_7_;
   wire add_2072_SUM_8_;
   wire add_2072_SUM_9_;
   wire add_2072_SUM_10_;
   wire add_2072_SUM_11_;
   wire add_2072_SUM_12_;
   wire add_2072_SUM_13_;
   wire add_2072_SUM_14_;
   wire add_2072_SUM_15_;
   wire add_2072_SUM_16_;
   wire add_2072_SUM_17_;
   wire add_2072_SUM_18_;
   wire add_2072_SUM_19_;
   wire add_2072_SUM_20_;
   wire add_2072_SUM_21_;
   wire add_2072_SUM_22_;
   wire add_2072_SUM_23_;
   wire add_2072_SUM_24_;
   wire add_2072_SUM_25_;
   wire add_2072_SUM_26_;
   wire add_2072_SUM_27_;
   wire add_2072_SUM_28_;
   wire add_2071_SUM_1_;
   wire add_2071_SUM_2_;
   wire add_2071_SUM_3_;
   wire add_2071_SUM_4_;
   wire add_2071_SUM_5_;
   wire add_2071_SUM_6_;
   wire add_2071_SUM_7_;
   wire add_2071_SUM_8_;
   wire add_2071_SUM_9_;
   wire add_2071_SUM_10_;
   wire add_2071_SUM_11_;
   wire add_2071_SUM_12_;
   wire add_2071_SUM_13_;
   wire add_2071_SUM_14_;
   wire add_2071_SUM_15_;
   wire add_2071_SUM_16_;
   wire add_2071_SUM_17_;
   wire add_2071_SUM_18_;
   wire add_2071_SUM_19_;
   wire add_2071_SUM_20_;
   wire add_2071_SUM_21_;
   wire add_2071_SUM_22_;
   wire add_2071_SUM_23_;
   wire add_2071_SUM_24_;
   wire add_2071_SUM_25_;
   wire add_2071_SUM_26_;
   wire add_2071_SUM_27_;
   wire add_2071_SUM_28_;
   wire add_2071_SUM_29_;
   wire sub_2069_carry_2_;
   wire sub_2069_carry_3_;
   wire sub_2069_carry_4_;
   wire sub_2069_carry_5_;
   wire sub_2069_carry_6_;
   wire sub_2069_carry_7_;
   wire sub_2069_carry_8_;
   wire sub_2069_SUM_1_;
   wire sub_2069_SUM_2_;
   wire sub_2069_SUM_3_;
   wire sub_2069_SUM_4_;
   wire sub_2069_SUM_5_;
   wire sub_2069_SUM_6_;
   wire sub_2069_SUM_7_;
   wire sub_2069_SUM_8_;
   wire sub_2069_A_1_;
   wire sub_2069_A_2_;
   wire sub_2069_A_3_;
   wire sub_2069_A_4_;
   wire sub_2069_A_5_;
   wire sub_2069_A_6_;
   wire sub_2069_A_7_;
   wire sub_2069_A_8_;
   wire sub_2068_carry_2_;
   wire sub_2068_carry_3_;
   wire sub_2068_carry_4_;
   wire sub_2068_carry_5_;
   wire sub_2068_carry_6_;
   wire sub_2068_carry_7_;
   wire sub_2068_carry_8_;
   wire sub_2068_carry_9_;
   wire sub_2068_carry_10_;
   wire sub_2068_carry_11_;
   wire sub_2068_carry_12_;
   wire sub_2068_carry_13_;
   wire sub_2068_carry_14_;
   wire sub_2068_carry_15_;
   wire sub_2068_carry_16_;
   wire sub_2068_carry_17_;
   wire sub_2068_carry_18_;
   wire sub_2068_carry_19_;
   wire sub_2068_carry_20_;
   wire sub_2068_carry_21_;
   wire sub_2068_carry_22_;
   wire sub_2068_carry_23_;
   wire sub_2068_SUM_1_;
   wire sub_2068_SUM_2_;
   wire sub_2068_SUM_3_;
   wire sub_2068_SUM_4_;
   wire sub_2068_SUM_5_;
   wire sub_2068_SUM_6_;
   wire sub_2068_SUM_7_;
   wire sub_2068_SUM_8_;
   wire sub_2068_SUM_9_;
   wire sub_2068_SUM_10_;
   wire sub_2068_SUM_11_;
   wire sub_2068_SUM_12_;
   wire sub_2068_SUM_13_;
   wire sub_2068_SUM_14_;
   wire sub_2068_SUM_15_;
   wire sub_2068_SUM_16_;
   wire sub_2068_SUM_17_;
   wire sub_2068_SUM_18_;
   wire sub_2068_SUM_19_;
   wire sub_2068_SUM_20_;
   wire sub_2068_SUM_21_;
   wire sub_2068_SUM_22_;
   wire sub_2068_A_0_;
   wire sub_2068_A_1_;
   wire sub_2068_A_2_;
   wire sub_2068_A_3_;
   wire sub_2068_A_4_;
   wire sub_2068_A_5_;
   wire sub_2068_A_6_;
   wire sub_2068_A_7_;
   wire sub_2068_A_8_;
   wire sub_2068_A_9_;
   wire sub_2068_A_10_;
   wire sub_2068_A_11_;
   wire sub_2068_A_12_;
   wire sub_2068_A_13_;
   wire sub_2068_A_14_;
   wire sub_2068_A_15_;
   wire sub_2068_A_16_;
   wire sub_2068_A_17_;
   wire sub_2068_A_18_;
   wire sub_2068_A_19_;
   wire sub_2068_A_20_;
   wire sub_2068_A_21_;
   wire sub_2068_A_22_;
   wire sub_2068_A_23_;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n33;
   wire n36;
   wire n37;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n44;
   wire n45;
   wire n46;
   wire n48;
   wire n49;
   wire n50;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n76;
   wire n77;
   wire n78;
   wire n80;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n104;
   wire n105;
   wire n106;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n113;
   wire n114;
   wire n115;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n122;
   wire n123;
   wire n124;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n131;
   wire n132;
   wire n133;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n140;
   wire n141;
   wire n142;
   wire n144;
   wire n145;
   wire n146;
   wire n148;
   wire n149;
   wire n150;
   wire n152;
   wire n153;
   wire n154;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n175;
   wire n176;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n264;
   wire n265;
   wire n266;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n320;
   wire n322;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n329;
   wire n330;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n440;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n471;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n510;
   wire n511;
   wire n512;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n522;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n788;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n863;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n994;
   wire n995;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1750;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2209;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2271;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2297;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2402;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2433;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2452;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2481;
   wire n2484;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2507;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2531;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2562;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2585;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2612;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2635;
   wire n2636;
   wire n2637;
   wire n2639;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2700;
   wire n2701;
   wire n2702;
   wire n2703;
   wire n2705;
   wire n2713;
   wire n2714;
   wire n2715;
   wire n2716;
   wire n2717;
   wire n2718;
   wire n2719;
   wire n2720;
   wire n2721;
   wire n2722;
   wire n2723;
   wire n2724;
   wire n2725;
   wire n2726;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2731;
   wire n2732;
   wire n2733;
   wire n2734;
   wire n2735;
   wire n2736;
   wire n2738;
   wire n2746;
   wire n2747;
   wire n2748;
   wire n2749;
   wire n2750;
   wire n2751;
   wire n2752;
   wire n2753;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2764;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2775;
   wire n2776;
   wire n2777;
   wire n2778;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2787;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2809;
   wire n2817;
   wire n2818;
   wire n2819;
   wire n2820;
   wire n2821;
   wire n2822;
   wire n2823;
   wire n2824;
   wire n2825;
   wire n2826;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2830;
   wire n2831;
   wire n2833;
   wire n2841;
   wire n2842;
   wire n2843;
   wire n2844;
   wire n2845;
   wire n2846;
   wire n2847;
   wire n2848;
   wire n2849;
   wire n2850;
   wire n2851;
   wire n2852;
   wire n2853;
   wire n2854;
   wire n2856;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2961;
   wire n2964;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3022;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3041;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3059;
   wire n3060;
   wire n3061;
   wire n3062;
   wire n3063;
   wire n3064;
   wire n3065;
   wire n3066;
   wire n3067;
   wire n3068;
   wire n3069;
   wire n3070;
   wire n3071;
   wire n3072;
   wire n3073;
   wire n3074;
   wire n3075;
   wire n3076;
   wire n3077;
   wire n3078;
   wire n3079;
   wire n3080;
   wire n3081;
   wire n3082;
   wire n3083;
   wire n3084;
   wire n3085;
   wire n3086;
   wire n3087;
   wire n3088;
   wire n3089;
   wire n3090;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3134;
   wire n3142;
   wire n3143;
   wire n3144;
   wire n3145;
   wire n3146;
   wire n3147;
   wire n3148;
   wire n3149;
   wire n3150;
   wire n3151;
   wire n3152;
   wire n3153;
   wire n3155;
   wire n3163;
   wire n3164;
   wire n3165;
   wire n3166;
   wire n3167;
   wire n3168;
   wire n3169;
   wire n3170;
   wire n3171;
   wire n3172;
   wire n3173;
   wire n3174;
   wire n3175;
   wire n3177;
   wire n3178;
   wire n3179;
   wire n3180;
   wire n3181;
   wire n3182;
   wire n3183;
   wire n3184;
   wire n3185;
   wire n3186;
   wire n3187;
   wire n3188;
   wire n3189;
   wire n3190;
   wire n3191;
   wire n3192;
   wire n3193;
   wire n3194;
   wire n3195;
   wire n3196;
   wire n3197;
   wire n3199;
   wire n3207;
   wire n3208;
   wire n3209;
   wire n3210;
   wire n3211;
   wire n3212;
   wire n3213;
   wire n3214;
   wire n3215;
   wire n3217;
   wire n3218;
   wire n3219;
   wire n3220;
   wire n3221;
   wire n3222;
   wire n3223;
   wire n3224;
   wire n3225;
   wire n3226;
   wire n3227;
   wire n3228;
   wire n3229;
   wire n3230;
   wire n3231;
   wire n3233;
   wire n3234;
   wire n3237;
   wire n3238;
   wire n3239;
   wire n3240;
   wire n3241;
   wire n3242;
   wire n3243;
   wire n3244;
   wire n3245;
   wire n3246;
   wire n3247;
   wire n3248;
   wire n3249;
   wire n3250;
   wire n3251;
   wire n3252;
   wire n3253;
   wire n3254;
   wire n3255;
   wire n3256;
   wire n3257;
   wire n3258;
   wire n3259;
   wire n3260;
   wire n3261;
   wire n3262;
   wire n3263;
   wire n3264;
   wire n3265;
   wire n3266;
   wire n3267;
   wire n3268;
   wire n3269;
   wire n3270;
   wire n3271;
   wire n3272;
   wire n3273;
   wire n3274;
   wire n3275;
   wire n3276;
   wire n3277;
   wire n3278;
   wire n3279;
   wire n3280;
   wire n3281;
   wire n3282;
   wire n3283;
   wire n3284;
   wire n3285;
   wire n3286;
   wire n3287;
   wire n3288;
   wire n3289;
   wire n3290;
   wire n3291;
   wire n3292;
   wire n3293;
   wire n3294;
   wire n3295;
   wire n3296;
   wire n3305;
   wire n3306;
   wire n3307;
   wire n3308;
   wire n3309;
   wire n3310;
   wire n3311;
   wire n3312;
   wire n3313;
   wire n3314;
   wire n3315;
   wire n3316;
   wire n3317;
   wire n3318;
   wire n3319;
   wire n3320;
   wire n3321;
   wire n3322;
   wire n3323;
   wire n3324;
   wire n3325;
   wire n3326;
   wire n3327;
   wire n3328;
   wire n3329;
   wire n3330;
   wire n3331;
   wire n3332;
   wire n3333;
   wire n3334;
   wire n3335;
   wire n3336;
   wire n3337;
   wire n3338;
   wire n3339;
   wire n3340;
   wire n3341;
   wire n3342;
   wire n3343;
   wire n3344;
   wire n3345;
   wire n3346;
   wire n3347;
   wire n3348;
   wire n3349;
   wire n3350;
   wire n3351;
   wire n3352;
   wire n3353;
   wire n3354;
   wire n3355;
   wire n3356;
   wire n3357;
   wire n3358;
   wire n3359;
   wire n3360;
   wire n3361;
   wire n3362;
   wire n3363;
   wire n3364;
   wire n3365;
   wire n3366;
   wire n3367;
   wire n3376;
   wire n3377;
   wire n3378;
   wire n3379;
   wire n3380;
   wire n3381;
   wire n3382;
   wire n3383;
   wire n3384;
   wire n3385;
   wire n3386;
   wire n3387;
   wire n3388;
   wire n3389;
   wire n3390;
   wire n3391;
   wire n3392;
   wire n3393;
   wire n3394;
   wire n3395;
   wire n3396;
   wire n3397;
   wire n3398;
   wire n3399;
   wire n3400;
   wire n3401;
   wire n3402;
   wire n3403;
   wire n3404;
   wire n3405;
   wire n3406;
   wire n3407;
   wire n3408;
   wire n3409;
   wire n3410;
   wire n3411;
   wire n3420;
   wire n3421;
   wire n3422;
   wire n3423;
   wire n3424;
   wire n3425;
   wire n3426;
   wire n3427;
   wire n3428;
   wire n3429;
   wire n3430;
   wire n3431;
   wire n3432;
   wire n3433;
   wire n3434;
   wire n3435;
   wire n3436;
   wire n3437;
   wire n3438;
   wire n3439;
   wire n3440;
   wire n3441;
   wire n3442;
   wire n3443;
   wire n3444;
   wire n3445;
   wire n3446;
   wire n3447;
   wire n3448;
   wire n3449;
   wire n3450;
   wire n3451;
   wire n3452;
   wire n3453;
   wire n3454;
   wire n3455;
   wire n3456;
   wire n3457;
   wire n3458;
   wire n3467;
   wire n3468;
   wire n3469;
   wire n3470;
   wire n3471;
   wire n3472;
   wire n3473;
   wire n3474;
   wire n3475;
   wire n3476;
   wire n3477;
   wire n3478;
   wire n3479;
   wire n3480;
   wire n3481;
   wire n3482;
   wire n3483;
   wire n3484;
   wire n3485;
   wire n3486;
   wire n3487;
   wire n3488;
   wire n3489;
   wire n3490;
   wire n3491;
   wire n3492;
   wire n3493;
   wire n3494;
   wire n3495;
   wire n3496;
   wire n3497;
   wire n3498;
   wire n3499;
   wire n3500;
   wire n3501;
   wire n3502;
   wire n3503;
   wire n3504;
   wire n3505;
   wire n3506;
   wire n3507;
   wire n3508;
   wire n3509;
   wire n3510;
   wire n3511;
   wire n3512;
   wire n3513;
   wire n3514;
   wire n3515;
   wire n3516;
   wire n3517;
   wire n3518;
   wire n3519;
   wire n3520;
   wire n3521;
   wire n3522;
   wire n3523;
   wire n3524;
   wire n3525;
   wire n3526;
   wire n3527;
   wire n3528;
   wire n3529;
   wire n3530;
   wire n3531;
   wire n3532;
   wire n3533;
   wire n3534;
   wire n3535;
   wire n3536;
   wire n3537;
   wire n3538;
   wire n3539;
   wire n3540;
   wire n3541;
   wire n3542;
   wire n3543;
   wire n3544;
   wire n3545;
   wire n3546;
   wire n3547;
   wire n3548;
   wire n3549;
   wire n3550;
   wire n3551;
   wire n3552;
   wire n3553;
   wire n3554;
   wire n3555;
   wire n3556;
   wire n3557;
   wire n3558;
   wire n3559;
   wire n3560;
   wire n3561;
   wire n3562;
   wire n3563;
   wire n3564;
   wire n3565;
   wire n3566;
   wire n3567;
   wire n3568;
   wire n3569;
   wire n3570;
   wire n3571;
   wire n3572;
   wire n3573;
   wire n3574;
   wire n3575;
   wire n3576;
   wire n3577;
   wire n3578;
   wire n3579;
   wire n3580;
   wire n3581;
   wire n3582;
   wire n3583;
   wire n3584;
   wire n3585;
   wire n3586;
   wire n3587;
   wire n3588;
   wire n3592;
   wire n3593;
   wire n3597;
   wire n3598;
   wire n3601;
   wire n3602;
   wire n3603;
   wire n3604;
   wire n3605;
   wire n3606;
   wire n3607;
   wire n3608;
   wire n3609;
   wire n3610;
   wire n3611;
   wire n3612;
   wire n3613;
   wire n3614;
   wire n3615;
   wire n3616;
   wire n3617;
   wire n3618;
   wire n3620;
   wire n3621;
   wire n3622;
   wire n3623;
   wire n3624;
   wire n3625;
   wire n3626;
   wire n3627;
   wire n3628;
   wire n3629;
   wire n3634;
   wire n3645;
   wire n3646;
   wire n3647;
   wire n3650;
   wire n3655;
   wire n3656;
   wire n3657;
   wire n3660;
   wire n3665;
   wire n3666;
   wire n3667;
   wire n3670;
   wire n3675;
   wire n3676;
   wire n3677;
   wire n3678;
   wire n3681;
   wire n3686;
   wire n3687;
   wire n3688;
   wire n3691;
   wire n3696;
   wire n3697;
   wire n3698;
   wire n3701;
   wire n3706;
   wire n3707;
   wire n3708;
   wire n3711;
   wire n3716;
   wire n3717;
   wire n3718;
   wire n3719;
   wire n3720;
   wire n3721;
   wire n3722;
   wire n3723;
   wire n3724;
   wire n3725;
   wire n3726;
   wire n3727;
   wire n3728;
   wire n3729;
   wire n3730;
   wire n3731;
   wire n3732;
   wire n3733;
   wire n3734;
   wire n3735;
   wire n3736;
   wire n3737;
   wire n3738;
   wire n3739;
   wire n3740;
   wire n3741;
   wire n3742;
   wire n3743;
   wire n3744;
   wire n3745;
   wire n3746;
   wire n3747;
   wire n3748;
   wire n3749;
   wire n3750;
   wire n3751;
   wire n3752;
   wire n3753;
   wire n3754;
   wire n3755;
   wire n3756;
   wire n3757;
   wire n3758;
   wire n3759;
   wire n3760;
   wire n3761;
   wire n3762;
   wire n3763;
   wire n3764;
   wire n3765;
   wire n3766;
   wire n3767;
   wire n3768;
   wire n3769;
   wire n3770;
   wire n3771;
   wire n3772;
   wire n3774;
   wire n3775;
   wire n3776;
   wire n3777;
   wire n3778;
   wire n3779;
   wire n3780;
   wire n3781;
   wire n3782;
   wire n3783;
   wire n3784;
   wire n3785;
   wire n3786;
   wire n3787;
   wire n3788;
   wire n3789;
   wire n3790;
   wire n3791;
   wire n3792;
   wire n3793;
   wire n3794;
   wire n3795;
   wire n3796;
   wire n3797;
   wire n3798;
   wire n3799;
   wire n3800;
   wire n3801;
   wire n3802;
   wire n3803;
   wire n3804;
   wire n3805;
   wire n3806;
   wire n3807;
   wire n3808;
   wire n3809;
   wire n3810;
   wire n3811;
   wire n3812;
   wire n3813;
   wire n3814;
   wire n3815;
   wire n3816;
   wire n3817;
   wire n3818;
   wire n3819;
   wire n3820;
   wire n3821;
   wire n3822;
   wire n3823;
   wire n3824;
   wire n3825;
   wire n3826;
   wire n3827;
   wire n3828;
   wire n3829;
   wire n3830;
   wire n3831;
   wire n3832;
   wire n3833;
   wire n3834;
   wire n3835;
   wire n3836;
   wire n3837;
   wire n3838;
   wire n3839;
   wire n3840;
   wire n3841;
   wire n3842;
   wire n3843;
   wire n3844;
   wire n3845;
   wire n3846;
   wire n3847;
   wire n3848;
   wire n3849;
   wire n3850;
   wire n3851;
   wire n3852;
   wire n3853;
   wire n3854;
   wire n3855;
   wire n3856;
   wire n3857;
   wire n3858;
   wire n3859;
   wire n3860;
   wire n3861;
   wire n3862;
   wire n3863;
   wire n3864;
   wire n3865;
   wire n3866;
   wire n3867;
   wire n3868;
   wire n3869;
   wire n3870;
   wire n3871;
   wire n3872;
   wire n3873;
   wire n3874;
   wire n3875;
   wire n3876;
   wire n3877;
   wire n3878;
   wire n3879;
   wire n3880;
   wire n3883;
   wire n3888;
   wire n3889;
   wire n3890;
   wire n3893;
   wire n3898;
   wire n3899;
   wire n3900;
   wire n3903;
   wire n3908;
   wire n3909;
   wire n3910;
   wire n3913;
   wire n3918;
   wire n3919;
   wire n3920;
   wire n3921;
   wire n3924;
   wire n3929;
   wire n3930;
   wire n3931;
   wire n3934;
   wire n3939;
   wire n3940;
   wire n3941;
   wire n3944;
   wire n3949;
   wire n3950;
   wire n3951;
   wire n3954;
   wire n3959;
   wire n3960;
   wire n3961;
   wire n3962;
   wire n3963;
   wire n3964;
   wire n3965;
   wire n3966;
   wire n3967;
   wire n3968;
   wire n3969;
   wire n3970;
   wire n3971;
   wire n3972;
   wire n3973;
   wire n3974;
   wire n3977;
   wire n3982;
   wire n3983;
   wire n3984;
   wire n3987;
   wire n3992;
   wire n3993;
   wire n3994;
   wire n3997;
   wire n4002;
   wire n4003;
   wire n4004;
   wire n4007;
   wire n4012;
   wire n4013;
   wire n4014;
   wire n4015;
   wire n4018;
   wire n4023;
   wire n4024;
   wire n4025;
   wire n4028;
   wire n4033;
   wire n4034;
   wire n4035;
   wire n4038;
   wire n4043;
   wire n4044;
   wire n4045;
   wire n4046;
   wire n4049;
   wire n4054;
   wire n4055;
   wire n4056;
   wire n4057;
   wire n4058;
   wire n4059;
   wire n4060;
   wire n4061;
   wire n4062;
   wire n4063;
   wire n4064;
   wire n4065;
   wire n4066;
   wire n4067;
   wire n4068;
   wire n4069;
   wire n4070;
   wire n4071;
   wire n4072;
   wire n4073;
   wire n4074;
   wire n4075;
   wire n4076;
   wire n4077;
   wire n4078;
   wire n4079;
   wire n4080;
   wire n4081;
   wire n4084;
   wire n4089;
   wire n4090;
   wire n4091;
   wire n4094;
   wire n4099;
   wire n4100;
   wire n4101;
   wire n4104;
   wire n4109;
   wire n4110;
   wire n4111;
   wire n4114;
   wire n4119;
   wire n4120;
   wire n4121;
   wire n4122;
   wire n4125;
   wire n4130;
   wire n4131;
   wire n4132;
   wire n4133;
   wire n4134;
   wire n4137;
   wire n4142;
   wire n4143;
   wire n4144;
   wire n4145;
   wire n4148;
   wire n4153;
   wire n4154;
   wire n4155;
   wire n4156;
   wire n4157;
   wire n4158;
   wire n4161;
   wire n4162;
   wire n4163;
   wire n4168;
   wire n4169;
   wire n4170;
   wire n4171;
   wire n4172;
   wire n4173;
   wire n4174;
   wire n4175;
   wire n4176;
   wire n4177;
   wire n4178;
   wire n4179;
   wire n4180;
   wire n4181;
   wire n4182;
   wire n4183;
   wire n4184;
   wire n4185;
   wire n4186;
   wire n4187;
   wire n4188;
   wire n4189;
   wire n4190;
   wire n4191;
   wire n4192;
   wire n4193;
   wire n4194;
   wire n4195;
   wire n4196;
   wire n4197;
   wire n4198;
   wire n4199;
   wire n4200;
   wire n4201;
   wire n4202;
   wire n4203;
   wire n4204;
   wire n4205;
   wire n4206;
   wire n4207;
   wire n4210;
   wire n4211;
   wire n4216;
   wire n4221;
   wire n4224;
   wire n4227;
   wire n4230;
   wire n4231;
   wire n4232;
   wire n4233;
   wire n4234;
   wire n4235;
   wire n4236;
   wire n4238;
   wire n4239;
   wire n4240;
   wire n4241;
   wire n4242;
   wire n4243;
   wire n4244;
   wire n4245;
   wire n4246;
   wire n4247;
   wire n4248;
   wire n4250;
   wire n4251;
   wire n4252;
   wire n4253;
   wire n4254;
   wire n4255;
   wire n4256;
   wire n4257;
   wire n4259;
   wire n4260;
   wire n4261;
   wire n4262;
   wire n4263;
   wire n4264;
   wire n4265;
   wire n4266;
   wire n4267;
   wire n4268;
   wire n4270;
   wire n4271;
   wire n4272;
   wire n4273;
   wire n4274;
   wire n4275;
   wire n4276;
   wire n4277;
   wire n4278;
   wire n4279;
   wire n4281;
   wire n4282;
   wire n4283;
   wire n4284;
   wire n4285;
   wire n4286;
   wire n4287;
   wire n4288;
   wire n4290;
   wire n4291;
   wire n4292;
   wire n4293;
   wire n4294;
   wire n4295;
   wire n4296;
   wire n4297;
   wire n4299;
   wire n4300;
   wire n4301;
   wire n4302;
   wire n4303;
   wire n4304;
   wire n4305;
   wire n4306;
   wire n4307;
   wire n4308;
   wire n4309;
   wire n4310;
   wire n4311;
   wire n4312;
   wire n4313;
   wire n4314;
   wire n4315;
   wire n4316;
   wire n4317;
   wire n4318;
   wire n4319;
   wire n4320;
   wire n4321;
   wire n4322;
   wire n4323;
   wire n4324;
   wire n4325;
   wire n4326;
   wire n4327;
   wire n4328;
   wire n4329;
   wire n4330;
   wire n4331;
   wire n4332;
   wire n4333;
   wire n4334;
   wire n4335;
   wire n4336;
   wire n4337;
   wire n4338;
   wire n4339;
   wire n4340;
   wire n4341;
   wire n4342;
   wire n4343;
   wire n4344;
   wire n4345;
   wire n4346;
   wire n4347;
   wire n4348;
   wire n4349;
   wire n4350;
   wire n4351;
   wire n4352;
   wire n4353;
   wire n4354;
   wire n4355;
   wire n4356;
   wire n4357;
   wire n4358;
   wire n4359;
   wire n4360;
   wire n4361;
   wire n4362;
   wire n4363;
   wire n4364;
   wire n4365;
   wire n4366;
   wire n4367;
   wire n4368;
   wire n4369;
   wire n4370;
   wire n4371;
   wire n4372;
   wire n4373;
   wire n4374;
   wire n4375;
   wire n4376;
   wire n4377;
   wire n4378;
   wire n4379;
   wire n4380;
   wire n4381;
   wire n4382;
   wire n4383;
   wire n4384;
   wire n4385;
   wire n4386;
   wire n4387;
   wire n4388;
   wire n4389;
   wire n4390;
   wire n4391;
   wire n4392;
   wire n4393;
   wire n4394;
   wire n4395;
   wire n4396;
   wire n4397;
   wire n4398;
   wire n4399;
   wire n4400;
   wire n4401;
   wire n4402;
   wire n4403;
   wire n4404;
   wire n4405;
   wire n4406;
   wire n4407;
   wire n4408;
   wire n4410;
   wire n4411;
   wire n4412;
   wire n4413;
   wire n4414;
   wire n4420;
   wire n4421;
   wire n4422;
   wire n4426;
   wire n4427;
   wire n4428;
   wire n4429;
   wire n4430;
   wire n4431;
   wire n4432;
   wire n4433;
   wire n4434;
   wire n4435;
   wire n4436;
   wire n4437;
   wire n4438;
   wire n4439;
   wire n4440;
   wire n4441;
   wire n4442;
   wire n4443;
   wire n4445;
   wire n4446;
   wire n4447;
   wire n4448;
   wire n4449;
   wire n4450;
   wire n4451;
   wire n4452;
   wire n4453;
   wire n4454;
   wire n4456;
   wire n4457;
   wire n4458;
   wire n4459;
   wire n4460;
   wire n4461;
   wire n4462;
   wire n4463;
   wire n4464;
   wire n4466;
   wire n4467;
   wire n4468;
   wire n4469;
   wire n4472;
   wire n4474;
   wire n4475;
   wire n4476;
   wire n4479;
   wire n4480;
   wire n4481;
   wire n4482;
   wire n4484;
   wire n4486;
   wire n4487;
   wire n4488;
   wire n4491;
   wire n4492;
   wire n4493;
   wire n4494;
   wire n4495;
   wire n4496;
   wire n4497;
   wire n4498;
   wire n4500;
   wire n4501;
   wire n4502;
   wire n4503;
   wire n4504;
   wire n4505;
   wire n4506;
   wire n4507;
   wire n4509;
   wire n4510;
   wire n4511;
   wire n4512;
   wire n4513;
   wire n4514;
   wire n4515;
   wire n4516;
   wire n4519;
   wire n4520;
   wire n4521;
   wire n4522;
   wire n4523;
   wire n4524;
   wire n4525;
   wire n4526;
   wire n4528;
   wire n4529;
   wire n4530;
   wire n4531;
   wire n4532;
   wire n4533;
   wire n4534;
   wire n4535;
   wire n4538;
   wire n4539;
   wire n4540;
   wire n4541;
   wire n4542;
   wire n4543;
   wire n4544;
   wire n4545;
   wire n4547;
   wire n4548;
   wire n4549;
   wire n4550;
   wire n4551;
   wire n4552;
   wire n4553;
   wire n4554;
   wire n4557;
   wire n4558;
   wire n4559;
   wire n4560;
   wire n4561;
   wire n4562;
   wire n4563;
   wire n4564;
   wire n4566;
   wire n4567;
   wire n4568;
   wire n4569;
   wire n4570;
   wire n4571;
   wire n4572;
   wire n4573;
   wire n4574;
   wire n4577;
   wire n4578;
   wire n4579;
   wire n4580;
   wire n4581;
   wire n4582;
   wire n4583;
   wire n4584;
   wire n4587;
   wire n4588;
   wire n4589;
   wire n4590;
   wire n4591;
   wire n4592;
   wire n4593;
   wire n4594;
   wire n4595;
   wire n4596;
   wire n4597;
   wire n4599;
   wire n4600;
   wire n4601;
   wire n4602;
   wire n4603;
   wire n4604;
   wire n4605;
   wire n4606;
   wire n4607;
   wire n4609;
   wire n4610;
   wire n4611;
   wire n4612;
   wire n4613;
   wire n4614;
   wire n4615;
   wire n4616;
   wire n4617;
   wire n4619;
   wire n4620;
   wire n4621;
   wire n4622;
   wire n4623;
   wire n4624;
   wire n4625;
   wire n4626;
   wire n4627;
   wire n4629;
   wire n4630;
   wire n4631;
   wire n4632;
   wire n4633;
   wire n4634;
   wire n4635;
   wire n4636;
   wire n4637;
   wire n4639;
   wire n4640;
   wire n4641;
   wire n4642;
   wire n4643;
   wire n4644;
   wire n4645;
   wire n4646;
   wire n4647;
   wire n4649;
   wire n4650;
   wire n4651;
   wire n4652;
   wire n4653;
   wire n4654;
   wire n4655;
   wire n4656;
   wire n4657;
   wire n4658;
   wire n4659;
   wire n4660;
   wire n4661;
   wire n4662;
   wire n4663;
   wire n4664;
   wire n4665;
   wire n4666;
   wire n4668;
   wire n4669;
   wire n4670;
   wire n4671;
   wire n4672;
   wire n4673;
   wire n4674;
   wire n4675;
   wire n4676;
   wire n4677;
   wire n4678;
   wire n4679;
   wire n4680;
   wire n4681;
   wire n4682;
   wire n4683;
   wire n4684;
   wire n4685;
   wire n4686;
   wire n4687;
   wire n4688;
   wire n4689;
   wire n4690;
   wire n4691;
   wire n4692;
   wire n4693;
   wire n4694;
   wire n4695;
   wire n4696;
   wire n4697;
   wire n4698;
   wire n4699;
   wire n4700;
   wire n4701;
   wire n4702;
   wire n4703;
   wire n4704;
   wire n4705;
   wire n4706;
   wire n4707;
   wire n4708;
   wire n4709;
   wire n4710;
   wire n4711;
   wire n4712;
   wire n4713;
   wire n4714;
   wire n4715;
   wire n4716;
   wire n4717;
   wire n4718;
   wire n4719;
   wire n4720;
   wire n4721;
   wire n4722;
   wire n4723;
   wire n4724;
   wire n4725;
   wire n4726;
   wire n4727;
   wire n4728;
   wire n4729;
   wire n4730;
   wire n4731;
   wire n4732;
   wire n4733;
   wire n4734;
   wire n4735;
   wire n4736;
   wire n4737;
   wire n4738;
   wire n4739;
   wire n4740;
   wire n4741;
   wire n4742;
   wire n4743;
   wire n4744;
   wire n4745;
   wire n4746;
   wire n4747;
   wire n4748;
   wire n4749;
   wire n4750;
   wire n4751;
   wire n4752;
   wire n4753;
   wire n4755;
   wire n4761;
   wire n4762;
   wire n4763;
   wire n4764;
   wire n4765;
   wire n4766;
   wire n4767;
   wire n4768;
   wire n4769;
   wire n4770;
   wire n4771;
   wire n4772;
   wire n4773;
   wire n4774;
   wire n4777;
   wire n4778;
   wire n4779;
   wire n4780;
   wire n4781;
   wire n4782;
   wire n4783;
   wire n4784;
   wire n4785;
   wire n4786;
   wire n4787;
   wire n4788;
   wire n4789;
   wire n4790;
   wire n4791;
   wire n4792;
   wire n4795;
   wire n4796;
   wire n4797;
   wire n4798;
   wire n4799;
   wire n4800;
   wire n4801;
   wire n4802;
   wire n4804;
   wire n4806;
   wire n4811;
   wire n4812;
   wire n4813;
   wire n4814;
   wire n4815;
   wire n4816;
   wire n4817;
   wire n4819;
   wire n4820;
   wire n4821;
   wire n4822;
   wire n4824;
   wire n4825;
   wire n4826;
   wire n4827;
   wire n4828;
   wire n4829;
   wire n4830;
   wire n4831;
   wire n4832;
   wire n4833;
   wire n4834;
   wire n4843;
   wire n4845;
   wire n4846;
   wire n4847;
   wire n4848;
   wire n4850;
   wire n4851;
   wire n4852;
   wire n4853;
   wire n4854;
   wire n4855;
   wire n4856;
   wire n4857;
   wire n4858;
   wire n4859;
   wire n4860;
   wire n4861;
   wire n4862;
   wire n4863;
   wire n4864;
   wire n4865;
   wire n4866;
   wire n4867;
   wire n4868;
   wire n4869;
   wire n4870;
   wire n4871;
   wire n4872;
   wire n4873;
   wire n4874;
   wire n4875;
   wire n4876;
   wire n4878;
   wire n4879;
   wire n4880;
   wire n4881;
   wire n4882;
   wire n4883;
   wire n4884;
   wire n4885;
   wire n4886;
   wire n4887;
   wire n4888;
   wire n4889;
   wire n4890;
   wire n4891;
   wire n4892;
   wire n4893;
   wire n4894;
   wire n4895;
   wire n4896;
   wire n4897;
   wire n4898;
   wire n4899;
   wire n4900;
   wire n4901;
   wire n4902;
   wire n4903;
   wire n4904;
   wire n4905;
   wire n4906;
   wire n4907;
   wire n4908;
   wire n4909;
   wire n4910;
   wire n4911;
   wire n4912;
   wire n4913;
   wire n4914;
   wire n4915;
   wire n4916;
   wire n4917;
   wire n4918;
   wire n4919;
   wire n4920;
   wire n4921;
   wire n4922;
   wire n4923;
   wire n4924;
   wire n4925;
   wire n4926;
   wire n4927;
   wire n4928;
   wire n4929;
   wire n4930;
   wire n4931;
   wire n4932;
   wire n4933;
   wire n4934;
   wire n4935;
   wire n4936;
   wire n4937;
   wire n4938;
   wire n4939;
   wire n4940;
   wire n4941;
   wire n4942;
   wire n4943;
   wire n4944;
   wire n4945;
   wire n4947;
   wire n4948;
   wire n4949;
   wire n4950;
   wire n4951;
   wire n4952;
   wire n4953;
   wire n4954;
   wire n4955;
   wire n4956;
   wire n4959;
   wire n4960;
   wire n4961;
   wire n4962;
   wire n4963;
   wire n4964;
   wire n4965;
   wire n4966;
   wire n4967;
   wire n4968;
   wire n4969;
   wire n4970;
   wire n4971;
   wire n4972;
   wire n4973;
   wire n4974;
   wire n4978;
   wire n4979;
   wire n4980;
   wire n4981;
   wire n4982;
   wire n4983;
   wire n4984;
   wire n4985;
   wire n4986;
   wire n4987;
   wire n4988;
   wire n4989;
   wire n4990;
   wire n4991;
   wire n4992;
   wire n4993;
   wire n4994;
   wire n4995;
   wire n4996;
   wire n4997;
   wire n4998;
   wire n5003;
   wire n5004;
   wire n5005;
   wire n5006;
   wire n5007;
   wire n5008;
   wire n5009;
   wire n5010;
   wire n5011;
   wire n5012;
   wire n5013;
   wire n5014;
   wire n5015;
   wire n5016;
   wire n5017;
   wire n5018;
   wire n5019;
   wire n5020;
   wire n5021;
   wire n5022;
   wire n5023;
   wire n5024;
   wire n5025;
   wire n5026;
   wire n5027;
   wire n5028;
   wire n5029;
   wire n5030;
   wire n5031;
   wire n5032;
   wire n5033;
   wire n5034;
   wire n5036;
   wire n5037;
   wire n5038;
   wire n5039;
   wire n5040;
   wire n5041;
   wire n5042;
   wire n5043;
   wire n5044;
   wire n5045;
   wire n5046;
   wire n5047;
   wire n5048;
   wire n5049;
   wire n5050;
   wire n5051;
   wire n5052;
   wire n5053;
   wire n5055;
   wire n5056;
   wire n5057;
   wire n5058;
   wire n5059;
   wire n5060;
   wire n5061;
   wire n5062;
   wire n5063;
   wire n5064;
   wire n5065;
   wire n5066;
   wire n5067;
   wire n5068;
   wire n5069;
   wire n5070;
   wire n5071;
   wire n5072;
   wire n5073;
   wire n5074;
   wire n5075;
   wire n5076;
   wire n5077;
   wire n5078;
   wire n5079;
   wire n5080;
   wire n5081;
   wire n5082;
   wire n5083;
   wire n5084;
   wire n5085;
   wire n5086;
   wire n5087;
   wire n5088;
   wire n5089;
   wire n5090;
   wire n5091;
   wire n5092;
   wire n5093;
   wire n5094;
   wire n5095;
   wire n5096;
   wire n5097;
   wire n5098;
   wire n5099;
   wire n5100;
   wire n5101;
   wire n5102;
   wire n5103;
   wire n5104;
   wire n5105;
   wire n5106;
   wire n5107;
   wire n5108;
   wire n5109;
   wire n5110;
   wire n5111;
   wire n5112;
   wire n5113;
   wire n5114;
   wire n5115;
   wire n5116;
   wire n5117;
   wire n5118;
   wire n5120;
   wire n5121;
   wire n5122;
   wire n5123;
   wire n5124;
   wire n5125;
   wire n5126;
   wire n5127;
   wire n5128;
   wire n5129;
   wire n5130;
   wire n5131;
   wire n5132;
   wire n5133;
   wire n5134;
   wire n5135;
   wire n5136;
   wire n5137;
   wire n5138;
   wire n5139;
   wire n5140;
   wire n5141;
   wire n5142;
   wire n5143;
   wire n5144;
   wire n5145;
   wire n5146;
   wire n5147;
   wire n5148;
   wire n5149;
   wire n5150;
   wire n5151;
   wire n5152;
   wire n5153;
   wire n5154;
   wire n5155;
   wire n5156;
   wire n5157;
   wire n5158;
   wire n5159;
   wire n5160;
   wire n5161;
   wire n5162;
   wire n5165;
   wire n5167;
   wire n5168;
   wire n5169;
   wire n5170;
   wire n5171;
   wire n5172;
   wire n5173;
   wire n5174;
   wire n5175;
   wire n5176;
   wire n5177;
   wire n5178;
   wire n5179;
   wire n5180;
   wire n5181;
   wire n5182;
   wire n5183;
   wire n5184;
   wire n5185;
   wire n5186;
   wire n5187;
   wire n5188;
   wire n5189;
   wire n5190;
   wire n5191;
   wire n5192;
   wire n5193;
   wire n5194;
   wire n5195;
   wire n5196;
   wire n5197;
   wire n5198;
   wire n5199;
   wire n5200;
   wire n5201;
   wire n5202;
   wire n5203;
   wire n5204;
   wire n5205;
   wire n5206;
   wire n5207;
   wire n5208;
   wire n5209;
   wire n5210;
   wire n5211;
   wire n5212;
   wire n5213;
   wire n5214;
   wire n5215;
   wire n5216;
   wire n5217;
   wire n5218;
   wire n5219;
   wire n5220;
   wire n5221;
   wire n5222;
   wire n5223;
   wire n5224;
   wire n5225;
   wire n5226;
   wire n5227;
   wire n5228;
   wire n5229;
   wire n5230;
   wire n5231;
   wire n5233;
   wire n5234;
   wire n5235;
   wire n5236;
   wire n5237;
   wire n5238;
   wire n5239;
   wire n5240;
   wire n5241;
   wire n5243;
   wire n5244;
   wire n5252;
   wire n5253;
   wire n5254;
   wire n5255;
   wire n5256;
   wire n5257;
   wire n5258;
   wire n5259;
   wire n5260;
   wire n5261;
   wire n5262;
   wire n5263;
   wire n5264;
   wire n5265;
   wire n5266;
   wire n5267;
   wire n5268;
   wire n5269;
   wire n5270;
   wire n5271;
   wire n5272;
   wire n5273;
   wire n5274;
   wire n5275;
   wire n5276;
   wire n5277;
   wire n5278;
   wire n5279;
   wire n5280;
   wire n5281;
   wire n5282;
   wire n5283;
   wire n5284;
   wire n5285;
   wire n5286;
   wire n5287;
   wire n5288;
   wire n5289;
   wire n5290;
   wire n5291;
   wire n5292;
   wire n5293;
   wire n5294;
   wire n5295;
   wire n5296;
   wire n5297;
   wire n5298;
   wire n5299;
   wire n5300;
   wire n5301;
   wire n5302;
   wire n5303;
   wire n5304;
   wire n5305;
   wire n5306;
   wire n5307;
   wire n5308;
   wire n5309;
   wire n5310;
   wire n5311;
   wire n5312;
   wire n5313;
   wire n5314;
   wire n5315;
   wire n5316;
   wire n5317;
   wire n5318;
   wire n5319;
   wire n5320;
   wire n5321;
   wire n5322;
   wire n5323;
   wire n5324;
   wire n5325;
   wire n5326;
   wire n5327;
   wire n5328;
   wire n5329;
   wire n5330;
   wire n5331;
   wire n5332;
   wire n5333;
   wire n5334;
   wire n5335;
   wire n5336;
   wire n5337;
   wire n5338;
   wire n5339;
   wire n5340;
   wire n5341;
   wire n5342;
   wire n5343;
   wire n5344;
   wire n5345;
   wire n5346;
   wire n5347;
   wire n5348;
   wire n5349;
   wire n5350;
   wire n5351;
   wire n5352;
   wire n5353;
   wire n5354;
   wire n5355;
   wire n5356;
   wire n5357;
   wire n5358;
   wire n5359;
   wire n5360;
   wire n5361;
   wire n5362;
   wire n5363;
   wire n5364;
   wire n5365;
   wire n5366;
   wire n5367;
   wire n5368;
   wire n5369;
   wire n5370;
   wire n5371;
   wire n5372;
   wire n5373;
   wire n5374;
   wire n5375;
   wire n5376;
   wire n5377;
   wire n5378;
   wire n5379;
   wire n5380;
   wire n5381;
   wire n5382;
   wire n5383;
   wire n5384;
   wire n5385;
   wire n5386;
   wire n5387;
   wire n5388;
   wire n5389;
   wire n5390;
   wire n5391;
   wire n5392;
   wire n5393;
   wire n5394;
   wire n5395;
   wire n5396;
   wire n5397;
   wire n5398;
   wire n5399;
   wire n5400;
   wire n5401;
   wire n5402;
   wire n5403;
   wire n5404;
   wire n5405;
   wire n5406;
   wire n5407;
   wire n5408;
   wire n5409;
   wire n5410;
   wire n5411;
   wire n5412;
   wire n5413;
   wire n5414;
   wire n5415;
   wire n5416;
   wire n5417;
   wire n5418;
   wire n5419;
   wire n5420;
   wire n5421;
   wire n5422;
   wire n5423;
   wire n5424;
   wire n5425;
   wire n5426;
   wire n5427;
   wire n5428;
   wire n5429;
   wire n5430;
   wire n5431;
   wire n5432;
   wire n5433;
   wire n5434;
   wire n5435;
   wire n5436;
   wire n5437;
   wire n5438;
   wire n5439;
   wire n5440;
   wire n5441;
   wire n5442;
   wire n5443;
   wire n5444;
   wire n5445;
   wire n5446;
   wire n5447;
   wire n5448;
   wire n5449;
   wire n5450;
   wire n5451;
   wire n5452;
   wire n5453;
   wire n5454;
   wire n5455;
   wire n5456;
   wire n5457;
   wire n5458;
   wire n5459;
   wire n5460;
   wire n5461;
   wire n5462;
   wire n5463;
   wire n5464;
   wire n5465;
   wire n5466;
   wire n5467;
   wire n5468;
   wire n5469;
   wire n5470;
   wire n5471;
   wire n5472;
   wire n5473;
   wire n5474;
   wire n5475;
   wire n5476;
   wire n5477;
   wire n5478;
   wire n5479;
   wire n5480;
   wire n5481;
   wire n5482;
   wire n5483;
   wire n5484;
   wire n5485;
   wire n5486;
   wire n5487;
   wire n5488;
   wire n5489;
   wire n5490;
   wire n5491;
   wire n5492;
   wire n5493;
   wire n5494;
   wire n5495;
   wire n5496;
   wire n5497;
   wire n5498;
   wire n5499;
   wire n5500;
   wire n5501;
   wire n5502;
   wire n5503;
   wire n5504;
   wire n5505;
   wire n5506;
   wire n5507;
   wire n5508;
   wire n5509;
   wire n5510;
   wire n5511;
   wire n5512;
   wire n5513;
   wire n5514;
   wire n5515;
   wire n5516;
   wire n5517;
   wire n5518;
   wire n5519;
   wire n5520;
   wire n5521;
   wire n5522;
   wire n5523;
   wire n5524;
   wire n5525;
   wire n5526;
   wire n5527;
   wire n5528;
   wire n5529;
   wire n5530;
   wire n5531;
   wire n5532;
   wire n5533;
   wire n5534;
   wire n5535;
   wire n5536;
   wire n5537;
   wire n5538;
   wire n5539;
   wire n5540;
   wire n5541;
   wire n5542;
   wire n5543;
   wire n5544;
   wire n5545;
   wire n5546;
   wire n5547;
   wire n5548;
   wire n5549;
   wire n5550;
   wire n5551;
   wire n5552;
   wire n5553;
   wire n5554;
   wire n5555;
   wire n5556;
   wire n5557;
   wire n5558;
   wire n5559;
   wire n5560;
   wire n5561;
   wire n5562;
   wire n5563;
   wire n5564;
   wire n5565;
   wire n5566;
   wire n5567;
   wire n5568;
   wire n5569;
   wire n5570;
   wire n5571;
   wire n5572;
   wire n5573;
   wire n5574;
   wire n5575;
   wire n5576;
   wire n5577;
   wire n5578;
   wire n5579;
   wire n5580;
   wire n5581;
   wire n5582;
   wire n5583;
   wire n5584;
   wire n5585;
   wire n5586;
   wire n5587;
   wire n5588;
   wire n5589;
   wire n5590;
   wire n5591;
   wire n5592;
   wire n5593;
   wire n5594;
   wire n5595;
   wire n5596;
   wire n5597;
   wire n5598;
   wire n5599;
   wire n5600;
   wire n5601;
   wire n5602;
   wire n5603;
   wire n5604;
   wire n5605;
   wire n5606;
   wire n5607;
   wire n5608;
   wire n5609;
   wire n5610;
   wire n5611;
   wire n5612;
   wire n5613;
   wire n5614;
   wire n5615;
   wire n5616;
   wire n5617;
   wire n5618;
   wire n5619;
   wire n5620;
   wire n5621;
   wire n5622;
   wire n5623;
   wire n5624;
   wire n5625;
   wire n5626;
   wire n5627;
   wire n5628;
   wire n5629;
   wire n5630;
   wire n5631;
   wire n5632;
   wire n5633;
   wire n5634;
   wire n5635;
   wire n5636;
   wire n5637;
   wire n5638;
   wire n5639;
   wire n5640;
   wire n5641;
   wire n5642;
   wire n5643;
   wire n5644;
   wire n5645;
   wire n5646;
   wire n5647;
   wire n5648;
   wire n5649;
   wire n5650;
   wire n5651;
   wire n5652;
   wire n5653;
   wire n5654;
   wire n5655;
   wire n5656;
   wire n5657;
   wire n5658;
   wire n5659;
   wire n5660;
   wire n5661;
   wire n5662;
   wire n5663;
   wire n5664;
   wire n5665;
   wire n5666;
   wire n5667;
   wire n5668;
   wire n5669;
   wire n5670;
   wire n5671;
   wire n5672;
   wire n5673;
   wire n5674;
   wire n5675;
   wire n5676;
   wire n5677;
   wire n5678;
   wire n5679;
   wire n5680;
   wire n5681;
   wire n5682;
   wire n5683;
   wire n5684;
   wire n5685;
   wire n5686;
   wire n5687;
   wire n5688;
   wire n5689;
   wire n5690;
   wire n5691;
   wire n5692;
   wire n5693;
   wire n5694;
   wire n5695;
   wire n5696;
   wire n5697;
   wire n5698;
   wire n5699;
   wire n5700;
   wire n5701;
   wire n5702;
   wire n5703;
   wire n5704;
   wire n5705;
   wire n5706;
   wire n5707;
   wire n5708;
   wire n5709;
   wire n5710;
   wire n5711;
   wire n5712;
   wire n5713;
   wire n5714;
   wire n5715;
   wire n5716;
   wire n5717;
   wire n5718;
   wire n5719;
   wire n5720;
   wire n5721;
   wire n5722;
   wire n5723;
   wire n5724;
   wire n5725;
   wire n5726;
   wire n5727;
   wire n5728;
   wire n5729;
   wire n5730;
   wire n5731;
   wire n5732;
   wire n5733;
   wire n5734;
   wire n5735;
   wire n5736;
   wire n5737;
   wire n5738;
   wire n5739;
   wire n5740;
   wire n5741;
   wire n5742;
   wire n5743;
   wire n5744;
   wire n5745;
   wire n5746;
   wire n5747;
   wire n5748;
   wire n5749;
   wire n5750;
   wire n5751;
   wire n5752;
   wire n5753;
   wire n5754;
   wire n5755;
   wire n5756;
   wire n5757;
   wire n5758;
   wire n5759;
   wire n5760;
   wire n5761;
   wire n5762;
   wire n5763;
   wire n5764;
   wire n5765;
   wire n5766;
   wire n5767;
   wire n5768;
   wire n5769;
   wire n5770;
   wire n5771;
   wire n5772;
   wire n5773;
   wire n5774;
   wire n5775;
   wire n5776;
   wire n5777;
   wire n5778;
   wire n5779;
   wire n5780;
   wire n5781;
   wire n5782;
   wire n5783;
   wire n5784;
   wire n5785;
   wire n5786;
   wire n5787;
   wire n5788;
   wire n5789;
   wire n5790;
   wire n5791;
   wire n5792;
   wire n5793;
   wire n5794;
   wire n5795;
   wire n5796;
   wire n5797;
   wire n5798;
   wire n5799;
   wire n5800;
   wire n5801;
   wire n5802;
   wire n5803;
   wire n5804;
   wire n5805;
   wire n5806;
   wire n5807;
   wire n5808;
   wire n5809;
   wire n5810;
   wire n5811;
   wire n5812;
   wire n5813;
   wire n5814;
   wire n5815;
   wire n5816;
   wire n5817;
   wire n5818;
   wire n5819;
   wire n5820;
   wire n5821;
   wire n5822;
   wire n5823;
   wire n5824;
   wire n5825;
   wire n5826;
   wire n5827;
   wire n5828;
   wire n5829;
   wire n16644;
   wire n16645;
   wire n16646;
   wire n16647;
   wire n16648;
   wire n16649;
   wire n16650;
   wire n16651;
   wire n16652;
   wire n16653;
   wire n16654;
   wire n16655;
   wire n16656;
   wire n16657;
   wire n16658;
   wire n16659;
   wire n16660;
   wire n16661;
   wire n16662;
   wire n16663;
   wire n16664;
   wire n16665;
   wire n16666;
   wire n16667;
   wire n16668;
   wire n16669;
   wire n16670;
   wire n16671;
   wire n16672;
   wire n16673;
   wire n16674;
   wire n16675;
   wire n16676;
   wire n16677;
   wire n16678;
   wire n16679;
   wire n16680;
   wire n16681;
   wire n16682;
   wire n16683;
   wire n16684;
   wire n16685;
   wire n16686;
   wire n16687;
   wire n16688;
   wire n16689;
   wire n16690;
   wire n16691;
   wire n16692;
   wire n16693;
   wire n16694;
   wire n16695;
   wire n16696;
   wire n16697;
   wire n16698;
   wire n16699;
   wire n16700;
   wire n16701;
   wire n16702;
   wire n16703;
   wire n16704;
   wire n16705;
   wire n16706;
   wire n16707;
   wire n16708;
   wire n16709;
   wire n16710;
   wire n16711;
   wire n16712;
   wire n16713;
   wire n16714;
   wire n16715;
   wire n16716;
   wire n16717;
   wire n16718;
   wire n16719;
   wire n16720;
   wire n16721;
   wire n16722;
   wire n16723;
   wire n16725;
   wire n16726;
   wire n16727;
   wire n16728;
   wire n16729;
   wire n16730;
   wire n16731;
   wire n16732;
   wire n16733;
   wire n16734;
   wire n16735;
   wire n16736;
   wire n16737;
   wire n16738;
   wire n16739;
   wire n16740;
   wire n16741;
   wire n16742;
   wire n16743;
   wire n16744;
   wire n16745;
   wire n16746;
   wire n16747;
   wire n16748;
   wire n16749;
   wire n16750;
   wire n16751;
   wire n16752;
   wire n16753;
   wire n16754;
   wire n16755;
   wire n16756;
   wire n16757;
   wire n16758;
   wire n16759;
   wire n16760;
   wire n16761;
   wire n16762;
   wire n16763;
   wire n16764;
   wire n16765;
   wire n16766;
   wire n16767;
   wire n16768;
   wire n16769;
   wire n16770;
   wire n16771;
   wire n16772;
   wire n16773;
   wire n16774;
   wire n16775;
   wire n16776;
   wire n16777;
   wire n16778;
   wire n16779;
   wire n16780;
   wire n16781;
   wire n16782;
   wire n16783;
   wire n16784;
   wire n16785;
   wire n16787;
   wire n16788;
   wire n16792;
   wire n16794;
   wire n16795;
   wire n16796;
   wire n16797;
   wire n16798;
   wire n16799;
   wire n16800;
   wire n16801;
   wire n16802;
   wire n16803;
   wire n16804;
   wire n16805;
   wire n16806;
   wire n16807;
   wire n16808;
   wire n16809;
   wire n16810;
   wire n16811;
   wire n16812;
   wire n16813;
   wire n16814;
   wire n16816;
   wire n16817;
   wire n16818;
   wire n16820;
   wire n16821;
   wire n16822;
   wire n16824;
   wire n16825;
   wire n16826;
   wire n16827;
   wire n16828;
   wire n16831;
   wire n16833;
   wire n16834;
   wire n16835;
   wire n16836;
   wire n16837;
   wire n16838;
   wire n16839;
   wire n16840;
   wire n16842;
   wire n16843;
   wire n16844;
   wire n16845;
   wire n16846;
   wire n16847;
   wire n16848;
   wire n16849;
   wire n16850;
   wire n16851;
   wire n16852;
   wire n16854;
   wire n16855;
   wire n16856;
   wire n16857;
   wire n16859;
   wire n16860;
   wire n16861;
   wire n16862;
   wire n16863;
   wire n16864;
   wire n16865;
   wire n16867;
   wire n16868;
   wire n16870;
   wire n16871;
   wire n16872;
   wire n16873;
   wire n16875;
   wire n16877;
   wire n16882;
   wire n16885;
   wire n16886;
   wire n16891;
   wire n16893;
   wire n16895;
   wire n16897;
   wire n16902;
   wire n16905;
   wire n16908;
   wire n16910;
   wire n16911;
   wire n16913;
   wire n16916;
   wire n16918;
   wire n16919;
   wire n16921;
   wire n16922;
   wire n16924;
   wire n16925;
   wire n16927;
   wire n16930;
   wire n16931;
   wire n16933;
   wire n16934;
   wire n16936;
   wire n16939;
   wire n16942;
   wire n16945;
   wire n16948;
   wire n16951;
   wire n16954;
   wire n16955;
   wire n16956;
   wire n16957;
   wire n16958;
   wire n16959;
   wire n16960;
   wire n16961;
   wire n16962;
   wire n16963;
   wire n16964;
   wire n16965;
   wire n16966;
   wire n16967;
   wire n16968;
   wire n16969;
   wire n16970;
   wire n16971;
   wire n16972;
   wire n16973;
   wire n16974;
   wire n16975;
   wire n16976;
   wire n16977;
   wire n16979;
   wire n16980;
   wire n16982;
   wire n16983;
   wire n16984;
   wire n16985;
   wire n16986;
   wire n16987;
   wire n16988;
   wire n16989;
   wire n16990;
   wire n16991;
   wire n16992;
   wire n16994;
   wire n16996;
   wire n17000;
   wire n17001;
   wire n17005;
   wire n17008;
   wire n17013;
   wire n17017;
   wire n17018;
   wire n17022;
   wire n17023;
   wire n17027;
   wire n17028;
   wire n17031;
   wire n17033;
   wire n17037;
   wire n17038;
   wire n17042;
   wire n17043;
   wire n17046;
   wire n17048;
   wire n17052;
   wire n17053;
   wire n17057;
   wire n17058;
   wire n17062;
   wire n17063;
   wire n17067;
   wire n17068;
   wire n17071;
   wire n17074;
   wire n17077;
   wire n17078;
   wire n17082;
   wire n17083;
   wire n17088;
   wire n17090;
   wire n17092;
   wire n17094;
   wire n17095;
   wire n17096;
   wire n17097;
   wire n17098;
   wire n17099;
   wire n17102;
   wire n17103;
   wire n17104;
   wire n17106;
   wire n17107;
   wire n17108;
   wire n17109;
   wire n17116;
   wire n17117;
   wire n17120;
   wire n17122;
   wire n17124;
   wire n17126;
   wire n17127;
   wire [33:3] add_2082_carry;
   wire [29:2] add_2072_carry;
   wire [30:2] add_2071_carry;

   BUF_X4 FE_PSC671_n2057 (.Z(FE_PSN5239_n2057), 
	.A(n2057));
   BUF_X4 FE_PSC670_n3097 (.Z(FE_PSN5238_n3097), 
	.A(n3097));
   CLKBUF_X3 FE_PSC669_n2184 (.Z(FE_PSN5237_n2184), 
	.A(n2184));
   CLKBUF_X3 FE_PSC668_n16960 (.Z(FE_PSN5236_n16960), 
	.A(n16960));
   BUF_X1 FE_PHC5254_n1134 (.Z(FE_PHN5254_n1134), 
	.A(FE_PHN5245_n1134));
   CLKBUF_X1 FE_PHC5252_n389 (.Z(FE_PHN5252_n389), 
	.A(n389));
   CLKBUF_X1 FE_PHC5251_n5743 (.Z(FE_PHN5251_n5743), 
	.A(FE_PHN717_n5743));
   CLKBUF_X1 FE_PHC5250_n5747 (.Z(FE_PHN5250_n5747), 
	.A(FE_PHN707_n5747));
   CLKBUF_X1 FE_PHC5249_n5740 (.Z(FE_PHN5249_n5740), 
	.A(FE_PHN722_n5740));
   CLKBUF_X1 FE_PHC5248_n395 (.Z(FE_PHN5248_n395), 
	.A(n395));
   CLKBUF_X1 FE_PHC5247_n14432 (.Z(FE_PHN5247_n14432), 
	.A(FE_PHN928_n14432));
   BUF_X8 FE_PHC5246_n1137 (.Z(FE_PHN5246_n1137), 
	.A(n1137));
   CLKBUF_X1 FE_PHC5245_n1134 (.Z(FE_PHN5245_n1134), 
	.A(n1134));
   CLKBUF_X1 FE_PHC5244_n4915 (.Z(FE_PHN5244_n4915), 
	.A(FE_PHN5204_n4915));
   CLKBUF_X1 FE_PHC5243_n5745 (.Z(FE_PHN5243_n5745), 
	.A(FE_PHN738_n5745));
   CLKBUF_X1 FE_PHC5242_n5749 (.Z(FE_PHN5242_n5749), 
	.A(FE_PHN721_n5749));
   CLKBUF_X1 FE_PHC5238_n5748 (.Z(FE_PHN5238_n5748), 
	.A(FE_PHN733_n5748));
   BUF_X8 FE_PHC5236_n5742 (.Z(FE_PHN5236_n5742), 
	.A(FE_PHN701_n5742));
   BUF_X32 FE_PHC5233_n5760 (.Z(FE_PHN5233_n5760), 
	.A(FE_PHN830_n5760));
   BUF_X32 FE_PHC5232_n385 (.Z(FE_PHN5232_n385), 
	.A(n385));
   BUF_X32 FE_PHC5231_n1136 (.Z(FE_PHN5231_n1136), 
	.A(n1136));
   BUF_X32 FE_PHC5230_n419 (.Z(FE_PHN5230_n419), 
	.A(n419));
   BUF_X32 FE_PHC5229_n1135 (.Z(FE_PHN5229_n1135), 
	.A(n1135));
   BUF_X32 FE_PHC5228_n1141 (.Z(FE_PHN5228_n1141), 
	.A(n1141));
   BUF_X32 FE_PHC5227_n1138 (.Z(FE_PHN5227_n1138), 
	.A(n1138));
   CLKBUF_X1 FE_PHC5226_U227_Z_0 (.Z(FE_PHN5226_U227_Z_0), 
	.A(U227_Z_0));
   BUF_X16 FE_PHC5225_n5746 (.Z(FE_PHN5225_n5746), 
	.A(n5746));
   BUF_X16 FE_PHC5224_n5751 (.Z(FE_PHN5224_n5751), 
	.A(FE_PHN739_n5751));
   BUF_X32 FE_PHC5223_n5752 (.Z(FE_PHN5223_n5752), 
	.A(FE_PHN704_n5752));
   BUF_X32 FE_PHC5222_n5750 (.Z(FE_PHN5222_n5750), 
	.A(FE_PHN730_n5750));
   BUF_X32 FE_PHC5221_n5763 (.Z(FE_PHN5221_n5763), 
	.A(FE_PHN852_n5763));
   BUF_X32 FE_PHC5220_n5754 (.Z(FE_PHN5220_n5754), 
	.A(FE_PHN715_n5754));
   BUF_X32 FE_PHC5219_n5756 (.Z(FE_PHN5219_n5756), 
	.A(FE_PHN829_n5756));
   BUF_X32 FE_PHC5217_n380 (.Z(FE_PHN5217_n380), 
	.A(n380));
   BUF_X32 FE_PHC5216_n1146 (.Z(FE_PHN5216_n1146), 
	.A(n1146));
   BUF_X32 FE_PHC5215_n387 (.Z(FE_PHN5215_n387), 
	.A(n387));
   BUF_X32 FE_PHC5214_n1133 (.Z(FE_PHN5214_n1133), 
	.A(n1133));
   BUF_X32 FE_PHC5213_n1132 (.Z(FE_PHN5213_n1132), 
	.A(n1132));
   BUF_X32 FE_PHC5212_n1130 (.Z(FE_PHN5212_n1130), 
	.A(n1130));
   BUF_X32 FE_PHC5211_n1139 (.Z(FE_PHN5211_n1139), 
	.A(n1139));
   BUF_X32 FE_PHC5210_n395 (.Z(FE_PHN5210_n395), 
	.A(FE_PHN5248_n395));
   BUF_X32 FE_PHC5209_n14432 (.Z(FE_PHN5209_n14432), 
	.A(FE_PHN5247_n14432));
   BUF_X32 FE_PHC5208_n389 (.Z(FE_PHN5208_n389), 
	.A(FE_PHN5252_n389));
   BUF_X32 FE_PHC5207_n1134 (.Z(FE_PHN5207_n1134), 
	.A(FE_PHN5254_n1134));
   BUF_X32 FE_PHC5206_n1137 (.Z(FE_PHN5206_n1137), 
	.A(FE_PHN5246_n1137));
   CLKBUF_X1 FE_PHC5205_n5761 (.Z(FE_PHN5205_n5761), 
	.A(FE_PHN1038_n5761));
   CLKBUF_X1 FE_PHC5204_n4915 (.Z(FE_PHN5204_n4915), 
	.A(FE_PHN846_n4915));
   BUF_X32 FE_PHC5202_n5741 (.Z(FE_PHN5202_n5741), 
	.A(FE_PHN723_n5741));
   BUF_X32 FE_PHC5201_n5744 (.Z(FE_PHN5201_n5744), 
	.A(FE_PHN737_n5744));
   BUF_X32 FE_PHC5200_n5753 (.Z(FE_PHN5200_n5753), 
	.A(FE_PHN716_n5753));
   BUF_X32 FE_PHC5199_n5766 (.Z(FE_PHN5199_n5766), 
	.A(FE_PHN1010_n5766));
   BUF_X32 FE_PHC5198_n5739 (.Z(FE_PHN5198_n5739), 
	.A(FE_PHN720_n5739));
   BUF_X32 FE_PHC5197_n5765 (.Z(FE_PHN5197_n5765), 
	.A(FE_PHN1009_n5765));
   BUF_X32 FE_PHC5196_n5745 (.Z(FE_PHN5196_n5745), 
	.A(FE_PHN5243_n5745));
   BUF_X32 FE_PHC5195_n5749 (.Z(FE_PHN5195_n5749), 
	.A(FE_PHN5242_n5749));
   BUF_X32 FE_PHC5194_n5742 (.Z(FE_PHN5194_n5742), 
	.A(FE_PHN5236_n5742));
   BUF_X1 FE_PHC5193_n4389 (.Z(FE_PHN5193_n4389), 
	.A(FE_PHN4673_n4389));
   CLKBUF_X1 FE_PHC5192_n17126 (.Z(FE_PHN5192_n17126), 
	.A(FE_PHN2911_n17126));
   BUF_X32 FE_PHC5188_n5768 (.Z(FE_PHN5188_n5768), 
	.A(FE_PHN1007_n5768));
   BUF_X32 FE_PHC5187_n5767 (.Z(FE_PHN5187_n5767), 
	.A(FE_PHN1008_n5767));
   BUF_X32 FE_PHC5186_n5769 (.Z(FE_PHN5186_n5769), 
	.A(FE_PHN1006_n5769));
   BUF_X32 FE_PHC5185_n5743 (.Z(FE_PHN5185_n5743), 
	.A(FE_PHN5251_n5743));
   BUF_X32 FE_PHC5184_n5748 (.Z(FE_PHN5184_n5748), 
	.A(FE_PHN5238_n5748));
   BUF_X32 FE_PHC5183_n5747 (.Z(FE_PHN5183_n5747), 
	.A(FE_PHN5250_n5747));
   BUF_X32 FE_PHC5182_n5740 (.Z(FE_PHN5182_n5740), 
	.A(FE_PHN5249_n5740));
   CLKBUF_X1 FE_PHC5178_IRQ_15_ (.Z(FE_PHN5178_IRQ_15_), 
	.A(FE_PHN4630_IRQ_15_));
   BUF_X1 FE_PHC5177_IRQ_11_ (.Z(FE_PHN5177_IRQ_11_), 
	.A(FE_PHN4638_IRQ_11_));
   CLKBUF_X1 FE_PHC5170_U591_Z_0 (.Z(FE_PHN5170_U591_Z_0), 
	.A(FE_PHN2085_U591_Z_0));
   CLKBUF_X1 FE_PHC5169_n5349 (.Z(FE_PHN5169_n5349), 
	.A(FE_PHN4090_n5349));
   CLKBUF_X1 FE_PHC5168_n5352 (.Z(FE_PHN5168_n5352), 
	.A(FE_PHN4089_n5352));
   CLKBUF_X1 FE_PHC5167_n5081 (.Z(FE_PHN5167_n5081), 
	.A(FE_PHN4258_n5081));
   CLKBUF_X1 FE_PHC5166_U503_Z_0 (.Z(FE_PHN5166_U503_Z_0), 
	.A(FE_PHN3868_U503_Z_0));
   CLKBUF_X1 FE_PHC5163_n5262 (.Z(FE_PHN5163_n5262), 
	.A(FE_PHN3886_n5262));
   CLKBUF_X1 FE_PHC5161_n4874 (.Z(FE_PHN5161_n4874), 
	.A(FE_PHN4133_n4874));
   CLKBUF_X1 FE_PHC5160_n5362 (.Z(FE_PHN5160_n5362), 
	.A(FE_PHN4150_n5362));
   CLKBUF_X1 FE_PHC5158_n4979 (.Z(FE_PHN5158_n4979), 
	.A(FE_PHN4219_n4979));
   CLKBUF_X1 FE_PHC5156_n5361 (.Z(FE_PHN5156_n5361), 
	.A(FE_PHN4220_n5361));
   CLKBUF_X1 FE_PHC5155_n5483 (.Z(FE_PHN5155_n5483), 
	.A(FE_PHN4266_n5483));
   CLKBUF_X2 FE_PHC5151_n5128 (.Z(FE_PHN5151_n5128), 
	.A(FE_PHN4032_n5128));
   CLKBUF_X2 FE_PHC5150_n5378 (.Z(FE_PHN5150_n5378), 
	.A(FE_PHN4057_n5378));
   CLKBUF_X2 FE_PHC5149_n5347 (.Z(FE_PHN5149_n5347), 
	.A(FE_PHN4083_n5347));
   CLKBUF_X2 FE_PHC5146_n5159 (.Z(FE_PHN5146_n5159), 
	.A(FE_PHN4271_n5159));
   BUF_X1 FE_PHC5145_U769_Z_0 (.Z(FE_PHN5145_U769_Z_0), 
	.A(FE_PHN3869_U769_Z_0));
   CLKBUF_X1 FE_PHC5141_n4875 (.Z(FE_PHN5141_n4875), 
	.A(FE_PHN3934_n4875));
   CLKBUF_X1 FE_PHC5139_n5319 (.Z(FE_PHN5139_n5319), 
	.A(FE_PHN4170_n5319));
   CLKBUF_X1 FE_PHC5137_n5610 (.Z(FE_PHN5137_n5610), 
	.A(FE_PHN4180_n5610));
   CLKBUF_X1 FE_PHC5136_n5360 (.Z(FE_PHN5136_n5360), 
	.A(FE_PHN4221_n5360));
   CLKBUF_X1 FE_PHC5135_n5391 (.Z(FE_PHN5135_n5391), 
	.A(FE_PHN4213_n5391));
   CLKBUF_X1 FE_PHC5134_n5413 (.Z(FE_PHN5134_n5413), 
	.A(FE_PHN4235_n5413));
   BUF_X1 FE_PHC5131_U247_Z_0 (.Z(FE_PHN5131_U247_Z_0), 
	.A(FE_PHN1741_U247_Z_0));
   CLKBUF_X2 FE_PHC5130_n5369 (.Z(FE_PHN5130_n5369), 
	.A(FE_PHN4199_n5369));
   CLKBUF_X2 FE_PHC5129_n5491 (.Z(FE_PHN5129_n5491), 
	.A(FE_PHN4059_n5491));
   BUF_X1 FE_PHC5127_n5018 (.Z(FE_PHN5127_n5018), 
	.A(FE_PHN4191_n5018));
   CLKBUF_X2 FE_PHC5126_n5280 (.Z(FE_PHN5126_n5280), 
	.A(FE_PHN4165_n5280));
   BUF_X1 FE_PHC5125_n5443 (.Z(FE_PHN5125_n5443), 
	.A(FE_PHN4231_n5443));
   CLKBUF_X2 FE_PHC5124_n5308 (.Z(FE_PHN5124_n5308), 
	.A(FE_PHN4249_n5308));
   CLKBUF_X1 FE_PHC5123_n4848 (.Z(FE_PHN5123_n4848), 
	.A(FE_PHN3620_n4848));
   CLKBUF_X1 FE_PHC5122_n5052 (.Z(FE_PHN5122_n5052), 
	.A(FE_PHN4040_n5052));
   CLKBUF_X1 FE_PHC5121_n5089 (.Z(FE_PHN5121_n5089), 
	.A(FE_PHN4058_n5089));
   CLKBUF_X1 FE_PHC5120_n5617 (.Z(FE_PHN5120_n5617), 
	.A(FE_PHN4021_n5617));
   CLKBUF_X1 FE_PHC5119_U528_Z_0 (.Z(FE_PHN5119_U528_Z_0), 
	.A(FE_PHN2057_U528_Z_0));
   CLKBUF_X1 FE_PHC5114_n5279 (.Z(FE_PHN5114_n5279), 
	.A(FE_PHN4147_n5279));
   CLKBUF_X1 FE_PHC5113_U761_Z_0 (.Z(FE_PHN5113_U761_Z_0), 
	.A(FE_PHN4229_U761_Z_0));
   CLKBUF_X2 FE_PHC5108_n5133 (.Z(FE_PHN5108_n5133), 
	.A(FE_PHN4166_n5133));
   CLKBUF_X2 FE_PHC5107_n5538 (.Z(FE_PHN5107_n5538), 
	.A(FE_PHN4205_n5538));
   CLKBUF_X2 FE_PHC5106_n5364 (.Z(FE_PHN5106_n5364), 
	.A(FE_PHN4240_n5364));
   BUF_X1 FE_PHC5105_n5204 (.Z(FE_PHN5105_n5204), 
	.A(FE_PHN3921_n5204));
   CLKBUF_X1 FE_PHC5104_U583_Z_0 (.Z(FE_PHN5104_U583_Z_0), 
	.A(FE_PHN2088_U583_Z_0));
   CLKBUF_X1 FE_PHC5099_n5611 (.Z(FE_PHN5099_n5611), 
	.A(FE_PHN4139_n5611));
   CLKBUF_X1 FE_PHC5097_U646_Z_0 (.Z(FE_PHN5097_U646_Z_0), 
	.A(FE_PHN3863_U646_Z_0));
   CLKBUF_X1 FE_PHC5096_U428_Z_0 (.Z(FE_PHN5096_U428_Z_0), 
	.A(FE_PHN3864_U428_Z_0));
   CLKBUF_X1 FE_PHC5094_n5142 (.Z(FE_PHN5094_n5142), 
	.A(FE_PHN3874_n5142));
   CLKBUF_X1 FE_PHC5093_n5220 (.Z(FE_PHN5093_n5220), 
	.A(FE_PHN4031_n5220));
   CLKBUF_X1 FE_PHC5091_U359_Z_0 (.Z(FE_PHN5091_U359_Z_0), 
	.A(FE_PHN4232_U359_Z_0));
   CLKBUF_X1 FE_PHC5090_n5201 (.Z(FE_PHN5090_n5201), 
	.A(FE_PHN4129_n5201));
   CLKBUF_X1 FE_PHC5089_U644_Z_0 (.Z(FE_PHN5089_U644_Z_0), 
	.A(FE_PHN3903_U644_Z_0));
   CLKBUF_X2 FE_PHC5088_n5355 (.Z(FE_PHN5088_n5355), 
	.A(FE_PHN4052_n5355));
   CLKBUF_X2 FE_PHC5086_n5202 (.Z(FE_PHN5086_n5202), 
	.A(FE_PHN4218_n5202));
   BUF_X1 FE_PHC5085_n5337 (.Z(FE_PHN5085_n5337), 
	.A(FE_PHN4026_n5337));
   CLKBUF_X2 FE_PHC5084_U275_Z_0 (.Z(FE_PHN5084_U275_Z_0), 
	.A(FE_PHN4196_U275_Z_0));
   BUF_X1 FE_PHC5080_U711_Z_0 (.Z(FE_PHN5080_U711_Z_0), 
	.A(FE_PHN3862_U711_Z_0));
   CLKBUF_X1 FE_PHC5077_U589_Z_0 (.Z(FE_PHN5077_U589_Z_0), 
	.A(FE_PHN2069_U589_Z_0));
   CLKBUF_X1 FE_PHC5076_U595_Z_0 (.Z(FE_PHN5076_U595_Z_0), 
	.A(FE_PHN2062_U595_Z_0));
   CLKBUF_X1 FE_PHC5074_n5260 (.Z(FE_PHN5074_n5260), 
	.A(FE_PHN3982_n5260));
   CLKBUF_X1 FE_PHC5066_n5653 (.Z(FE_PHN5066_n5653), 
	.A(FE_PHN1875_n5653));
   CLKBUF_X1 FE_PHC5065_n5223 (.Z(FE_PHN5065_n5223), 
	.A(FE_PHN3571_n5223));
   CLKBUF_X1 FE_PHC5061_n5042 (.Z(FE_PHN5061_n5042), 
	.A(FE_PHN3973_n5042));
   CLKBUF_X1 FE_PHC5060_n5136 (.Z(FE_PHN5060_n5136), 
	.A(FE_PHN4168_n5136));
   CLKBUF_X1 FE_PHC5059_n5367 (.Z(FE_PHN5059_n5367), 
	.A(FE_PHN4172_n5367));
   CLKBUF_X2 FE_PHC5055_n5209 (.Z(FE_PHN5055_n5209), 
	.A(FE_PHN4198_n5209));
   BUF_X1 FE_PHC5053_n5271 (.Z(FE_PHN5053_n5271), 
	.A(FE_PHN4044_n5271));
   BUF_X1 FE_PHC5052_n5383 (.Z(FE_PHN5052_n5383), 
	.A(FE_PHN4148_n5383));
   CLKBUF_X2 FE_PHC5050_n5511 (.Z(FE_PHN5050_n5511), 
	.A(FE_PHN4185_n5511));
   CLKBUF_X1 FE_PHC5049_U677_Z_0 (.Z(FE_PHN5049_U677_Z_0), 
	.A(FE_PHN3856_U677_Z_0));
   CLKBUF_X1 FE_PHC5046_n4963 (.Z(FE_PHN5046_n4963), 
	.A(FE_PHN3883_n4963));
   CLKBUF_X1 FE_PHC5045_n5200 (.Z(FE_PHN5045_n5200), 
	.A(FE_PHN4175_n5200));
   CLKBUF_X1 FE_PHC5044_n5339 (.Z(FE_PHN5044_n5339), 
	.A(FE_PHN4135_n5339));
   CLKBUF_X1 FE_PHC5043_n4878 (.Z(FE_PHN5043_n4878), 
	.A(FE_PHN4104_n4878));
   CLKBUF_X1 FE_PHC5039_U441_Z_0 (.Z(FE_PHN5039_U441_Z_0), 
	.A(FE_PHN4039_U441_Z_0));
   CLKBUF_X1 FE_PHC5035_n5602 (.Z(FE_PHN5035_n5602), 
	.A(FE_PHN4012_n5602));
   CLKBUF_X1 FE_PHC5034_n5104 (.Z(FE_PHN5034_n5104), 
	.A(FE_PHN4002_n5104));
   CLKBUF_X1 FE_PHC5031_U784_Z_0 (.Z(FE_PHN5031_U784_Z_0), 
	.A(FE_PHN4202_U784_Z_0));
   CLKBUF_X1 FE_PHC5029_n5084 (.Z(FE_PHN5029_n5084), 
	.A(FE_PHN4117_n5084));
   CLKBUF_X1 FE_PHC5028_n4995 (.Z(FE_PHN5028_n4995), 
	.A(FE_PHN4187_n4995));
   CLKBUF_X1 FE_PHC5027_n5384 (.Z(FE_PHN5027_n5384), 
	.A(FE_PHN4192_n5384));
   CLKBUF_X1 FE_PHC5026_U363_Z_0 (.Z(FE_PHN5026_U363_Z_0), 
	.A(FE_PHN3857_U363_Z_0));
   BUF_X1 FE_PHC5025_U309_Z_0 (.Z(FE_PHN5025_U309_Z_0), 
	.A(FE_PHN2058_U309_Z_0));
   BUF_X1 FE_PHC5023_n5381 (.Z(FE_PHN5023_n5381), 
	.A(FE_PHN3974_n5381));
   BUF_X1 FE_PHC5019_n5492 (.Z(FE_PHN5019_n5492), 
	.A(FE_PHN4094_n5492));
   BUF_X1 FE_PHC5018_n5493 (.Z(FE_PHN5018_n5493), 
	.A(FE_PHN4093_n5493));
   BUF_X1 FE_PHC5017_n5221 (.Z(FE_PHN5017_n5221), 
	.A(FE_PHN4072_n5221));
   BUF_X1 FE_PHC5015_n5489 (.Z(FE_PHN5015_n5489), 
	.A(FE_PHN4122_n5489));
   BUF_X1 FE_PHC5014_n5294 (.Z(FE_PHN5014_n5294), 
	.A(FE_PHN4119_n5294));
   CLKBUF_X1 FE_PHC5013_n5307 (.Z(FE_PHN5013_n5307), 
	.A(FE_PHN3943_n5307));
   CLKBUF_X1 FE_PHC5010_n4924 (.Z(FE_PHN5010_n4924), 
	.A(FE_PHN1934_n4924));
   CLKBUF_X1 FE_PHC5008_n5019 (.Z(FE_PHN5008_n5019), 
	.A(FE_PHN4171_n5019));
   CLKBUF_X1 FE_PHC5006_n5640 (.Z(FE_PHN5006_n5640), 
	.A(FE_PHN4136_n5640));
   CLKBUF_X1 FE_PHC5002_n5643 (.Z(FE_PHN5002_n5643), 
	.A(FE_PHN4201_n5643));
   CLKBUF_X1 FE_PHC5001_n5376 (.Z(FE_PHN5001_n5376), 
	.A(FE_PHN4141_n5376));
   CLKBUF_X1 FE_PHC5000_n5508 (.Z(FE_PHN5000_n5508), 
	.A(FE_PHN4078_n5508));
   BUF_X2 FE_PHC4999_U320_Z_0 (.Z(FE_PHN4999_U320_Z_0), 
	.A(FE_PHN2210_U320_Z_0));
   BUF_X1 FE_PHC4997_n5490 (.Z(FE_PHN4997_n5490), 
	.A(FE_PHN3972_n5490));
   BUF_X1 FE_PHC4995_n5109 (.Z(FE_PHN4995_n5109), 
	.A(FE_PHN4102_n5109));
   CLKBUF_X2 FE_PHC4994_n5336 (.Z(FE_PHN4994_n5336), 
	.A(FE_PHN4043_n5336));
   BUF_X1 FE_PHC4991_U234_Z_0 (.Z(FE_PHN4991_U234_Z_0), 
	.A(FE_PHN3877_U234_Z_0));
   CLKBUF_X1 FE_PHC4990_n5092 (.Z(FE_PHN4990_n5092), 
	.A(FE_PHN3969_n5092));
   CLKBUF_X1 FE_PHC4989_n5496 (.Z(FE_PHN4989_n5496), 
	.A(FE_PHN4088_n5496));
   CLKBUF_X1 FE_PHC4988_n5218 (.Z(FE_PHN4988_n5218), 
	.A(FE_PHN4160_n5218));
   CLKBUF_X1 FE_PHC4986_U800_Z_0 (.Z(FE_PHN4986_U800_Z_0), 
	.A(FE_PHN3845_U800_Z_0));
   CLKBUF_X1 FE_PHC4985_n5792 (.Z(FE_PHN4985_n5792), 
	.A(FE_PHN2415_n5792));
   CLKBUF_X1 FE_PHC4984_U305_Z_0 (.Z(FE_PHN4984_U305_Z_0), 
	.A(FE_PHN2066_U305_Z_0));
   CLKBUF_X1 FE_PHC4983_U557_Z_0 (.Z(FE_PHN4983_U557_Z_0), 
	.A(FE_PHN2074_U557_Z_0));
   CLKBUF_X1 FE_PHC4982_U606_Z_0 (.Z(FE_PHN4982_U606_Z_0), 
	.A(FE_PHN4034_U606_Z_0));
   CLKBUF_X1 FE_PHC4980_n5283 (.Z(FE_PHN4980_n5283), 
	.A(FE_PHN3961_n5283));
   CLKBUF_X1 FE_PHC4977_n5353 (.Z(FE_PHN4977_n5353), 
	.A(FE_PHN3958_n5353));
   CLKBUF_X1 FE_PHC4976_n5599 (.Z(FE_PHN4976_n5599), 
	.A(FE_PHN4108_n5599));
   BUF_X1 FE_PHC4974_n5634 (.Z(FE_PHN4974_n5634), 
	.A(FE_PHN3962_n5634));
   BUF_X1 FE_PHC4972_n5261 (.Z(FE_PHN4972_n5261), 
	.A(FE_PHN4169_n5261));
   BUF_X1 FE_PHC4971_n5380 (.Z(FE_PHN4971_n5380), 
	.A(FE_PHN3915_n5380));
   BUF_X1 FE_PHC4970_n5365 (.Z(FE_PHN4970_n5365), 
	.A(FE_PHN4142_n5365));
   CLKBUF_X2 FE_PHC4969_n5198 (.Z(FE_PHN4969_n5198), 
	.A(FE_PHN3948_n5198));
   BUF_X1 FE_PHC4967_n5394 (.Z(FE_PHN4967_n5394), 
	.A(FE_PHN4176_n5394));
   CLKBUF_X1 FE_PHC4963_n5356 (.Z(FE_PHN4963_n5356), 
	.A(FE_PHN4124_n5356));
   BUF_X2 FE_PHC4960_U324_Z_0 (.Z(FE_PHN4960_U324_Z_0), 
	.A(FE_PHN2072_U324_Z_0));
   CLKBUF_X1 FE_PHC4959_n5350 (.Z(FE_PHN4959_n5350), 
	.A(FE_PHN4022_n5350));
   CLKBUF_X1 FE_PHC4958_U411_Z_0 (.Z(FE_PHN4958_U411_Z_0), 
	.A(FE_PHN4024_U411_Z_0));
   CLKBUF_X1 FE_PHC4956_n5073 (.Z(FE_PHN4956_n5073), 
	.A(FE_PHN3916_n5073));
   CLKBUF_X1 FE_PHC4955_n5214 (.Z(FE_PHN4955_n5214), 
	.A(FE_PHN4041_n5214));
   CLKBUF_X1 FE_PHC4954_U471_Z_0 (.Z(FE_PHN4954_U471_Z_0), 
	.A(FE_PHN3847_U471_Z_0));
   CLKBUF_X1 FE_PHC4953_n5066 (.Z(FE_PHN4953_n5066), 
	.A(FE_PHN3872_n5066));
   CLKBUF_X1 FE_PHC4950_n5403 (.Z(FE_PHN4950_n5403), 
	.A(FE_PHN4120_n5403));
   BUF_X1 FE_PHC4949_n5515 (.Z(FE_PHN4949_n5515), 
	.A(FE_PHN3928_n5515));
   CLKBUF_X2 FE_PHC4947_n5357 (.Z(FE_PHN4947_n5357), 
	.A(FE_PHN4146_n5357));
   BUF_X1 FE_PHC4946_n5372 (.Z(FE_PHN4946_n5372), 
	.A(FE_PHN4042_n5372));
   BUF_X2 FE_PHC4944_U323_Z_0 (.Z(FE_PHN4944_U323_Z_0), 
	.A(FE_PHN2056_U323_Z_0));
   CLKBUF_X1 FE_PHC4943_U566_Z_0 (.Z(FE_PHN4943_U566_Z_0), 
	.A(FE_PHN1742_U566_Z_0));
   CLKBUF_X1 FE_PHC4941_n5275 (.Z(FE_PHN4941_n5275), 
	.A(FE_PHN3930_n5275));
   CLKBUF_X1 FE_PHC4940_n5379 (.Z(FE_PHN4940_n5379), 
	.A(FE_PHN4017_n5379));
   CLKBUF_X1 FE_PHC4937_n5788 (.Z(FE_PHN4937_n5788), 
	.A(FE_PHN1450_n5788));
   CLKBUF_X1 FE_PHC4935_n5390 (.Z(FE_PHN4935_n5390), 
	.A(FE_PHN3875_n5390));
   CLKBUF_X1 FE_PHC4933_n5226 (.Z(FE_PHN4933_n5226), 
	.A(FE_PHN3917_n5226));
   CLKBUF_X1 FE_PHC4932_U506_Z_0 (.Z(FE_PHN4932_U506_Z_0), 
	.A(FE_PHN4096_U506_Z_0));
   CLKBUF_X1 FE_PHC4931_n5273 (.Z(FE_PHN4931_n5273), 
	.A(FE_PHN4177_n5273));
   CLKBUF_X1 FE_PHC4930_U563_Z_0 (.Z(FE_PHN4930_U563_Z_0), 
	.A(FE_PHN2059_U563_Z_0));
   BUF_X2 FE_PHC4927_U395_Z_0 (.Z(FE_PHN4927_U395_Z_0), 
	.A(FE_PHN3976_U395_Z_0));
   BUF_X1 FE_PHC4924_n5286 (.Z(FE_PHN4924_n5286), 
	.A(FE_PHN4051_n5286));
   BUF_X2 FE_PHC4923_U318_Z_0 (.Z(FE_PHN4923_U318_Z_0), 
	.A(FE_PHN2060_U318_Z_0));
   CLKBUF_X1 FE_PHC4921_U673_Z_0 (.Z(FE_PHN4921_U673_Z_0), 
	.A(FE_PHN4023_U673_Z_0));
   CLKBUF_X1 FE_PHC4920_U726_Z_0 (.Z(FE_PHN4920_U726_Z_0), 
	.A(FE_PHN4048_U726_Z_0));
   CLKBUF_X1 FE_PHC4919_n5494 (.Z(FE_PHN4919_n5494), 
	.A(FE_PHN3907_n5494));
   CLKBUF_X1 FE_PHC4916_n5738 (.Z(FE_PHN4916_n5738), 
	.A(FE_PHN1472_n5738));
   BUF_X1 FE_PHC4912_n5335 (.Z(FE_PHN4912_n5335), 
	.A(FE_PHN4115_n5335));
   BUF_X1 FE_PHC4911_n5210 (.Z(FE_PHN4911_n5210), 
	.A(FE_PHN3892_n5210));
   BUF_X1 FE_PHC4910_n5497 (.Z(FE_PHN4910_n5497), 
	.A(FE_PHN3986_n5497));
   BUF_X1 FE_PHC4909_n5277 (.Z(FE_PHN4909_n5277), 
	.A(FE_PHN4118_n5277));
   CLKBUF_X1 FE_PHC4907_U619_Z_0 (.Z(FE_PHN4907_U619_Z_0), 
	.A(FE_PHN3843_U619_Z_0));
   CLKBUF_X1 FE_PHC4906_n5541 (.Z(FE_PHN4906_n5541), 
	.A(FE_PHN4020_n5541));
   CLKBUF_X1 FE_PHC4905_U692_Z_0 (.Z(FE_PHN4905_U692_Z_0), 
	.A(FE_PHN3076_U692_Z_0));
   CLKBUF_X1 FE_PHC4904_n5374 (.Z(FE_PHN4904_n5374), 
	.A(FE_PHN4085_n5374));
   CLKBUF_X1 FE_PHC4902_n5479 (.Z(FE_PHN4902_n5479), 
	.A(FE_PHN4084_n5479));
   CLKBUF_X1 FE_PHC4900_U263_Z_0 (.Z(FE_PHN4900_U263_Z_0), 
	.A(FE_PHN3842_U263_Z_0));
   BUF_X1 FE_PHC4898_n5495 (.Z(FE_PHN4898_n5495), 
	.A(FE_PHN3977_n5495));
   CLKBUF_X1 FE_PHC4897_U513_Z_0 (.Z(FE_PHN4897_U513_Z_0), 
	.A(FE_PHN3811_U513_Z_0));
   BUF_X1 FE_PHC4896_n5134 (.Z(FE_PHN4896_n5134), 
	.A(FE_PHN3780_n5134));
   CLKBUF_X1 FE_PHC4895_U745_Z_0 (.Z(FE_PHN4895_U745_Z_0), 
	.A(FE_PHN3839_U745_Z_0));
   CLKBUF_X1 FE_PHC4891_U663_Z_0 (.Z(FE_PHN4891_U663_Z_0), 
	.A(FE_PHN3806_U663_Z_0));
   CLKBUF_X1 FE_PHC4890_U481_Z_0 (.Z(FE_PHN4890_U481_Z_0), 
	.A(FE_PHN3821_U481_Z_0));
   CLKBUF_X1 FE_PHC4888_n4998 (.Z(FE_PHN4888_n4998), 
	.A(FE_PHN4005_n4998));
   CLKBUF_X1 FE_PHC4887_n5341 (.Z(FE_PHN4887_n5341), 
	.A(FE_PHN3893_n5341));
   CLKBUF_X1 FE_PHC4886_n5216 (.Z(FE_PHN4886_n5216), 
	.A(FE_PHN3987_n5216));
   CLKBUF_X1 FE_PHC4885_n5559 (.Z(FE_PHN4885_n5559), 
	.A(FE_PHN3981_n5559));
   CLKBUF_X1 FE_PHC4884_U504_Z_0 (.Z(FE_PHN4884_U504_Z_0), 
	.A(FE_PHN3851_U504_Z_0));
   CLKBUF_X1 FE_PHC4883_n5354 (.Z(FE_PHN4883_n5354), 
	.A(FE_PHN3884_n5354));
   BUF_X1 FE_PHC4882_U660_Z_0 (.Z(FE_PHN4882_U660_Z_0), 
	.A(FE_PHN4053_U660_Z_0));
   CLKBUF_X1 FE_PHC4876_n5480 (.Z(FE_PHN4876_n5480), 
	.A(FE_PHN4077_n5480));
   CLKBUF_X1 FE_PHC4874_n5630 (.Z(FE_PHN4874_n5630), 
	.A(FE_PHN4061_n5630));
   CLKBUF_X1 FE_PHC4873_n5566 (.Z(FE_PHN4873_n5566), 
	.A(FE_PHN4018_n5566));
   CLKBUF_X1 FE_PHC4870_n5334 (.Z(FE_PHN4870_n5334), 
	.A(FE_PHN4082_n5334));
   CLKBUF_X1 FE_PHC4869_U475_Z_0 (.Z(FE_PHN4869_U475_Z_0), 
	.A(FE_PHN4054_U475_Z_0));
   BUF_X1 FE_PHC4868_n5608 (.Z(FE_PHN4868_n5608), 
	.A(FE_PHN3959_n5608));
   BUF_X1 FE_PHC4867_n5506 (.Z(FE_PHN4867_n5506), 
	.A(FE_PHN3871_n5506));
   BUF_X1 FE_PHC4866_n5037 (.Z(FE_PHN4866_n5037), 
	.A(FE_PHN3970_n5037));
   CLKBUF_X1 FE_PHC4865_U500_Z_0 (.Z(FE_PHN4865_U500_Z_0), 
	.A(FE_PHN3775_U500_Z_0));
   CLKBUF_X1 FE_PHC4864_U585_Z_0 (.Z(FE_PHN4864_U585_Z_0), 
	.A(FE_PHN3823_U585_Z_0));
   CLKBUF_X1 FE_PHC4863_U466_Z_0 (.Z(FE_PHN4863_U466_Z_0), 
	.A(FE_PHN3882_U466_Z_0));
   BUF_X2 FE_PHC4862_U291_Z_0 (.Z(FE_PHN4862_U291_Z_0), 
	.A(FE_PHN3971_U291_Z_0));
   CLKBUF_X1 FE_PHC4861_n5278 (.Z(FE_PHN4861_n5278), 
	.A(FE_PHN4060_n5278));
   CLKBUF_X1 FE_PHC4860_U779_Z_0 (.Z(FE_PHN4860_U779_Z_0), 
	.A(FE_PHN4035_U779_Z_0));
   CLKBUF_X1 FE_PHC4859_n5563 (.Z(FE_PHN4859_n5563), 
	.A(FE_PHN3942_n5563));
   CLKBUF_X1 FE_PHC4857_U667_Z_0 (.Z(FE_PHN4857_U667_Z_0), 
	.A(FE_PHN3785_U667_Z_0));
   CLKBUF_X1 FE_PHC4854_n5276 (.Z(FE_PHN4854_n5276), 
	.A(FE_PHN3911_n5276));
   CLKBUF_X1 FE_PHC4853_n5063 (.Z(FE_PHN4853_n5063), 
	.A(FE_PHN4003_n5063));
   CLKBUF_X1 FE_PHC4850_n5168 (.Z(FE_PHN4850_n5168), 
	.A(FE_PHN3828_n5168));
   BUF_X1 FE_PHC4847_n5382 (.Z(FE_PHN4847_n5382), 
	.A(FE_PHN3949_n5382));
   CLKBUF_X1 FE_PHC4844_U712_Z_0 (.Z(FE_PHN4844_U712_Z_0), 
	.A(FE_PHN3887_U712_Z_0));
   CLKBUF_X1 FE_PHC4840_n5577 (.Z(FE_PHN4840_n5577), 
	.A(FE_PHN3985_n5577));
   CLKBUF_X1 FE_PHC4839_n5569 (.Z(FE_PHN4839_n5569), 
	.A(FE_PHN3954_n5569));
   CLKBUF_X1 FE_PHC4838_n5131 (.Z(FE_PHN4838_n5131), 
	.A(FE_PHN3937_n5131));
   CLKBUF_X1 FE_PHC4835_U454_Z_0 (.Z(FE_PHN4835_U454_Z_0), 
	.A(FE_PHN3798_U454_Z_0));
   CLKBUF_X1 FE_PHC4834_U743_Z_0 (.Z(FE_PHN4834_U743_Z_0), 
	.A(FE_PHN3778_U743_Z_0));
   CLKBUF_X1 FE_PHC4833_n5343 (.Z(FE_PHN4833_n5343), 
	.A(FE_PHN4027_n5343));
   CLKBUF_X1 FE_PHC4831_n4982 (.Z(FE_PHN4831_n4982), 
	.A(FE_PHN3793_n4982));
   CLKBUF_X1 FE_PHC4830_U748_Z_0 (.Z(FE_PHN4830_U748_Z_0), 
	.A(FE_PHN3803_U748_Z_0));
   CLKBUF_X1 FE_PHC4829_n5791 (.Z(FE_PHN4829_n5791), 
	.A(FE_PHN3209_n5791));
   CLKBUF_X1 FE_PHC4828_n5574 (.Z(FE_PHN4828_n5574), 
	.A(FE_PHN3926_n5574));
   CLKBUF_X1 FE_PHC4827_n5087 (.Z(FE_PHN4827_n5087), 
	.A(FE_PHN4001_n5087));
   BUF_X1 FE_PHC4823_n5631 (.Z(FE_PHN4823_n5631), 
	.A(FE_PHN3960_n5631));
   CLKBUF_X1 FE_PHC4822_n5389 (.Z(FE_PHN4822_n5389), 
	.A(FE_PHN3898_n5389));
   CLKBUF_X1 FE_PHC4821_n5607 (.Z(FE_PHN4821_n5607), 
	.A(FE_PHN3924_n5607));
   CLKBUF_X1 FE_PHC4820_U242_Z_0 (.Z(FE_PHN4820_U242_Z_0), 
	.A(FE_PHN3787_U242_Z_0));
   CLKBUF_X1 FE_PHC4815_U651_Z_0 (.Z(FE_PHN4815_U651_Z_0), 
	.A(FE_PHN3784_U651_Z_0));
   CLKBUF_X1 FE_PHC4814_U445_Z_0 (.Z(FE_PHN4814_U445_Z_0), 
	.A(FE_PHN3753_U445_Z_0));
   CLKBUF_X1 FE_PHC4813_n5683 (.Z(FE_PHN4813_n5683), 
	.A(FE_PHN936_n5683));
   CLKBUF_X1 FE_PHC4810_U708_Z_0 (.Z(FE_PHN4810_U708_Z_0), 
	.A(FE_PHN3774_U708_Z_0));
   CLKBUF_X1 FE_PHC4809_n5264 (.Z(FE_PHN4809_n5264), 
	.A(FE_PHN3918_n5264));
   CLKBUF_X1 FE_PHC4808_n5345 (.Z(FE_PHN4808_n5345), 
	.A(FE_PHN3896_n5345));
   CLKBUF_X1 FE_PHC4807_n5340 (.Z(FE_PHN4807_n5340), 
	.A(FE_PHN3879_n5340));
   CLKBUF_X1 FE_PHC4804_n14928 (.Z(FE_PHN4804_n14928), 
	.A(FE_PHN892_n14928));
   CLKBUF_X1 FE_PHC4802_n5263 (.Z(FE_PHN4802_n5263), 
	.A(FE_PHN3983_n5263));
   CLKBUF_X1 FE_PHC4801_n5543 (.Z(FE_PHN4801_n5543), 
	.A(FE_PHN3908_n5543));
   BUF_X1 FE_PHC4797_U325_Z_0 (.Z(FE_PHN4797_U325_Z_0), 
	.A(FE_PHN3950_U325_Z_0));
   CLKBUF_X1 FE_PHC4796_n5122 (.Z(FE_PHN4796_n5122), 
	.A(FE_PHN3919_n5122));
   CLKBUF_X1 FE_PHC4795_n5368 (.Z(FE_PHN4795_n5368), 
	.A(FE_PHN3931_n5368));
   CLKBUF_X1 FE_PHC4794_n5215 (.Z(FE_PHN4794_n5215), 
	.A(FE_PHN3909_n5215));
   CLKBUF_X1 FE_PHC4790_n5125 (.Z(FE_PHN4790_n5125), 
	.A(FE_PHN3963_n5125));
   CLKBUF_X1 FE_PHC4788_U496_Z_0 (.Z(FE_PHN4788_U496_Z_0), 
	.A(FE_PHN3762_U496_Z_0));
   CLKBUF_X1 FE_PHC4784_n5627 (.Z(FE_PHN4784_n5627), 
	.A(FE_PHN3922_n5627));
   CLKBUF_X1 FE_PHC4783_n4938 (.Z(FE_PHN4783_n4938), 
	.A(FE_PHN1978_n4938));
   CLKBUF_X1 FE_PHC4782_n5548 (.Z(FE_PHN4782_n5548), 
	.A(FE_PHN3941_n5548));
   CLKBUF_X1 FE_PHC4781_U728_Z_0 (.Z(FE_PHN4781_U728_Z_0), 
	.A(FE_PHN3782_U728_Z_0));
   CLKBUF_X1 FE_PHC4779_n4937 (.Z(FE_PHN4779_n4937), 
	.A(FE_PHN1910_n4937));
   CLKBUF_X1 FE_PHC4778_n5614 (.Z(FE_PHN4778_n5614), 
	.A(FE_PHN3888_n5614));
   CLKBUF_X1 FE_PHC4774_U683_Z_0 (.Z(FE_PHN4774_U683_Z_0), 
	.A(FE_PHN3765_U683_Z_0));
   CLKBUF_X1 FE_PHC4772_U628_Z_0 (.Z(FE_PHN4772_U628_Z_0), 
	.A(FE_PHN3853_U628_Z_0));
   CLKBUF_X1 FE_PHC4767_n5265 (.Z(FE_PHN4767_n5265), 
	.A(FE_PHN3866_n5265));
   CLKBUF_X1 FE_PHC4761_U634_Z_0 (.Z(FE_PHN4761_U634_Z_0), 
	.A(FE_PHN3682_U634_Z_0));
   CLKBUF_X1 FE_PHC4756_n5056 (.Z(FE_PHN4756_n5056), 
	.A(FE_PHN3699_n5056));
   CLKBUF_X1 FE_PHC4750_n5565 (.Z(FE_PHN4750_n5565), 
	.A(n5565));
   CLKBUF_X1 FE_PHC4749_n4925 (.Z(FE_PHN4749_n4925), 
	.A(FE_PHN1908_n4925));
   CLKBUF_X1 FE_PHC4748_n276 (.Z(FE_PHN4748_n276), 
	.A(FE_PHN3662_n276));
   CLKBUF_X1 FE_PHC4743_U656_Z_0 (.Z(FE_PHN4743_U656_Z_0), 
	.A(FE_PHN3663_U656_Z_0));
   CLKBUF_X1 FE_PHC4739_n5586 (.Z(FE_PHN4739_n5586), 
	.A(FE_PHN3617_n5586));
   CLKBUF_X1 FE_PHC4737_n5712 (.Z(FE_PHN4737_n5712), 
	.A(FE_PHN1919_n5712));
   CLKBUF_X1 FE_PHC4735_n4939 (.Z(FE_PHN4735_n4939), 
	.A(FE_PHN1174_n4939));
   CLKBUF_X1 FE_PHC4734_n5555 (.Z(FE_PHN4734_n5555), 
	.A(n5555));
   CLKBUF_X1 FE_PHC4733_n4935 (.Z(FE_PHN4733_n4935), 
	.A(FE_PHN1920_n4935));
   CLKBUF_X1 FE_PHC4732_n5561 (.Z(FE_PHN4732_n5561), 
	.A(n5561));
   CLKBUF_X1 FE_PHC4731_n4936 (.Z(FE_PHN4731_n4936), 
	.A(FE_PHN1915_n4936));
   CLKBUF_X1 FE_PHC4730_n4926 (.Z(FE_PHN4730_n4926), 
	.A(FE_PHN1912_n4926));
   CLKBUF_X1 FE_PHC4729_n4942 (.Z(FE_PHN4729_n4942), 
	.A(FE_PHN1914_n4942));
   BUF_X32 FE_PHC4726_n5760 (.Z(FE_PHN4726_n5760), 
	.A(FE_PHN5233_n5760));
   BUF_X32 FE_PHC4725_n385 (.Z(FE_PHN4725_n385), 
	.A(FE_PHN5232_n385));
   BUF_X32 FE_PHC4724_n1136 (.Z(FE_PHN4724_n1136), 
	.A(FE_PHN5231_n1136));
   BUF_X32 FE_PHC4723_n419 (.Z(FE_PHN4723_n419), 
	.A(FE_PHN5230_n419));
   BUF_X32 FE_PHC4722_n1135 (.Z(FE_PHN4722_n1135), 
	.A(FE_PHN5229_n1135));
   BUF_X32 FE_PHC4721_n1141 (.Z(FE_PHN4721_n1141), 
	.A(FE_PHN5228_n1141));
   BUF_X32 FE_PHC4720_n1138 (.Z(FE_PHN4720_n1138), 
	.A(FE_PHN5227_n1138));
   CLKBUF_X1 FE_PHC4712_n4923 (.Z(FE_PHN4712_n4923), 
	.A(FE_PHN3290_n4923));
   BUF_X32 FE_PHC4711_U227_Z_0 (.Z(FE_PHN4711_U227_Z_0), 
	.A(FE_PHN5226_U227_Z_0));
   BUF_X32 FE_PHC4710_n5751 (.Z(FE_PHN4710_n5751), 
	.A(FE_PHN5224_n5751));
   BUF_X32 FE_PHC4709_n5752 (.Z(FE_PHN4709_n5752), 
	.A(FE_PHN5223_n5752));
   BUF_X32 FE_PHC4708_n5746 (.Z(FE_PHN4708_n5746), 
	.A(FE_PHN5225_n5746));
   BUF_X32 FE_PHC4707_n5750 (.Z(FE_PHN4707_n5750), 
	.A(FE_PHN5222_n5750));
   BUF_X32 FE_PHC4706_n5763 (.Z(FE_PHN4706_n5763), 
	.A(FE_PHN5221_n5763));
   BUF_X32 FE_PHC4704_n5754 (.Z(FE_PHN4704_n5754), 
	.A(FE_PHN5220_n5754));
   BUF_X32 FE_PHC4703_n5756 (.Z(FE_PHN4703_n5756), 
	.A(FE_PHN5219_n5756));
   BUF_X32 FE_PHC4702_n1146 (.Z(FE_PHN4702_n1146), 
	.A(FE_PHN5216_n1146));
   BUF_X32 FE_PHC4701_n380 (.Z(FE_PHN4701_n380), 
	.A(FE_PHN5217_n380));
   BUF_X32 FE_PHC4700_n387 (.Z(FE_PHN4700_n387), 
	.A(FE_PHN5215_n387));
   BUF_X32 FE_PHC4699_n1132 (.Z(FE_PHN4699_n1132), 
	.A(FE_PHN5213_n1132));
   BUF_X32 FE_PHC4698_n1133 (.Z(FE_PHN4698_n1133), 
	.A(FE_PHN5214_n1133));
   BUF_X32 FE_PHC4697_n1130 (.Z(FE_PHN4697_n1130), 
	.A(FE_PHN5212_n1130));
   BUF_X32 FE_PHC4696_n1139 (.Z(FE_PHN4696_n1139), 
	.A(FE_PHN5211_n1139));
   BUF_X32 FE_PHC4695_n395 (.Z(FE_PHN4695_n395), 
	.A(FE_PHN5210_n395));
   BUF_X32 FE_PHC4694_n14432 (.Z(FE_PHN4694_n14432), 
	.A(FE_PHN5209_n14432));
   BUF_X32 FE_PHC4693_n389 (.Z(FE_PHN4693_n389), 
	.A(FE_PHN5208_n389));
   BUF_X32 FE_PHC4692_n4917 (.Z(FE_PHN4692_n4917), 
	.A(n4917));
   BUF_X32 FE_PHC4691_n4919 (.Z(FE_PHN4691_n4919), 
	.A(n4919));
   BUF_X32 FE_PHC4690_n4918 (.Z(FE_PHN4690_n4918), 
	.A(n4918));
   BUF_X32 FE_PHC4689_n5761 (.Z(FE_PHN4689_n5761), 
	.A(FE_PHN5205_n5761));
   BUF_X32 FE_PHC4688_n4915 (.Z(FE_PHN4688_n4915), 
	.A(FE_PHN5244_n4915));
   BUF_X32 FE_PHC4687_n5741 (.Z(FE_PHN4687_n5741), 
	.A(FE_PHN5202_n5741));
   BUF_X32 FE_PHC4686_n5744 (.Z(FE_PHN4686_n5744), 
	.A(FE_PHN5201_n5744));
   BUF_X32 FE_PHC4685_n5753 (.Z(FE_PHN4685_n5753), 
	.A(FE_PHN5200_n5753));
   BUF_X32 FE_PHC4684_n5766 (.Z(FE_PHN4684_n5766), 
	.A(FE_PHN5199_n5766));
   BUF_X32 FE_PHC4683_n5739 (.Z(FE_PHN4683_n5739), 
	.A(FE_PHN5198_n5739));
   BUF_X32 FE_PHC4682_n5765 (.Z(FE_PHN4682_n5765), 
	.A(FE_PHN5197_n5765));
   BUF_X32 FE_PHC4681_n5745 (.Z(FE_PHN4681_n5745), 
	.A(FE_PHN5196_n5745));
   BUF_X32 FE_PHC4680_n5749 (.Z(FE_PHN4680_n5749), 
	.A(FE_PHN5195_n5749));
   BUF_X32 FE_PHC4679_n5742 (.Z(FE_PHN4679_n5742), 
	.A(FE_PHN5194_n5742));
   CLKBUF_X1 FE_PHC4675_n4902 (.Z(FE_PHN4675_n4902), 
	.A(n4902));
   BUF_X16 FE_PHC4674_n4394 (.Z(FE_PHN4674_n4394), 
	.A(n4394));
   BUF_X16 FE_PHC4673_n4389 (.Z(FE_PHN4673_n4389), 
	.A(n4389));
   BUF_X32 FE_PHC4672_n4300 (.Z(FE_PHN4672_n4300), 
	.A(n4300));
   BUF_X32 FE_PHC4671_n4903 (.Z(FE_PHN4671_n4903), 
	.A(n4903));
   BUF_X32 FE_PHC4670_n4193 (.Z(FE_PHN4670_n4193), 
	.A(n4193));
   BUF_X32 FE_PHC4669_n4324 (.Z(FE_PHN4669_n4324), 
	.A(n4324));
   BUF_X32 FE_PHC4668_n4391 (.Z(FE_PHN4668_n4391), 
	.A(n4391));
   BUF_X32 FE_PHC4667_n4397 (.Z(FE_PHN4667_n4397), 
	.A(n4397));
   BUF_X32 FE_PHC4666_n4190 (.Z(FE_PHN4666_n4190), 
	.A(n4190));
   BUF_X32 FE_PHC4662_n5768 (.Z(FE_PHN4662_n5768), 
	.A(FE_PHN5188_n5768));
   BUF_X32 FE_PHC4661_n5767 (.Z(FE_PHN4661_n5767), 
	.A(FE_PHN5187_n5767));
   BUF_X32 FE_PHC4660_n5769 (.Z(FE_PHN4660_n5769), 
	.A(FE_PHN5186_n5769));
   BUF_X32 FE_PHC4659_n5743 (.Z(FE_PHN4659_n5743), 
	.A(FE_PHN5185_n5743));
   BUF_X32 FE_PHC4658_n5747 (.Z(FE_PHN4658_n5747), 
	.A(FE_PHN5183_n5747));
   BUF_X32 FE_PHC4657_n5748 (.Z(FE_PHN4657_n5748), 
	.A(FE_PHN5184_n5748));
   BUF_X32 FE_PHC4656_n5740 (.Z(FE_PHN4656_n5740), 
	.A(FE_PHN5182_n5740));
   BUF_X32 FE_PHC4655_n4909 (.Z(FE_PHN4655_n4909), 
	.A(FE_PHN819_n4909));
   BUF_X32 FE_PHC4654_n4912 (.Z(FE_PHN4654_n4912), 
	.A(FE_PHN818_n4912));
   CLKBUF_X1 FE_PHC4653_n3273 (.Z(FE_PHN4653_n3273), 
	.A(n3273));
   BUF_X16 FE_PHC4652_n4920 (.Z(FE_PHN4652_n4920), 
	.A(n4920));
   BUF_X16 FE_PHC4641_IRQ_14_ (.Z(FE_PHN4641_IRQ_14_), 
	.A(FE_PHN3018_IRQ_14_));
   CLKBUF_X1 FE_PHC4639_n5692 (.Z(FE_PHN4639_n5692), 
	.A(FE_PHN2927_n5692));
   BUF_X16 FE_PHC4638_IRQ_11_ (.Z(FE_PHN4638_IRQ_11_), 
	.A(FE_PHN2994_IRQ_11_));
   BUF_X32 FE_PHC4637_IRQ_9_ (.Z(FE_PHN4637_IRQ_9_), 
	.A(FE_PHN2988_IRQ_9_));
   BUF_X32 FE_PHC4634_IRQ_1_ (.Z(FE_PHN4634_IRQ_1_), 
	.A(FE_PHN2983_IRQ_1_));
   CLKBUF_X1 FE_PHC4631_NMI (.Z(FE_PHN4631_NMI), 
	.A(FE_PHN2982_NMI));
   CLKBUF_X1 FE_PHC4630_IRQ_15_ (.Z(FE_PHN4630_IRQ_15_), 
	.A(FE_PHN2980_IRQ_15_));
   BUF_X32 FE_PHC4629_n17127 (.Z(FE_PHN4629_n17127), 
	.A(FE_PHN2912_n17127));
   BUF_X32 FE_PHC4624_n17126 (.Z(FE_PHN4624_n17126), 
	.A(FE_PHN5192_n17126));
   CLKBUF_X1 FE_PHC4615_U762_Z_0 (.Z(FE_PHN4615_U762_Z_0), 
	.A(U762_Z_0));
   CLKBUF_X1 FE_PHC4611_n5710 (.Z(FE_PHN4611_n5710), 
	.A(FE_PHN2898_n5710));
   CLKBUF_X1 FE_PHC4608_U802_Z_0 (.Z(FE_PHN4608_U802_Z_0), 
	.A(U802_Z_0));
   CLKBUF_X1 FE_PHC4607_n5652 (.Z(FE_PHN4607_n5652), 
	.A(n5652));
   CLKBUF_X1 FE_PHC4602_n4890 (.Z(FE_PHN4602_n4890), 
	.A(n4890));
   CLKBUF_X1 FE_PHC4601_U317_Z_0 (.Z(FE_PHN4601_U317_Z_0), 
	.A(FE_PHN1898_U317_Z_0));
   CLKBUF_X1 FE_PHC4597_U789_Z_0 (.Z(FE_PHN4597_U789_Z_0), 
	.A(U789_Z_0));
   CLKBUF_X1 FE_PHC4596_U781_Z_0 (.Z(FE_PHN4596_U781_Z_0), 
	.A(U781_Z_0));
   CLKBUF_X1 FE_PHC4595_U791_Z_0 (.Z(FE_PHN4595_U791_Z_0), 
	.A(FE_PHN2890_U791_Z_0));
   CLKBUF_X1 FE_PHC4590_U518_Z_0 (.Z(FE_PHN4590_U518_Z_0), 
	.A(U518_Z_0));
   CLKBUF_X1 FE_PHC4588_n5704 (.Z(FE_PHN4588_n5704), 
	.A(n5704));
   CLKBUF_X1 FE_PHC4586_n5097 (.Z(FE_PHN4586_n5097), 
	.A(n5097));
   CLKBUF_X1 FE_PHC4585_n5706 (.Z(FE_PHN4585_n5706), 
	.A(FE_PHN2901_n5706));
   CLKBUF_X1 FE_PHC4584_n5737 (.Z(FE_PHN4584_n5737), 
	.A(FE_PHN1588_n5737));
   CLKBUF_X1 FE_PHC4583_n5651 (.Z(FE_PHN4583_n5651), 
	.A(n5651));
   CLKBUF_X1 FE_PHC4580_U763_Z_0 (.Z(FE_PHN4580_U763_Z_0), 
	.A(FE_PHN2897_U763_Z_0));
   CLKBUF_X1 FE_PHC4579_n5705 (.Z(FE_PHN4579_n5705), 
	.A(n5705));
   CLKBUF_X1 FE_PHC4577_n5612 (.Z(FE_PHN4577_n5612), 
	.A(n5612));
   CLKBUF_X1 FE_PHC4576_U782_Z_0 (.Z(FE_PHN4576_U782_Z_0), 
	.A(U782_Z_0));
   CLKBUF_X1 FE_PHC4575_n4862 (.Z(FE_PHN4575_n4862), 
	.A(n4862));
   CLKBUF_X1 FE_PHC4573_n5130 (.Z(FE_PHN4573_n5130), 
	.A(n5130));
   CLKBUF_X1 FE_PHC4572_U783_Z_0 (.Z(FE_PHN4572_U783_Z_0), 
	.A(U783_Z_0));
   CLKBUF_X1 FE_PHC4571_U144_Z_0 (.Z(FE_PHN4571_U144_Z_0), 
	.A(FE_PHN2039_U144_Z_0));
   CLKBUF_X1 FE_PHC4570_n5568 (.Z(FE_PHN4570_n5568), 
	.A(n5568));
   CLKBUF_X1 FE_PHC4569_n5103 (.Z(FE_PHN4569_n5103), 
	.A(n5103));
   CLKBUF_X1 FE_PHC4567_n5172 (.Z(FE_PHN4567_n5172), 
	.A(n5172));
   CLKBUF_X1 FE_PHC4566_U771_Z_0 (.Z(FE_PHN4566_U771_Z_0), 
	.A(U771_Z_0));
   CLKBUF_X1 FE_PHC4565_n5015 (.Z(FE_PHN4565_n5015), 
	.A(n5015));
   CLKBUF_X1 FE_PHC4564_n5012 (.Z(FE_PHN4564_n5012), 
	.A(n5012));
   CLKBUF_X1 FE_PHC4563_n5450 (.Z(FE_PHN4563_n5450), 
	.A(n5450));
   CLKBUF_X1 FE_PHC4562_n5702 (.Z(FE_PHN4562_n5702), 
	.A(FE_PHN2900_n5702));
   CLKBUF_X1 FE_PHC4561_n4857 (.Z(FE_PHN4561_n4857), 
	.A(n4857));
   CLKBUF_X1 FE_PHC4560_n5267 (.Z(FE_PHN4560_n5267), 
	.A(n5267));
   CLKBUF_X1 FE_PHC4559_n5457 (.Z(FE_PHN4559_n5457), 
	.A(n5457));
   CLKBUF_X1 FE_PHC4557_n5299 (.Z(FE_PHN4557_n5299), 
	.A(n5299));
   CLKBUF_X1 FE_PHC4556_n5396 (.Z(FE_PHN4556_n5396), 
	.A(n5396));
   CLKBUF_X1 FE_PHC4555_U772_Z_0 (.Z(FE_PHN4555_U772_Z_0), 
	.A(U772_Z_0));
   CLKBUF_X1 FE_PHC4554_n5178 (.Z(FE_PHN4554_n5178), 
	.A(n5178));
   CLKBUF_X1 FE_PHC4553_n5604 (.Z(FE_PHN4553_n5604), 
	.A(n5604));
   CLKBUF_X1 FE_PHC4552_n4885 (.Z(FE_PHN4552_n4885), 
	.A(n4885));
   CLKBUF_X1 FE_PHC4550_n4856 (.Z(FE_PHN4550_n4856), 
	.A(n4856));
   CLKBUF_X1 FE_PHC4549_n5284 (.Z(FE_PHN4549_n5284), 
	.A(n5284));
   CLKBUF_X1 FE_PHC4548_n5449 (.Z(FE_PHN4548_n5449), 
	.A(n5449));
   CLKBUF_X1 FE_PHC4545_n5420 (.Z(FE_PHN4545_n5420), 
	.A(n5420));
   CLKBUF_X1 FE_PHC4544_n5770 (.Z(FE_PHN4544_n5770), 
	.A(FE_PHN1283_n5770));
   CLKBUF_X1 FE_PHC4541_n5772 (.Z(FE_PHN4541_n5772), 
	.A(FE_PHN1538_n5772));
   CLKBUF_X1 FE_PHC4540_n5297 (.Z(FE_PHN4540_n5297), 
	.A(n5297));
   CLKBUF_X1 FE_PHC4539_n5428 (.Z(FE_PHN4539_n5428), 
	.A(n5428));
   CLKBUF_X1 FE_PHC4538_n5187 (.Z(FE_PHN4538_n5187), 
	.A(n5187));
   CLKBUF_X1 FE_PHC4536_n5603 (.Z(FE_PHN4536_n5603), 
	.A(n5603));
   CLKBUF_X1 FE_PHC4535_n5641 (.Z(FE_PHN4535_n5641), 
	.A(n5641));
   CLKBUF_X1 FE_PHC4534_n5072 (.Z(FE_PHN4534_n5072), 
	.A(n5072));
   CLKBUF_X1 FE_PHC4533_n5062 (.Z(FE_PHN4533_n5062), 
	.A(n5062));
   CLKBUF_X1 FE_PHC4532_n5135 (.Z(FE_PHN4532_n5135), 
	.A(n5135));
   CLKBUF_X1 FE_PHC4531_n5174 (.Z(FE_PHN4531_n5174), 
	.A(n5174));
   CLKBUF_X1 FE_PHC4529_n5300 (.Z(FE_PHN4529_n5300), 
	.A(n5300));
   CLKBUF_X1 FE_PHC4526_U788_Z_0 (.Z(FE_PHN4526_U788_Z_0), 
	.A(U788_Z_0));
   CLKBUF_X1 FE_PHC4525_n5433 (.Z(FE_PHN4525_n5433), 
	.A(n5433));
   CLKBUF_X1 FE_PHC4524_U691_Z_0 (.Z(FE_PHN4524_U691_Z_0), 
	.A(U691_Z_0));
   CLKBUF_X1 FE_PHC4523_n5487 (.Z(FE_PHN4523_n5487), 
	.A(n5487));
   CLKBUF_X1 FE_PHC4518_n5141 (.Z(FE_PHN4518_n5141), 
	.A(n5141));
   CLKBUF_X1 FE_PHC4517_n5115 (.Z(FE_PHN4517_n5115), 
	.A(n5115));
   CLKBUF_X1 FE_PHC4516_n5288 (.Z(FE_PHN4516_n5288), 
	.A(n5288));
   CLKBUF_X1 FE_PHC4515_n5083 (.Z(FE_PHN4515_n5083), 
	.A(n5083));
   CLKBUF_X1 FE_PHC4514_n5468 (.Z(FE_PHN4514_n5468), 
	.A(n5468));
   CLKBUF_X1 FE_PHC4512_U770_Z_0 (.Z(FE_PHN4512_U770_Z_0), 
	.A(U770_Z_0));
   CLKBUF_X1 FE_PHC4511_n5170 (.Z(FE_PHN4511_n5170), 
	.A(n5170));
   CLKBUF_X1 FE_PHC4510_n5040 (.Z(FE_PHN4510_n5040), 
	.A(n5040));
   CLKBUF_X1 FE_PHC4509_n5622 (.Z(FE_PHN4509_n5622), 
	.A(n5622));
   CLKBUF_X1 FE_PHC4508_n5463 (.Z(FE_PHN4508_n5463), 
	.A(n5463));
   CLKBUF_X1 FE_PHC4506_n5470 (.Z(FE_PHN4506_n5470), 
	.A(n5470));
   CLKBUF_X1 FE_PHC4505_n5169 (.Z(FE_PHN4505_n5169), 
	.A(n5169));
   CLKBUF_X1 FE_PHC4504_n5181 (.Z(FE_PHN4504_n5181), 
	.A(n5181));
   CLKBUF_X1 FE_PHC4500_n5039 (.Z(FE_PHN4500_n5039), 
	.A(n5039));
   CLKBUF_X1 FE_PHC4499_n5138 (.Z(FE_PHN4499_n5138), 
	.A(n5138));
   CLKBUF_X1 FE_PHC4496_n5461 (.Z(FE_PHN4496_n5461), 
	.A(n5461));
   CLKBUF_X1 FE_PHC4495_n5075 (.Z(FE_PHN4495_n5075), 
	.A(n5075));
   CLKBUF_X1 FE_PHC4494_n5472 (.Z(FE_PHN4494_n5472), 
	.A(n5472));
   CLKBUF_X1 FE_PHC4493_n5557 (.Z(FE_PHN4493_n5557), 
	.A(n5557));
   CLKBUF_X1 FE_PHC4492_n5186 (.Z(FE_PHN4492_n5186), 
	.A(n5186));
   CLKBUF_X1 FE_PHC4490_n5453 (.Z(FE_PHN4490_n5453), 
	.A(n5453));
   CLKBUF_X1 FE_PHC4488_n4884 (.Z(FE_PHN4488_n4884), 
	.A(n4884));
   CLKBUF_X1 FE_PHC4487_n5478 (.Z(FE_PHN4487_n5478), 
	.A(n5478));
   CLKBUF_X1 FE_PHC4486_n4969 (.Z(FE_PHN4486_n4969), 
	.A(n4969));
   CLKBUF_X1 FE_PHC4485_n5196 (.Z(FE_PHN4485_n5196), 
	.A(n5196));
   CLKBUF_X1 FE_PHC4484_n4985 (.Z(FE_PHN4484_n4985), 
	.A(n4985));
   CLKBUF_X1 FE_PHC4482_n5455 (.Z(FE_PHN4482_n5455), 
	.A(n5455));
   CLKBUF_X1 FE_PHC4481_n5459 (.Z(FE_PHN4481_n5459), 
	.A(n5459));
   CLKBUF_X1 FE_PHC4479_U787_Z_0 (.Z(FE_PHN4479_U787_Z_0), 
	.A(U787_Z_0));
   CLKBUF_X1 FE_PHC4478_U775_Z_0 (.Z(FE_PHN4478_U775_Z_0), 
	.A(U775_Z_0));
   CLKBUF_X1 FE_PHC4477_n5173 (.Z(FE_PHN4477_n5173), 
	.A(n5173));
   CLKBUF_X1 FE_PHC4476_n5633 (.Z(FE_PHN4476_n5633), 
	.A(n5633));
   CLKBUF_X1 FE_PHC4475_n5597 (.Z(FE_PHN4475_n5597), 
	.A(n5597));
   CLKBUF_X1 FE_PHC4474_n5427 (.Z(FE_PHN4474_n5427), 
	.A(n5427));
   CLKBUF_X1 FE_PHC4472_n4869 (.Z(FE_PHN4472_n4869), 
	.A(n4869));
   CLKBUF_X1 FE_PHC4471_n5190 (.Z(FE_PHN4471_n5190), 
	.A(n5190));
   CLKBUF_X1 FE_PHC4468_n5426 (.Z(FE_PHN4468_n5426), 
	.A(n5426));
   CLKBUF_X1 FE_PHC4467_n5553 (.Z(FE_PHN4467_n5553), 
	.A(n5553));
   CLKBUF_X1 FE_PHC4466_n5312 (.Z(FE_PHN4466_n5312), 
	.A(n5312));
   CLKBUF_X1 FE_PHC4463_n5161 (.Z(FE_PHN4463_n5161), 
	.A(n5161));
   CLKBUF_X1 FE_PHC4462_n5564 (.Z(FE_PHN4462_n5564), 
	.A(n5564));
   CLKBUF_X1 FE_PHC4460_n5469 (.Z(FE_PHN4460_n5469), 
	.A(n5469));
   CLKBUF_X1 FE_PHC4459_n5401 (.Z(FE_PHN4459_n5401), 
	.A(n5401));
   CLKBUF_X1 FE_PHC4458_n5437 (.Z(FE_PHN4458_n5437), 
	.A(n5437));
   CLKBUF_X1 FE_PHC4457_n5121 (.Z(FE_PHN4457_n5121), 
	.A(n5121));
   CLKBUF_X1 FE_PHC4456_n5197 (.Z(FE_PHN4456_n5197), 
	.A(n5197));
   CLKBUF_X1 FE_PHC4454_U786_Z_0 (.Z(FE_PHN4454_U786_Z_0), 
	.A(U786_Z_0));
   CLKBUF_X1 FE_PHC4453_U459_Z_0 (.Z(FE_PHN4453_U459_Z_0), 
	.A(U459_Z_0));
   CLKBUF_X1 FE_PHC4452_n5296 (.Z(FE_PHN4452_n5296), 
	.A(n5296));
   CLKBUF_X1 FE_PHC4451_n5598 (.Z(FE_PHN4451_n5598), 
	.A(n5598));
   CLKBUF_X1 FE_PHC4450_n5486 (.Z(FE_PHN4450_n5486), 
	.A(n5486));
   CLKBUF_X1 FE_PHC4449_n5021 (.Z(FE_PHN4449_n5021), 
	.A(n5021));
   CLKBUF_X1 FE_PHC4448_n5576 (.Z(FE_PHN4448_n5576), 
	.A(n5576));
   CLKBUF_X1 FE_PHC4447_n5567 (.Z(FE_PHN4447_n5567), 
	.A(n5567));
   CLKBUF_X1 FE_PHC4446_n5093 (.Z(FE_PHN4446_n5093), 
	.A(n5093));
   CLKBUF_X1 FE_PHC4444_n5447 (.Z(FE_PHN4444_n5447), 
	.A(n5447));
   CLKBUF_X1 FE_PHC4441_U764_Z_0 (.Z(FE_PHN4441_U764_Z_0), 
	.A(FE_PHN2874_U764_Z_0));
   CLKBUF_X1 FE_PHC4440_n5616 (.Z(FE_PHN4440_n5616), 
	.A(n5616));
   CLKBUF_X1 FE_PHC4439_n5600 (.Z(FE_PHN4439_n5600), 
	.A(n5600));
   CLKBUF_X1 FE_PHC4438_n5636 (.Z(FE_PHN4438_n5636), 
	.A(n5636));
   CLKBUF_X1 FE_PHC4437_n5046 (.Z(FE_PHN4437_n5046), 
	.A(n5046));
   CLKBUF_X1 FE_PHC4436_n5464 (.Z(FE_PHN4436_n5464), 
	.A(n5464));
   CLKBUF_X1 FE_PHC4433_n5579 (.Z(FE_PHN4433_n5579), 
	.A(n5579));
   CLKBUF_X1 FE_PHC4432_n5086 (.Z(FE_PHN4432_n5086), 
	.A(n5086));
   CLKBUF_X1 FE_PHC4431_n4865 (.Z(FE_PHN4431_n4865), 
	.A(n4865));
   CLKBUF_X1 FE_PHC4430_n5485 (.Z(FE_PHN4430_n5485), 
	.A(n5485));
   CLKBUF_X1 FE_PHC4427_n5020 (.Z(FE_PHN4427_n5020), 
	.A(n5020));
   CLKBUF_X1 FE_PHC4426_n5366 (.Z(FE_PHN4426_n5366), 
	.A(n5366));
   CLKBUF_X1 FE_PHC4425_n5558 (.Z(FE_PHN4425_n5558), 
	.A(n5558));
   CLKBUF_X1 FE_PHC4422_n5392 (.Z(FE_PHN4422_n5392), 
	.A(n5392));
   CLKBUF_X1 FE_PHC4421_n5477 (.Z(FE_PHN4421_n5477), 
	.A(n5477));
   CLKBUF_X1 FE_PHC4420_n5539 (.Z(FE_PHN4420_n5539), 
	.A(n5539));
   CLKBUF_X1 FE_PHC4419_n5444 (.Z(FE_PHN4419_n5444), 
	.A(n5444));
   CLKBUF_X1 FE_PHC4418_n5022 (.Z(FE_PHN4418_n5022), 
	.A(n5022));
   CLKBUF_X1 FE_PHC4417_n5398 (.Z(FE_PHN4417_n5398), 
	.A(n5398));
   CLKBUF_X1 FE_PHC4416_n5067 (.Z(FE_PHN4416_n5067), 
	.A(n5067));
   CLKBUF_X1 FE_PHC4413_n5430 (.Z(FE_PHN4413_n5430), 
	.A(n5430));
   CLKBUF_X1 FE_PHC4412_n5442 (.Z(FE_PHN4412_n5442), 
	.A(n5442));
   CLKBUF_X1 FE_PHC4411_n5434 (.Z(FE_PHN4411_n5434), 
	.A(n5434));
   CLKBUF_X1 FE_PHC4407_n4870 (.Z(FE_PHN4407_n4870), 
	.A(n4870));
   CLKBUF_X1 FE_PHC4406_n5432 (.Z(FE_PHN4406_n5432), 
	.A(n5432));
   CLKBUF_X1 FE_PHC4405_n5476 (.Z(FE_PHN4405_n5476), 
	.A(n5476));
   CLKBUF_X1 FE_PHC4404_n5171 (.Z(FE_PHN4404_n5171), 
	.A(n5171));
   CLKBUF_X1 FE_PHC4403_n5438 (.Z(FE_PHN4403_n5438), 
	.A(n5438));
   CLKBUF_X1 FE_PHC4402_n5033 (.Z(FE_PHN4402_n5033), 
	.A(n5033));
   CLKBUF_X1 FE_PHC4401_n5287 (.Z(FE_PHN4401_n5287), 
	.A(n5287));
   CLKBUF_X1 FE_PHC4400_n5397 (.Z(FE_PHN4400_n5397), 
	.A(n5397));
   CLKBUF_X1 FE_PHC4399_n5606 (.Z(FE_PHN4399_n5606), 
	.A(n5606));
   CLKBUF_X1 FE_PHC4396_n5452 (.Z(FE_PHN4396_n5452), 
	.A(n5452));
   CLKBUF_X1 FE_PHC4394_U774_Z_0 (.Z(FE_PHN4394_U774_Z_0), 
	.A(FE_PHN2895_U774_Z_0));
   CLKBUF_X1 FE_PHC4393_n5462 (.Z(FE_PHN4393_n5462), 
	.A(n5462));
   CLKBUF_X1 FE_PHC4392_n5575 (.Z(FE_PHN4392_n5575), 
	.A(n5575));
   CLKBUF_X1 FE_PHC4387_n5069 (.Z(FE_PHN4387_n5069), 
	.A(n5069));
   CLKBUF_X1 FE_PHC4386_n5439 (.Z(FE_PHN4386_n5439), 
	.A(n5439));
   CLKBUF_X1 FE_PHC4385_n5182 (.Z(FE_PHN4385_n5182), 
	.A(n5182));
   CLKBUF_X1 FE_PHC4383_n4891 (.Z(FE_PHN4383_n4891), 
	.A(n4891));
   CLKBUF_X1 FE_PHC4382_n5424 (.Z(FE_PHN4382_n5424), 
	.A(n5424));
   CLKBUF_X1 FE_PHC4380_n5550 (.Z(FE_PHN4380_n5550), 
	.A(n5550));
   CLKBUF_X1 FE_PHC4379_n5412 (.Z(FE_PHN4379_n5412), 
	.A(n5412));
   CLKBUF_X1 FE_PHC4378_n5448 (.Z(FE_PHN4378_n5448), 
	.A(n5448));
   CLKBUF_X1 FE_PHC4377_n5421 (.Z(FE_PHN4377_n5421), 
	.A(n5421));
   CLKBUF_X1 FE_PHC4376_n5184 (.Z(FE_PHN4376_n5184), 
	.A(n5184));
   CLKBUF_X1 FE_PHC4375_n5466 (.Z(FE_PHN4375_n5466), 
	.A(n5466));
   CLKBUF_X1 FE_PHC4374_n5298 (.Z(FE_PHN4374_n5298), 
	.A(n5298));
   CLKBUF_X1 FE_PHC4373_n5030 (.Z(FE_PHN4373_n5030), 
	.A(n5030));
   CLKBUF_X1 FE_PHC4372_n5010 (.Z(FE_PHN4372_n5010), 
	.A(n5010));
   CLKBUF_X1 FE_PHC4371_n5175 (.Z(FE_PHN4371_n5175), 
	.A(n5175));
   CLKBUF_X1 FE_PHC4369_n5041 (.Z(FE_PHN4369_n5041), 
	.A(n5041));
   CLKBUF_X1 FE_PHC4368_n5123 (.Z(FE_PHN4368_n5123), 
	.A(n5123));
   CLKBUF_X1 FE_PHC4367_n5411 (.Z(FE_PHN4367_n5411), 
	.A(n5411));
   CLKBUF_X1 FE_PHC4366_n5414 (.Z(FE_PHN4366_n5414), 
	.A(n5414));
   CLKBUF_X1 FE_PHC4364_n5074 (.Z(FE_PHN4364_n5074), 
	.A(n5074));
   CLKBUF_X1 FE_PHC4363_n5108 (.Z(FE_PHN4363_n5108), 
	.A(n5108));
   CLKBUF_X1 FE_PHC4362_n5043 (.Z(FE_PHN4362_n5043), 
	.A(n5043));
   CLKBUF_X1 FE_PHC4361_n4987 (.Z(FE_PHN4361_n4987), 
	.A(n4987));
   CLKBUF_X1 FE_PHC4358_n4872 (.Z(FE_PHN4358_n4872), 
	.A(n4872));
   CLKBUF_X1 FE_PHC4357_n5192 (.Z(FE_PHN4357_n5192), 
	.A(n5192));
   CLKBUF_X1 FE_PHC4356_n5191 (.Z(FE_PHN4356_n5191), 
	.A(n5191));
   CLKBUF_X1 FE_PHC4355_n5441 (.Z(FE_PHN4355_n5441), 
	.A(n5441));
   CLKBUF_X1 FE_PHC4352_n5473 (.Z(FE_PHN4352_n5473), 
	.A(n5473));
   CLKBUF_X1 FE_PHC4351_n5051 (.Z(FE_PHN4351_n5051), 
	.A(n5051));
   CLKBUF_X1 FE_PHC4350_n5091 (.Z(FE_PHN4350_n5091), 
	.A(n5091));
   CLKBUF_X1 FE_PHC4348_n5410 (.Z(FE_PHN4348_n5410), 
	.A(n5410));
   CLKBUF_X1 FE_PHC4346_n5316 (.Z(FE_PHN4346_n5316), 
	.A(n5316));
   CLKBUF_X1 FE_PHC4343_n5419 (.Z(FE_PHN4343_n5419), 
	.A(n5419));
   CLKBUF_X1 FE_PHC4340_n5106 (.Z(FE_PHN4340_n5106), 
	.A(n5106));
   CLKBUF_X1 FE_PHC4338_n5132 (.Z(FE_PHN4338_n5132), 
	.A(n5132));
   CLKBUF_X1 FE_PHC4337_n5509 (.Z(FE_PHN4337_n5509), 
	.A(n5509));
   CLKBUF_X1 FE_PHC4336_n5304 (.Z(FE_PHN4336_n5304), 
	.A(n5304));
   CLKBUF_X1 FE_PHC4335_n5386 (.Z(FE_PHN4335_n5386), 
	.A(n5386));
   CLKBUF_X1 FE_PHC4334_n5393 (.Z(FE_PHN4334_n5393), 
	.A(n5393));
   CLKBUF_X1 FE_PHC4333_n5395 (.Z(FE_PHN4333_n5395), 
	.A(n5395));
   CLKBUF_X1 FE_PHC4332_n5180 (.Z(FE_PHN4332_n5180), 
	.A(n5180));
   CLKBUF_X1 FE_PHC4331_n5399 (.Z(FE_PHN4331_n5399), 
	.A(n5399));
   CLKBUF_X1 FE_PHC4330_n5435 (.Z(FE_PHN4330_n5435), 
	.A(n5435));
   CLKBUF_X1 FE_PHC4329_n5205 (.Z(FE_PHN4329_n5205), 
	.A(n5205));
   CLKBUF_X1 FE_PHC4327_n5183 (.Z(FE_PHN4327_n5183), 
	.A(n5183));
   CLKBUF_X1 FE_PHC4326_U279_Z_0 (.Z(FE_PHN4326_U279_Z_0), 
	.A(U279_Z_0));
   CLKBUF_X1 FE_PHC4325_n4986 (.Z(FE_PHN4325_n4986), 
	.A(n4986));
   CLKBUF_X1 FE_PHC4324_U105_Z_0 (.Z(FE_PHN4324_U105_Z_0), 
	.A(FE_PHN1654_U105_Z_0));
   CLKBUF_X1 FE_PHC4322_U780_Z_0 (.Z(FE_PHN4322_U780_Z_0), 
	.A(U780_Z_0));
   CLKBUF_X1 FE_PHC4320_n5451 (.Z(FE_PHN4320_n5451), 
	.A(n5451));
   BUF_X1 FE_PHC4319_n5189 (.Z(FE_PHN4319_n5189), 
	.A(n5189));
   CLKBUF_X1 FE_PHC4318_n5521 (.Z(FE_PHN4318_n5521), 
	.A(n5521));
   CLKBUF_X1 FE_PHC4317_n5289 (.Z(FE_PHN4317_n5289), 
	.A(n5289));
   CLKBUF_X1 FE_PHC4316_n5799 (.Z(FE_PHN4316_n5799), 
	.A(FE_PHN2899_n5799));
   CLKBUF_X1 FE_PHC4314_n5629 (.Z(FE_PHN4314_n5629), 
	.A(n5629));
   CLKBUF_X1 FE_PHC4313_n5596 (.Z(FE_PHN4313_n5596), 
	.A(n5596));
   CLKBUF_X1 FE_PHC4312_n5199 (.Z(FE_PHN4312_n5199), 
	.A(n5199));
   CLKBUF_X1 FE_PHC4311_n5195 (.Z(FE_PHN4311_n5195), 
	.A(n5195));
   CLKBUF_X1 FE_PHC4305_n5422 (.Z(FE_PHN4305_n5422), 
	.A(n5422));
   CLKBUF_X1 FE_PHC4303_U766_Z_0 (.Z(FE_PHN4303_U766_Z_0), 
	.A(FE_PHN2857_U766_Z_0));
   CLKBUF_X1 FE_PHC4302_n5440 (.Z(FE_PHN4302_n5440), 
	.A(n5440));
   CLKBUF_X1 FE_PHC4301_n5409 (.Z(FE_PHN4301_n5409), 
	.A(n5409));
   CLKBUF_X1 FE_PHC4298_U785_Z_0 (.Z(FE_PHN4298_U785_Z_0), 
	.A(U785_Z_0));
   CLKBUF_X1 FE_PHC4297_U261_Z_0 (.Z(FE_PHN4297_U261_Z_0), 
	.A(U261_Z_0));
   CLKBUF_X1 FE_PHC4295_n5436 (.Z(FE_PHN4295_n5436), 
	.A(n5436));
   CLKBUF_X1 FE_PHC4291_n5207 (.Z(FE_PHN4291_n5207), 
	.A(n5207));
   CLKBUF_X1 FE_PHC4289_n4854 (.Z(FE_PHN4289_n4854), 
	.A(n4854));
   CLKBUF_X1 FE_PHC4288_n1319 (.Z(FE_PHN4288_n1319), 
	.A(n1319));
   CLKBUF_X1 FE_PHC4287_n5415 (.Z(FE_PHN4287_n5415), 
	.A(n5415));
   CLKBUF_X1 FE_PHC4283_n5309 (.Z(FE_PHN4283_n5309), 
	.A(n5309));
   CLKBUF_X1 FE_PHC4282_n5418 (.Z(FE_PHN4282_n5418), 
	.A(n5418));
   CLKBUF_X1 FE_PHC4280_n5624 (.Z(FE_PHN4280_n5624), 
	.A(n5624));
   CLKBUF_X1 FE_PHC4279_n5301 (.Z(FE_PHN4279_n5301), 
	.A(n5301));
   CLKBUF_X1 FE_PHC4274_n5176 (.Z(FE_PHN4274_n5176), 
	.A(n5176));
   CLKBUF_X1 FE_PHC4273_n5225 (.Z(FE_PHN4273_n5225), 
	.A(n5225));
   CLKBUF_X1 FE_PHC4272_U479_Z_0 (.Z(FE_PHN4272_U479_Z_0), 
	.A(U479_Z_0));
   CLKBUF_X1 FE_PHC4271_n5159 (.Z(FE_PHN4271_n5159), 
	.A(n5159));
   CLKBUF_X1 FE_PHC4270_U509_Z_0 (.Z(FE_PHN4270_U509_Z_0), 
	.A(U509_Z_0));
   CLKBUF_X1 FE_PHC4269_U429_Z_0 (.Z(FE_PHN4269_U429_Z_0), 
	.A(U429_Z_0));
   CLKBUF_X1 FE_PHC4267_n5363 (.Z(FE_PHN4267_n5363), 
	.A(n5363));
   CLKBUF_X1 FE_PHC4266_n5483 (.Z(FE_PHN4266_n5483), 
	.A(n5483));
   CLKBUF_X1 FE_PHC4264_U777_Z_0 (.Z(FE_PHN4264_U777_Z_0), 
	.A(U777_Z_0));
   CLKBUF_X1 FE_PHC4263_n5028 (.Z(FE_PHN4263_n5028), 
	.A(n5028));
   CLKBUF_X1 FE_PHC4262_n5013 (.Z(FE_PHN4262_n5013), 
	.A(n5013));
   CLKBUF_X1 FE_PHC4261_n5481 (.Z(FE_PHN4261_n5481), 
	.A(n5481));
   CLKBUF_X1 FE_PHC4260_n5045 (.Z(FE_PHN4260_n5045), 
	.A(n5045));
   CLKBUF_X1 FE_PHC4259_n5049 (.Z(FE_PHN4259_n5049), 
	.A(n5049));
   CLKBUF_X1 FE_PHC4258_n5081 (.Z(FE_PHN4258_n5081), 
	.A(n5081));
   CLKBUF_X1 FE_PHC4257_n5318 (.Z(FE_PHN4257_n5318), 
	.A(n5318));
   CLKBUF_X1 FE_PHC4249_n5308 (.Z(FE_PHN4249_n5308), 
	.A(n5308));
   CLKBUF_X1 FE_PHC4248_n5203 (.Z(FE_PHN4248_n5203), 
	.A(n5203));
   CLKBUF_X1 FE_PHC4247_n5270 (.Z(FE_PHN4247_n5270), 
	.A(n5270));
   CLKBUF_X1 FE_PHC4240_n5364 (.Z(FE_PHN4240_n5364), 
	.A(n5364));
   CLKBUF_X1 FE_PHC4237_n5076 (.Z(FE_PHN4237_n5076), 
	.A(n5076));
   CLKBUF_X1 FE_PHC4235_n5413 (.Z(FE_PHN4235_n5413), 
	.A(n5413));
   BUF_X1 FE_PHC4234_n5224 (.Z(FE_PHN4234_n5224), 
	.A(n5224));
   CLKBUF_X1 FE_PHC4233_n5542 (.Z(FE_PHN4233_n5542), 
	.A(n5542));
   CLKBUF_X1 FE_PHC4232_U359_Z_0 (.Z(FE_PHN4232_U359_Z_0), 
	.A(U359_Z_0));
   CLKBUF_X1 FE_PHC4231_n5443 (.Z(FE_PHN4231_n5443), 
	.A(n5443));
   CLKBUF_X1 FE_PHC4230_n5268 (.Z(FE_PHN4230_n5268), 
	.A(n5268));
   CLKBUF_X1 FE_PHC4229_U761_Z_0 (.Z(FE_PHN4229_U761_Z_0), 
	.A(U761_Z_0));
   CLKBUF_X1 FE_PHC4227_n5317 (.Z(FE_PHN4227_n5317), 
	.A(n5317));
   CLKBUF_X1 FE_PHC4221_n5360 (.Z(FE_PHN4221_n5360), 
	.A(n5360));
   CLKBUF_X1 FE_PHC4220_n5361 (.Z(FE_PHN4220_n5361), 
	.A(n5361));
   CLKBUF_X1 FE_PHC4219_n4979 (.Z(FE_PHN4219_n4979), 
	.A(n4979));
   CLKBUF_X1 FE_PHC4218_n5202 (.Z(FE_PHN4218_n5202), 
	.A(n5202));
   CLKBUF_X1 FE_PHC4217_n5079 (.Z(FE_PHN4217_n5079), 
	.A(n5079));
   CLKBUF_X1 FE_PHC4216_n5514 (.Z(FE_PHN4216_n5514), 
	.A(n5514));
   CLKBUF_X1 FE_PHC4215_n5638 (.Z(FE_PHN4215_n5638), 
	.A(n5638));
   CLKBUF_X1 FE_PHC4214_n5621 (.Z(FE_PHN4214_n5621), 
	.A(n5621));
   CLKBUF_X1 FE_PHC4213_n5391 (.Z(FE_PHN4213_n5391), 
	.A(n5391));
   CLKBUF_X1 FE_PHC4212_U590_Z_0 (.Z(FE_PHN4212_U590_Z_0), 
	.A(U590_Z_0));
   CLKBUF_X1 FE_PHC4205_n5538 (.Z(FE_PHN4205_n5538), 
	.A(n5538));
   CLKBUF_X1 FE_PHC4202_U784_Z_0 (.Z(FE_PHN4202_U784_Z_0), 
	.A(U784_Z_0));
   CLKBUF_X1 FE_PHC4201_n5643 (.Z(FE_PHN4201_n5643), 
	.A(n5643));
   CLKBUF_X1 FE_PHC4200_n5112 (.Z(FE_PHN4200_n5112), 
	.A(n5112));
   CLKBUF_X1 FE_PHC4199_n5369 (.Z(FE_PHN4199_n5369), 
	.A(n5369));
   CLKBUF_X1 FE_PHC4198_n5209 (.Z(FE_PHN4198_n5209), 
	.A(n5209));
   CLKBUF_X1 FE_PHC4196_U275_Z_0 (.Z(FE_PHN4196_U275_Z_0), 
	.A(U275_Z_0));
   CLKBUF_X1 FE_PHC4193_n5266 (.Z(FE_PHN4193_n5266), 
	.A(n5266));
   CLKBUF_X1 FE_PHC4192_n5384 (.Z(FE_PHN4192_n5384), 
	.A(n5384));
   CLKBUF_X1 FE_PHC4191_n5018 (.Z(FE_PHN4191_n5018), 
	.A(n5018));
   CLKBUF_X1 FE_PHC4187_n4995 (.Z(FE_PHN4187_n4995), 
	.A(n4995));
   CLKBUF_X1 FE_PHC4185_n5511 (.Z(FE_PHN4185_n5511), 
	.A(n5511));
   CLKBUF_X1 FE_PHC4182_n5348 (.Z(FE_PHN4182_n5348), 
	.A(n5348));
   CLKBUF_X1 FE_PHC4181_n5554 (.Z(FE_PHN4181_n5554), 
	.A(n5554));
   CLKBUF_X1 FE_PHC4180_n5610 (.Z(FE_PHN4180_n5610), 
	.A(n5610));
   CLKBUF_X1 FE_PHC4178_n5070 (.Z(FE_PHN4178_n5070), 
	.A(n5070));
   CLKBUF_X1 FE_PHC4177_n5273 (.Z(FE_PHN4177_n5273), 
	.A(n5273));
   CLKBUF_X1 FE_PHC4176_n5394 (.Z(FE_PHN4176_n5394), 
	.A(n5394));
   CLKBUF_X1 FE_PHC4175_n5200 (.Z(FE_PHN4175_n5200), 
	.A(n5200));
   CLKBUF_X1 FE_PHC4174_U243_Z_0 (.Z(FE_PHN4174_U243_Z_0), 
	.A(U243_Z_0));
   CLKBUF_X1 FE_PHC4172_n5367 (.Z(FE_PHN4172_n5367), 
	.A(n5367));
   CLKBUF_X1 FE_PHC4171_n5019 (.Z(FE_PHN4171_n5019), 
	.A(n5019));
   CLKBUF_X1 FE_PHC4170_n5319 (.Z(FE_PHN4170_n5319), 
	.A(n5319));
   CLKBUF_X1 FE_PHC4169_n5261 (.Z(FE_PHN4169_n5261), 
	.A(n5261));
   CLKBUF_X1 FE_PHC4168_n5136 (.Z(FE_PHN4168_n5136), 
	.A(n5136));
   CLKBUF_X1 FE_PHC4167_n5139 (.Z(FE_PHN4167_n5139), 
	.A(n5139));
   CLKBUF_X1 FE_PHC4166_n5133 (.Z(FE_PHN4166_n5133), 
	.A(n5133));
   CLKBUF_X1 FE_PHC4165_n5280 (.Z(FE_PHN4165_n5280), 
	.A(n5280));
   CLKBUF_X1 FE_PHC4161_n5107 (.Z(FE_PHN4161_n5107), 
	.A(n5107));
   CLKBUF_X1 FE_PHC4160_n5218 (.Z(FE_PHN4160_n5218), 
	.A(n5218));
   CLKBUF_X1 FE_PHC4154_n5213 (.Z(FE_PHN4154_n5213), 
	.A(n5213));
   CLKBUF_X1 FE_PHC4150_n5362 (.Z(FE_PHN4150_n5362), 
	.A(n5362));
   CLKBUF_X1 FE_PHC4149_n5560 (.Z(FE_PHN4149_n5560), 
	.A(n5560));
   CLKBUF_X1 FE_PHC4148_n5383 (.Z(FE_PHN4148_n5383), 
	.A(n5383));
   CLKBUF_X1 FE_PHC4147_n5279 (.Z(FE_PHN4147_n5279), 
	.A(n5279));
   CLKBUF_X1 FE_PHC4146_n5357 (.Z(FE_PHN4146_n5357), 
	.A(n5357));
   CLKBUF_X1 FE_PHC4145_n5405 (.Z(FE_PHN4145_n5405), 
	.A(n5405));
   CLKBUF_X1 FE_PHC4142_n5365 (.Z(FE_PHN4142_n5365), 
	.A(n5365));
   CLKBUF_X1 FE_PHC4141_n5376 (.Z(FE_PHN4141_n5376), 
	.A(n5376));
   CLKBUF_X1 FE_PHC4140_n5217 (.Z(FE_PHN4140_n5217), 
	.A(n5217));
   CLKBUF_X1 FE_PHC4139_n5611 (.Z(FE_PHN4139_n5611), 
	.A(n5611));
   BUF_X2 FE_PHC4138_U295_Z_0 (.Z(FE_PHN4138_U295_Z_0), 
	.A(U295_Z_0));
   CLKBUF_X1 FE_PHC4136_n5640 (.Z(FE_PHN4136_n5640), 
	.A(n5640));
   CLKBUF_X1 FE_PHC4135_n5339 (.Z(FE_PHN4135_n5339), 
	.A(n5339));
   CLKBUF_X1 FE_PHC4133_n4874 (.Z(FE_PHN4133_n4874), 
	.A(n4874));
   CLKBUF_X1 FE_PHC4132_n5517 (.Z(FE_PHN4132_n5517), 
	.A(n5517));
   CLKBUF_X1 FE_PHC4129_n5201 (.Z(FE_PHN4129_n5201), 
	.A(n5201));
   BUF_X8 FE_PHC4126_n5776 (.Z(FE_PHN4126_n5776), 
	.A(FE_PHN2028_n5776));
   CLKBUF_X1 FE_PHC4124_n5356 (.Z(FE_PHN4124_n5356), 
	.A(n5356));
   CLKBUF_X1 FE_PHC4123_n5124 (.Z(FE_PHN4123_n5124), 
	.A(n5124));
   CLKBUF_X1 FE_PHC4122_n5489 (.Z(FE_PHN4122_n5489), 
	.A(n5489));
   CLKBUF_X1 FE_PHC4120_n5403 (.Z(FE_PHN4120_n5403), 
	.A(n5403));
   CLKBUF_X1 FE_PHC4119_n5294 (.Z(FE_PHN4119_n5294), 
	.A(n5294));
   CLKBUF_X1 FE_PHC4118_n5277 (.Z(FE_PHN4118_n5277), 
	.A(n5277));
   CLKBUF_X1 FE_PHC4117_n5084 (.Z(FE_PHN4117_n5084), 
	.A(n5084));
   CLKBUF_X1 FE_PHC4115_n5335 (.Z(FE_PHN4115_n5335), 
	.A(n5335));
   CLKBUF_X1 FE_PHC4109_n5219 (.Z(FE_PHN4109_n5219), 
	.A(n5219));
   CLKBUF_X1 FE_PHC4108_n5599 (.Z(FE_PHN4108_n5599), 
	.A(n5599));
   CLKBUF_X1 FE_PHC4104_n4878 (.Z(FE_PHN4104_n4878), 
	.A(n4878));
   CLKBUF_X1 FE_PHC4102_n5109 (.Z(FE_PHN4102_n5109), 
	.A(n5109));
   CLKBUF_X1 FE_PHC4101_n5562 (.Z(FE_PHN4101_n5562), 
	.A(n5562));
   CLKBUF_X1 FE_PHC4096_U506_Z_0 (.Z(FE_PHN4096_U506_Z_0), 
	.A(U506_Z_0));
   CLKBUF_X1 FE_PHC4094_n5492 (.Z(FE_PHN4094_n5492), 
	.A(n5492));
   CLKBUF_X1 FE_PHC4093_n5493 (.Z(FE_PHN4093_n5493), 
	.A(n5493));
   CLKBUF_X1 FE_PHC4090_n5349 (.Z(FE_PHN4090_n5349), 
	.A(n5349));
   CLKBUF_X1 FE_PHC4089_n5352 (.Z(FE_PHN4089_n5352), 
	.A(n5352));
   CLKBUF_X1 FE_PHC4088_n5496 (.Z(FE_PHN4088_n5496), 
	.A(n5496));
   CLKBUF_X1 FE_PHC4085_n5374 (.Z(FE_PHN4085_n5374), 
	.A(n5374));
   CLKBUF_X1 FE_PHC4084_n5479 (.Z(FE_PHN4084_n5479), 
	.A(n5479));
   CLKBUF_X1 FE_PHC4083_n5347 (.Z(FE_PHN4083_n5347), 
	.A(n5347));
   CLKBUF_X1 FE_PHC4082_n5334 (.Z(FE_PHN4082_n5334), 
	.A(n5334));
   CLKBUF_X1 FE_PHC4078_n5508 (.Z(FE_PHN4078_n5508), 
	.A(n5508));
   CLKBUF_X1 FE_PHC4077_n5480 (.Z(FE_PHN4077_n5480), 
	.A(n5480));
   CLKBUF_X1 FE_PHC4076_n5044 (.Z(FE_PHN4076_n5044), 
	.A(n5044));
   CLKBUF_X1 FE_PHC4072_n5221 (.Z(FE_PHN4072_n5221), 
	.A(n5221));
   CLKBUF_X1 FE_PHC4067_n5292 (.Z(FE_PHN4067_n5292), 
	.A(n5292));
   CLKBUF_X1 FE_PHC4061_n5630 (.Z(FE_PHN4061_n5630), 
	.A(n5630));
   CLKBUF_X1 FE_PHC4060_n5278 (.Z(FE_PHN4060_n5278), 
	.A(n5278));
   CLKBUF_X1 FE_PHC4059_n5491 (.Z(FE_PHN4059_n5491), 
	.A(n5491));
   CLKBUF_X1 FE_PHC4058_n5089 (.Z(FE_PHN4058_n5089), 
	.A(n5089));
   CLKBUF_X1 FE_PHC4057_n5378 (.Z(FE_PHN4057_n5378), 
	.A(n5378));
   CLKBUF_X1 FE_PHC4054_U475_Z_0 (.Z(FE_PHN4054_U475_Z_0), 
	.A(U475_Z_0));
   CLKBUF_X1 FE_PHC4053_U660_Z_0 (.Z(FE_PHN4053_U660_Z_0), 
	.A(U660_Z_0));
   CLKBUF_X1 FE_PHC4052_n5355 (.Z(FE_PHN4052_n5355), 
	.A(n5355));
   CLKBUF_X1 FE_PHC4051_n5286 (.Z(FE_PHN4051_n5286), 
	.A(n5286));
   CLKBUF_X1 FE_PHC4050_n5635 (.Z(FE_PHN4050_n5635), 
	.A(n5635));
   CLKBUF_X1 FE_PHC4048_U726_Z_0 (.Z(FE_PHN4048_U726_Z_0), 
	.A(U726_Z_0));
   BUF_X8 FE_PHC4047_U257_Z_0 (.Z(FE_PHN4047_U257_Z_0), 
	.A(U257_Z_0));
   CLKBUF_X1 FE_PHC4044_n5271 (.Z(FE_PHN4044_n5271), 
	.A(n5271));
   CLKBUF_X1 FE_PHC4043_n5336 (.Z(FE_PHN4043_n5336), 
	.A(n5336));
   CLKBUF_X1 FE_PHC4042_n5372 (.Z(FE_PHN4042_n5372), 
	.A(n5372));
   CLKBUF_X1 FE_PHC4041_n5214 (.Z(FE_PHN4041_n5214), 
	.A(n5214));
   CLKBUF_X1 FE_PHC4040_n5052 (.Z(FE_PHN4040_n5052), 
	.A(n5052));
   CLKBUF_X1 FE_PHC4039_U441_Z_0 (.Z(FE_PHN4039_U441_Z_0), 
	.A(FE_PHN2879_U441_Z_0));
   CLKBUF_X1 FE_PHC4035_U779_Z_0 (.Z(FE_PHN4035_U779_Z_0), 
	.A(U779_Z_0));
   CLKBUF_X1 FE_PHC4034_U606_Z_0 (.Z(FE_PHN4034_U606_Z_0), 
	.A(U606_Z_0));
   CLKBUF_X1 FE_PHC4032_n5128 (.Z(FE_PHN4032_n5128), 
	.A(n5128));
   CLKBUF_X1 FE_PHC4031_n5220 (.Z(FE_PHN4031_n5220), 
	.A(n5220));
   CLKBUF_X1 FE_PHC4027_n5343 (.Z(FE_PHN4027_n5343), 
	.A(n5343));
   CLKBUF_X1 FE_PHC4026_n5337 (.Z(FE_PHN4026_n5337), 
	.A(n5337));
   CLKBUF_X1 FE_PHC4024_U411_Z_0 (.Z(FE_PHN4024_U411_Z_0), 
	.A(U411_Z_0));
   CLKBUF_X1 FE_PHC4023_U673_Z_0 (.Z(FE_PHN4023_U673_Z_0), 
	.A(U673_Z_0));
   CLKBUF_X1 FE_PHC4022_n5350 (.Z(FE_PHN4022_n5350), 
	.A(n5350));
   CLKBUF_X1 FE_PHC4021_n5617 (.Z(FE_PHN4021_n5617), 
	.A(n5617));
   CLKBUF_X1 FE_PHC4020_n5541 (.Z(FE_PHN4020_n5541), 
	.A(n5541));
   CLKBUF_X1 FE_PHC4018_n5566 (.Z(FE_PHN4018_n5566), 
	.A(n5566));
   CLKBUF_X1 FE_PHC4017_n5379 (.Z(FE_PHN4017_n5379), 
	.A(n5379));
   CLKBUF_X1 FE_PHC4012_n5602 (.Z(FE_PHN4012_n5602), 
	.A(n5602));
   CLKBUF_X1 FE_PHC4005_n4998 (.Z(FE_PHN4005_n4998), 
	.A(n4998));
   CLKBUF_X1 FE_PHC4004_n5211 (.Z(FE_PHN4004_n5211), 
	.A(n5211));
   CLKBUF_X1 FE_PHC4003_n5063 (.Z(FE_PHN4003_n5063), 
	.A(n5063));
   CLKBUF_X1 FE_PHC4002_n5104 (.Z(FE_PHN4002_n5104), 
	.A(n5104));
   CLKBUF_X1 FE_PHC4001_n5087 (.Z(FE_PHN4001_n5087), 
	.A(n5087));
   BUF_X8 FE_PHC4000_n4984 (.Z(FE_PHN4000_n4984), 
	.A(n4984));
   BUF_X8 FE_PHC3989_U448_Z_0 (.Z(FE_PHN3989_U448_Z_0), 
	.A(U448_Z_0));
   CLKBUF_X1 FE_PHC3987_n5216 (.Z(FE_PHN3987_n5216), 
	.A(n5216));
   CLKBUF_X1 FE_PHC3986_n5497 (.Z(FE_PHN3986_n5497), 
	.A(n5497));
   CLKBUF_X1 FE_PHC3985_n5577 (.Z(FE_PHN3985_n5577), 
	.A(n5577));
   CLKBUF_X1 FE_PHC3983_n5263 (.Z(FE_PHN3983_n5263), 
	.A(n5263));
   CLKBUF_X1 FE_PHC3982_n5260 (.Z(FE_PHN3982_n5260), 
	.A(n5260));
   CLKBUF_X1 FE_PHC3981_n5559 (.Z(FE_PHN3981_n5559), 
	.A(n5559));
   CLKBUF_X1 FE_PHC3977_n5495 (.Z(FE_PHN3977_n5495), 
	.A(n5495));
   CLKBUF_X2 FE_PHC3976_U395_Z_0 (.Z(FE_PHN3976_U395_Z_0), 
	.A(U395_Z_0));
   CLKBUF_X1 FE_PHC3975_n5385 (.Z(FE_PHN3975_n5385), 
	.A(n5385));
   CLKBUF_X1 FE_PHC3974_n5381 (.Z(FE_PHN3974_n5381), 
	.A(n5381));
   CLKBUF_X1 FE_PHC3973_n5042 (.Z(FE_PHN3973_n5042), 
	.A(n5042));
   CLKBUF_X1 FE_PHC3972_n5490 (.Z(FE_PHN3972_n5490), 
	.A(n5490));
   CLKBUF_X1 FE_PHC3971_U291_Z_0 (.Z(FE_PHN3971_U291_Z_0), 
	.A(U291_Z_0));
   CLKBUF_X1 FE_PHC3970_n5037 (.Z(FE_PHN3970_n5037), 
	.A(n5037));
   CLKBUF_X1 FE_PHC3969_n5092 (.Z(FE_PHN3969_n5092), 
	.A(n5092));
   CLKBUF_X1 FE_PHC3963_n5125 (.Z(FE_PHN3963_n5125), 
	.A(n5125));
   CLKBUF_X1 FE_PHC3962_n5634 (.Z(FE_PHN3962_n5634), 
	.A(n5634));
   CLKBUF_X1 FE_PHC3961_n5283 (.Z(FE_PHN3961_n5283), 
	.A(n5283));
   CLKBUF_X1 FE_PHC3960_n5631 (.Z(FE_PHN3960_n5631), 
	.A(n5631));
   CLKBUF_X1 FE_PHC3959_n5608 (.Z(FE_PHN3959_n5608), 
	.A(n5608));
   CLKBUF_X1 FE_PHC3958_n5353 (.Z(FE_PHN3958_n5353), 
	.A(n5353));
   CLKBUF_X1 FE_PHC3954_n5569 (.Z(FE_PHN3954_n5569), 
	.A(n5569));
   CLKBUF_X1 FE_PHC3950_U325_Z_0 (.Z(FE_PHN3950_U325_Z_0), 
	.A(U325_Z_0));
   CLKBUF_X1 FE_PHC3949_n5382 (.Z(FE_PHN3949_n5382), 
	.A(n5382));
   CLKBUF_X1 FE_PHC3948_n5198 (.Z(FE_PHN3948_n5198), 
	.A(n5198));
   CLKBUF_X1 FE_PHC3943_n5307 (.Z(FE_PHN3943_n5307), 
	.A(n5307));
   CLKBUF_X1 FE_PHC3942_n5563 (.Z(FE_PHN3942_n5563), 
	.A(n5563));
   CLKBUF_X1 FE_PHC3941_n5548 (.Z(FE_PHN3941_n5548), 
	.A(n5548));
   CLKBUF_X1 FE_PHC3937_n5131 (.Z(FE_PHN3937_n5131), 
	.A(n5131));
   BUF_X8 FE_PHC3934_n4875 (.Z(FE_PHN3934_n4875), 
	.A(n4875));
   CLKBUF_X1 FE_PHC3931_n5368 (.Z(FE_PHN3931_n5368), 
	.A(n5368));
   CLKBUF_X1 FE_PHC3930_n5275 (.Z(FE_PHN3930_n5275), 
	.A(n5275));
   CLKBUF_X1 FE_PHC3928_n5515 (.Z(FE_PHN3928_n5515), 
	.A(n5515));
   BUF_X8 FE_PHC3927_n5116 (.Z(FE_PHN3927_n5116), 
	.A(n5116));
   CLKBUF_X1 FE_PHC3926_n5574 (.Z(FE_PHN3926_n5574), 
	.A(n5574));
   BUF_X8 FE_PHC3925_U329_Z_0 (.Z(FE_PHN3925_U329_Z_0), 
	.A(U329_Z_0));
   CLKBUF_X1 FE_PHC3924_n5607 (.Z(FE_PHN3924_n5607), 
	.A(n5607));
   BUF_X8 FE_PHC3923_n5351 (.Z(FE_PHN3923_n5351), 
	.A(n5351));
   CLKBUF_X1 FE_PHC3922_n5627 (.Z(FE_PHN3922_n5627), 
	.A(n5627));
   BUF_X8 FE_PHC3921_n5204 (.Z(FE_PHN3921_n5204), 
	.A(n5204));
   CLKBUF_X1 FE_PHC3919_n5122 (.Z(FE_PHN3919_n5122), 
	.A(n5122));
   CLKBUF_X1 FE_PHC3918_n5264 (.Z(FE_PHN3918_n5264), 
	.A(n5264));
   CLKBUF_X1 FE_PHC3917_n5226 (.Z(FE_PHN3917_n5226), 
	.A(n5226));
   CLKBUF_X1 FE_PHC3916_n5073 (.Z(FE_PHN3916_n5073), 
	.A(n5073));
   CLKBUF_X1 FE_PHC3915_n5380 (.Z(FE_PHN3915_n5380), 
	.A(n5380));
   BUF_X8 FE_PHC3912_n5212 (.Z(FE_PHN3912_n5212), 
	.A(n5212));
   CLKBUF_X1 FE_PHC3911_n5276 (.Z(FE_PHN3911_n5276), 
	.A(n5276));
   BUF_X8 FE_PHC3910_n5370 (.Z(FE_PHN3910_n5370), 
	.A(n5370));
   CLKBUF_X1 FE_PHC3909_n5215 (.Z(FE_PHN3909_n5215), 
	.A(n5215));
   CLKBUF_X1 FE_PHC3908_n5543 (.Z(FE_PHN3908_n5543), 
	.A(n5543));
   CLKBUF_X1 FE_PHC3907_n5494 (.Z(FE_PHN3907_n5494), 
	.A(n5494));
   BUF_X8 FE_PHC3906_n5016 (.Z(FE_PHN3906_n5016), 
	.A(n5016));
   BUF_X8 FE_PHC3904_U624_Z_0 (.Z(FE_PHN3904_U624_Z_0), 
	.A(U624_Z_0));
   BUF_X8 FE_PHC3903_U644_Z_0 (.Z(FE_PHN3903_U644_Z_0), 
	.A(U644_Z_0));
   BUF_X8 FE_PHC3902_n5650 (.Z(FE_PHN3902_n5650), 
	.A(n5650));
   BUF_X8 FE_PHC3900_U386_Z_0 (.Z(FE_PHN3900_U386_Z_0), 
	.A(U386_Z_0));
   CLKBUF_X1 FE_PHC3898_n5389 (.Z(FE_PHN3898_n5389), 
	.A(n5389));
   CLKBUF_X1 FE_PHC3896_n5345 (.Z(FE_PHN3896_n5345), 
	.A(n5345));
   CLKBUF_X1 FE_PHC3893_n5341 (.Z(FE_PHN3893_n5341), 
	.A(n5341));
   CLKBUF_X1 FE_PHC3892_n5210 (.Z(FE_PHN3892_n5210), 
	.A(n5210));
   CLKBUF_X1 FE_PHC3888_n5614 (.Z(FE_PHN3888_n5614), 
	.A(n5614));
   CLKBUF_X2 FE_PHC3887_U712_Z_0 (.Z(FE_PHN3887_U712_Z_0), 
	.A(U712_Z_0));
   BUF_X8 FE_PHC3886_n5262 (.Z(FE_PHN3886_n5262), 
	.A(n5262));
   BUF_X8 FE_PHC3885_U239_Z_0 (.Z(FE_PHN3885_U239_Z_0), 
	.A(U239_Z_0));
   CLKBUF_X1 FE_PHC3884_n5354 (.Z(FE_PHN3884_n5354), 
	.A(n5354));
   CLKBUF_X1 FE_PHC3883_n4963 (.Z(FE_PHN3883_n4963), 
	.A(n4963));
   CLKBUF_X1 FE_PHC3882_U466_Z_0 (.Z(FE_PHN3882_U466_Z_0), 
	.A(U466_Z_0));
   BUF_X8 FE_PHC3880_n5738 (.Z(FE_PHN3880_n5738), 
	.A(FE_PHN4916_n5738));
   CLKBUF_X1 FE_PHC3879_n5340 (.Z(FE_PHN3879_n5340), 
	.A(n5340));
   BUF_X8 FE_PHC3878_U353_Z_0 (.Z(FE_PHN3878_U353_Z_0), 
	.A(FE_PHN2883_U353_Z_0));
   BUF_X8 FE_PHC3877_U234_Z_0 (.Z(FE_PHN3877_U234_Z_0), 
	.A(U234_Z_0));
   CLKBUF_X1 FE_PHC3875_n5390 (.Z(FE_PHN3875_n5390), 
	.A(n5390));
   BUF_X8 FE_PHC3874_n5142 (.Z(FE_PHN3874_n5142), 
	.A(n5142));
   BUF_X8 FE_PHC3872_n5066 (.Z(FE_PHN3872_n5066), 
	.A(n5066));
   CLKBUF_X1 FE_PHC3871_n5506 (.Z(FE_PHN3871_n5506), 
	.A(n5506));
   BUF_X8 FE_PHC3869_U769_Z_0 (.Z(FE_PHN3869_U769_Z_0), 
	.A(U769_Z_0));
   BUF_X8 FE_PHC3868_U503_Z_0 (.Z(FE_PHN3868_U503_Z_0), 
	.A(U503_Z_0));
   CLKBUF_X1 FE_PHC3866_n5265 (.Z(FE_PHN3866_n5265), 
	.A(n5265));
   CLKBUF_X3 FE_PHC3865_U345_Z_0 (.Z(FE_PHN3865_U345_Z_0), 
	.A(U345_Z_0));
   BUF_X8 FE_PHC3864_U428_Z_0 (.Z(FE_PHN3864_U428_Z_0), 
	.A(U428_Z_0));
   BUF_X8 FE_PHC3863_U646_Z_0 (.Z(FE_PHN3863_U646_Z_0), 
	.A(U646_Z_0));
   CLKBUF_X2 FE_PHC3862_U711_Z_0 (.Z(FE_PHN3862_U711_Z_0), 
	.A(U711_Z_0));
   BUF_X8 FE_PHC3857_U363_Z_0 (.Z(FE_PHN3857_U363_Z_0), 
	.A(FE_PHN2871_U363_Z_0));
   BUF_X8 FE_PHC3856_U677_Z_0 (.Z(FE_PHN3856_U677_Z_0), 
	.A(U677_Z_0));
   CLKBUF_X1 FE_PHC3853_U628_Z_0 (.Z(FE_PHN3853_U628_Z_0), 
	.A(U628_Z_0));
   BUF_X8 FE_PHC3851_U504_Z_0 (.Z(FE_PHN3851_U504_Z_0), 
	.A(U504_Z_0));
   BUF_X8 FE_PHC3847_U471_Z_0 (.Z(FE_PHN3847_U471_Z_0), 
	.A(U471_Z_0));
   BUF_X8 FE_PHC3845_U800_Z_0 (.Z(FE_PHN3845_U800_Z_0), 
	.A(FE_PHN2867_U800_Z_0));
   BUF_X8 FE_PHC3843_U619_Z_0 (.Z(FE_PHN3843_U619_Z_0), 
	.A(U619_Z_0));
   CLKBUF_X2 FE_PHC3842_U263_Z_0 (.Z(FE_PHN3842_U263_Z_0), 
	.A(U263_Z_0));
   CLKBUF_X2 FE_PHC3839_U745_Z_0 (.Z(FE_PHN3839_U745_Z_0), 
	.A(U745_Z_0));
   BUF_X16 FE_PHC3836_U612_Z_0 (.Z(FE_PHN3836_U612_Z_0), 
	.A(U612_Z_0));
   BUF_X8 FE_PHC3828_n5168 (.Z(FE_PHN3828_n5168), 
	.A(n5168));
   BUF_X8 FE_PHC3823_U585_Z_0 (.Z(FE_PHN3823_U585_Z_0), 
	.A(U585_Z_0));
   BUF_X8 FE_PHC3821_U481_Z_0 (.Z(FE_PHN3821_U481_Z_0), 
	.A(U481_Z_0));
   BUF_X16 FE_PHC3814_U425_Z_0 (.Z(FE_PHN3814_U425_Z_0), 
	.A(FE_PHN2868_U425_Z_0));
   BUF_X8 FE_PHC3811_U513_Z_0 (.Z(FE_PHN3811_U513_Z_0), 
	.A(FE_PHN2862_U513_Z_0));
   BUF_X16 FE_PHC3808_n270 (.Z(FE_PHN3808_n270), 
	.A(n270));
   BUF_X8 FE_PHC3806_U663_Z_0 (.Z(FE_PHN3806_U663_Z_0), 
	.A(U663_Z_0));
   CLKBUF_X2 FE_PHC3803_U748_Z_0 (.Z(FE_PHN3803_U748_Z_0), 
	.A(U748_Z_0));
   BUF_X16 FE_PHC3802_U490_Z_0 (.Z(FE_PHN3802_U490_Z_0), 
	.A(U490_Z_0));
   CLKBUF_X3 FE_PHC3799_U335_Z_0 (.Z(FE_PHN3799_U335_Z_0), 
	.A(U335_Z_0));
   BUF_X8 FE_PHC3798_U454_Z_0 (.Z(FE_PHN3798_U454_Z_0), 
	.A(U454_Z_0));
   BUF_X16 FE_PHC3797_U391_Z_0 (.Z(FE_PHN3797_U391_Z_0), 
	.A(U391_Z_0));
   BUF_X16 FE_PHC3796_U754_Z_0 (.Z(FE_PHN3796_U754_Z_0), 
	.A(U754_Z_0));
   BUF_X8 FE_PHC3793_n4982 (.Z(FE_PHN3793_n4982), 
	.A(n4982));
   BUF_X8 FE_PHC3787_U242_Z_0 (.Z(FE_PHN3787_U242_Z_0), 
	.A(U242_Z_0));
   BUF_X8 FE_PHC3785_U667_Z_0 (.Z(FE_PHN3785_U667_Z_0), 
	.A(FE_PHN2860_U667_Z_0));
   CLKBUF_X3 FE_PHC3784_U651_Z_0 (.Z(FE_PHN3784_U651_Z_0), 
	.A(U651_Z_0));
   CLKBUF_X2 FE_PHC3782_U728_Z_0 (.Z(FE_PHN3782_U728_Z_0), 
	.A(U728_Z_0));
   BUF_X8 FE_PHC3780_n5134 (.Z(FE_PHN3780_n5134), 
	.A(n5134));
   BUF_X16 FE_PHC3779_n286 (.Z(FE_PHN3779_n286), 
	.A(n286));
   CLKBUF_X2 FE_PHC3778_U743_Z_0 (.Z(FE_PHN3778_U743_Z_0), 
	.A(U743_Z_0));
   BUF_X8 FE_PHC3775_U500_Z_0 (.Z(FE_PHN3775_U500_Z_0), 
	.A(U500_Z_0));
   CLKBUF_X2 FE_PHC3774_U708_Z_0 (.Z(FE_PHN3774_U708_Z_0), 
	.A(U708_Z_0));
   BUF_X16 FE_PHC3769_U407_Z_0 (.Z(FE_PHN3769_U407_Z_0), 
	.A(FE_PHN2846_U407_Z_0));
   BUF_X8 FE_PHC3765_U683_Z_0 (.Z(FE_PHN3765_U683_Z_0), 
	.A(U683_Z_0));
   BUF_X16 FE_PHC3764_n5004 (.Z(FE_PHN3764_n5004), 
	.A(n5004));
   BUF_X16 FE_PHC3763_U233_Z_0 (.Z(FE_PHN3763_U233_Z_0), 
	.A(U233_Z_0));
   BUF_X8 FE_PHC3762_U496_Z_0 (.Z(FE_PHN3762_U496_Z_0), 
	.A(U496_Z_0));
   BUF_X16 FE_PHC3755_n8706 (.Z(FE_PHN3755_n8706), 
	.A(FE_PHN1566_n8706));
   BUF_X8 FE_PHC3753_U445_Z_0 (.Z(FE_PHN3753_U445_Z_0), 
	.A(U445_Z_0));
   BUF_X16 FE_PHC3744_U610_Z_0 (.Z(FE_PHN3744_U610_Z_0), 
	.A(FE_PHN2844_U610_Z_0));
   BUF_X16 FE_PHC3735_n284 (.Z(FE_PHN3735_n284), 
	.A(n284));
   BUF_X16 FE_PHC3733_U463_Z_0 (.Z(FE_PHN3733_U463_Z_0), 
	.A(FE_PHN2842_U463_Z_0));
   BUF_X16 FE_PHC3730_U497_Z_0 (.Z(FE_PHN3730_U497_Z_0), 
	.A(FE_PHN2855_U497_Z_0));
   BUF_X16 FE_PHC3726_n5193 (.Z(FE_PHN3726_n5193), 
	.A(n5193));
   BUF_X16 FE_PHC3725_U594_Z_0 (.Z(FE_PHN3725_U594_Z_0), 
	.A(FE_PHN2355_U594_Z_0));
   BUF_X16 FE_PHC3718_U680_Z_0 (.Z(FE_PHN3718_U680_Z_0), 
	.A(U680_Z_0));
   BUF_X16 FE_PHC3717_n278 (.Z(FE_PHN3717_n278), 
	.A(n278));
   BUF_X8 FE_PHC3699_n5056 (.Z(FE_PHN3699_n5056), 
	.A(n5056));
   BUF_X16 FE_PHC3690_n8698 (.Z(FE_PHN3690_n8698), 
	.A(FE_PHN1565_n8698));
   BUF_X8 FE_PHC3682_U634_Z_0 (.Z(FE_PHN3682_U634_Z_0), 
	.A(U634_Z_0));
   BUF_X16 FE_PHC3681_n5302 (.Z(FE_PHN3681_n5302), 
	.A(n5302));
   BUF_X8 FE_PHC3663_U656_Z_0 (.Z(FE_PHN3663_U656_Z_0), 
	.A(U656_Z_0));
   BUF_X8 FE_PHC3662_n276 (.Z(FE_PHN3662_n276), 
	.A(n276));
   BUF_X16 FE_PHC3661_n4852 (.Z(FE_PHN3661_n4852), 
	.A(n4852));
   BUF_X16 FE_PHC3654_n5733 (.Z(FE_PHN3654_n5733), 
	.A(FE_PHN1142_n5733));
   BUF_X16 FE_PHC3648_n5594 (.Z(FE_PHN3648_n5594), 
	.A(n5594));
   BUF_X16 FE_PHC3647_U493_Z_0 (.Z(FE_PHN3647_U493_Z_0), 
	.A(FE_PHN2838_U493_Z_0));
   BUF_X16 FE_PHC3642_n5179 (.Z(FE_PHN3642_n5179), 
	.A(n5179));
   BUF_X16 FE_PHC3641_n282 (.Z(FE_PHN3641_n282), 
	.A(n282));
   BUF_X16 FE_PHC3639_n5735 (.Z(FE_PHN3639_n5735), 
	.A(FE_PHN1255_n5735));
   BUF_X16 FE_PHC3637_n5429 (.Z(FE_PHN3637_n5429), 
	.A(n5429));
   BUF_X2 FE_PHC3636_U341_Z_0 (.Z(FE_PHN3636_U341_Z_0), 
	.A(U341_Z_0));
   BUF_X16 FE_PHC3635_n5645 (.Z(FE_PHN3635_n5645), 
	.A(n5645));
   BUF_X16 FE_PHC3634_n5475 (.Z(FE_PHN3634_n5475), 
	.A(n5475));
   BUF_X16 FE_PHC3633_n4989 (.Z(FE_PHN3633_n4989), 
	.A(n4989));
   BUF_X16 FE_PHC3631_n294 (.Z(FE_PHN3631_n294), 
	.A(n294));
   BUF_X16 FE_PHC3630_n5194 (.Z(FE_PHN3630_n5194), 
	.A(n5194));
   BUF_X16 FE_PHC3629_n5400 (.Z(FE_PHN3629_n5400), 
	.A(n5400));
   BUF_X16 FE_PHC3627_n5147 (.Z(FE_PHN3627_n5147), 
	.A(n5147));
   BUF_X16 FE_PHC3626_n5446 (.Z(FE_PHN3626_n5446), 
	.A(n5446));
   BUF_X16 FE_PHC3625_n5732 (.Z(FE_PHN3625_n5732), 
	.A(n5732));
   BUF_X16 FE_PHC3624_n4992 (.Z(FE_PHN3624_n4992), 
	.A(n4992));
   BUF_X16 FE_PHC3623_n5058 (.Z(FE_PHN3623_n5058), 
	.A(n5058));
   BUF_X16 FE_PHC3622_n5416 (.Z(FE_PHN3622_n5416), 
	.A(n5416));
   BUF_X16 FE_PHC3621_n5499 (.Z(FE_PHN3621_n5499), 
	.A(n5499));
   BUF_X16 FE_PHC3620_n4848 (.Z(FE_PHN3620_n4848), 
	.A(n4848));
   BUF_X8 FE_PHC3617_n5586 (.Z(FE_PHN3617_n5586), 
	.A(n5586));
   BUF_X32 FE_PHC3616_n4853 (.Z(FE_PHN3616_n4853), 
	.A(n4853));
   BUF_X16 FE_PHC3615_n4746 (.Z(FE_PHN3615_n4746), 
	.A(n4746));
   BUF_X16 FE_PHC3612_n5731 (.Z(FE_PHN3612_n5731), 
	.A(n5731));
   BUF_X32 FE_PHC3611_n288 (.Z(FE_PHN3611_n288), 
	.A(n288));
   BUF_X32 FE_PHC3610_n5725 (.Z(FE_PHN3610_n5725), 
	.A(n5725));
   BUF_X16 FE_PHC3609_n5327 (.Z(FE_PHN3609_n5327), 
	.A(n5327));
   BUF_X32 FE_PHC3608_n5784 (.Z(FE_PHN3608_n5784), 
	.A(n5784));
   BUF_X16 FE_PHC3606_U98_Z_0 (.Z(FE_PHN3606_U98_Z_0), 
	.A(FE_PHN1633_U98_Z_0));
   BUF_X16 FE_PHC3605_n5402 (.Z(FE_PHN3605_n5402), 
	.A(n5402));
   BUF_X32 FE_PHC3604_n5730 (.Z(FE_PHN3604_n5730), 
	.A(n5730));
   BUF_X16 FE_PHC3603_n5583 (.Z(FE_PHN3603_n5583), 
	.A(n5583));
   BUF_X16 FE_PHC3602_n4829 (.Z(FE_PHN3602_n4829), 
	.A(n4829));
   BUF_X16 FE_PHC3601_n5094 (.Z(FE_PHN3601_n5094), 
	.A(n5094));
   BUF_X32 FE_PHC3599_n5377 (.Z(FE_PHN3599_n5377), 
	.A(n5377));
   BUF_X32 FE_PHC3598_n5500 (.Z(FE_PHN3598_n5500), 
	.A(n5500));
   BUF_X32 FE_PHC3597_U721_Z_0 (.Z(FE_PHN3597_U721_Z_0), 
	.A(FE_PHN2816_U721_Z_0));
   BUF_X32 FE_PHC3596_n5145 (.Z(FE_PHN3596_n5145), 
	.A(n5145));
   BUF_X32 FE_PHC3595_n5720 (.Z(FE_PHN3595_n5720), 
	.A(n5720));
   BUF_X16 FE_PHC3594_n5330 (.Z(FE_PHN3594_n5330), 
	.A(n5330));
   BUF_X32 FE_PHC3593_n5269 (.Z(FE_PHN3593_n5269), 
	.A(n5269));
   BUF_X16 FE_PHC3592_n5714 (.Z(FE_PHN3592_n5714), 
	.A(n5714));
   BUF_X32 FE_PHC3591_n5726 (.Z(FE_PHN3591_n5726), 
	.A(n5726));
   BUF_X32 FE_PHC3590_n5588 (.Z(FE_PHN3590_n5588), 
	.A(n5588));
   BUF_X32 FE_PHC3589_n5059 (.Z(FE_PHN3589_n5059), 
	.A(n5059));
   BUF_X32 FE_PHC3587_n5359 (.Z(FE_PHN3587_n5359), 
	.A(n5359));
   BUF_X32 FE_PHC3586_n5293 (.Z(FE_PHN3586_n5293), 
	.A(n5293));
   BUF_X32 FE_PHC3585_n5734 (.Z(FE_PHN3585_n5734), 
	.A(FE_PHN1139_n5734));
   BUF_X32 FE_PHC3584_n4990 (.Z(FE_PHN3584_n4990), 
	.A(n4990));
   BUF_X16 FE_PHC3583_n4980 (.Z(FE_PHN3583_n4980), 
	.A(n4980));
   BUF_X32 FE_PHC3582_U453_Z_0 (.Z(FE_PHN3582_U453_Z_0), 
	.A(FE_PHN2800_U453_Z_0));
   BUF_X32 FE_PHC3581_n5032 (.Z(FE_PHN3581_n5032), 
	.A(n5032));
   BUF_X16 FE_PHC3580_n5148 (.Z(FE_PHN3580_n5148), 
	.A(n5148));
   BUF_X32 FE_PHC3578_n5406 (.Z(FE_PHN3578_n5406), 
	.A(n5406));
   BUF_X32 FE_PHC3577_n5295 (.Z(FE_PHN3577_n5295), 
	.A(n5295));
   BUF_X32 FE_PHC3576_U97_Z_0 (.Z(FE_PHN3576_U97_Z_0), 
	.A(FE_PHN1632_U97_Z_0));
   BUF_X32 FE_PHC3574_n5587 (.Z(FE_PHN3574_n5587), 
	.A(n5587));
   BUF_X16 FE_PHC3573_U320_Z_0 (.Z(FE_PHN3573_U320_Z_0), 
	.A(FE_PHN4999_U320_Z_0));
   BUF_X32 FE_PHC3572_n5590 (.Z(FE_PHN3572_n5590), 
	.A(n5590));
   BUF_X16 FE_PHC3571_n5223 (.Z(FE_PHN3571_n5223), 
	.A(n5223));
   BUF_X32 FE_PHC3570_n5222 (.Z(FE_PHN3570_n5222), 
	.A(n5222));
   BUF_X32 FE_PHC3569_n5282 (.Z(FE_PHN3569_n5282), 
	.A(n5282));
   BUF_X32 FE_PHC3568_n5556 (.Z(FE_PHN3568_n5556), 
	.A(n5556));
   BUF_X32 FE_PHC3567_n5342 (.Z(FE_PHN3567_n5342), 
	.A(n5342));
   BUF_X32 FE_PHC3566_n5031 (.Z(FE_PHN3566_n5031), 
	.A(n5031));
   BUF_X32 FE_PHC3565_n5404 (.Z(FE_PHN3565_n5404), 
	.A(n5404));
   BUF_X32 FE_PHC3564_n5375 (.Z(FE_PHN3564_n5375), 
	.A(n5375));
   BUF_X32 FE_PHC3563_n5482 (.Z(FE_PHN3563_n5482), 
	.A(n5482));
   BUF_X32 FE_PHC3562_n5371 (.Z(FE_PHN3562_n5371), 
	.A(n5371));
   BUF_X32 FE_PHC3561_U630_Z_0 (.Z(FE_PHN3561_U630_Z_0), 
	.A(FE_PHN1759_U630_Z_0));
   BUF_X32 FE_PHC3560_n5303 (.Z(FE_PHN3560_n5303), 
	.A(n5303));
   BUF_X32 FE_PHC3559_n5373 (.Z(FE_PHN3559_n5373), 
	.A(n5373));
   BUF_X32 FE_PHC3558_n5591 (.Z(FE_PHN3558_n5591), 
	.A(n5591));
   BUF_X32 FE_PHC3557_n5274 (.Z(FE_PHN3557_n5274), 
	.A(n5274));
   BUF_X32 FE_PHC3556_n5206 (.Z(FE_PHN3556_n5206), 
	.A(n5206));
   BUF_X32 FE_PHC3555_n5281 (.Z(FE_PHN3555_n5281), 
	.A(n5281));
   BUF_X32 FE_PHC3554_n5060 (.Z(FE_PHN3554_n5060), 
	.A(n5060));
   BUF_X32 FE_PHC3553_n5647 (.Z(FE_PHN3553_n5647), 
	.A(n5647));
   BUF_X32 FE_PHC3552_U246_Z_0 (.Z(FE_PHN3552_U246_Z_0), 
	.A(FE_PHN2101_U246_Z_0));
   BUF_X32 FE_PHC3551_n5593 (.Z(FE_PHN3551_n5593), 
	.A(n5593));
   BUF_X32 FE_PHC3550_n5417 (.Z(FE_PHN3550_n5417), 
	.A(n5417));
   BUF_X32 FE_PHC3548_U627_Z_0 (.Z(FE_PHN3548_U627_Z_0), 
	.A(FE_PHN2179_U627_Z_0));
   BUF_X32 FE_PHC3547_n5728 (.Z(FE_PHN3547_n5728), 
	.A(FE_PHN1133_n5728));
   BUF_X16 FE_PHC3546_U319_Z_0 (.Z(FE_PHN3546_U319_Z_0), 
	.A(FE_PHN1751_U319_Z_0));
   BUF_X32 FE_PHC3545_U586_Z_0 (.Z(FE_PHN3545_U586_Z_0), 
	.A(FE_PHN2114_U586_Z_0));
   BUF_X32 FE_PHC3544_n5716 (.Z(FE_PHN3544_n5716), 
	.A(FE_PHN1134_n5716));
   BUF_X32 FE_PHC3542_U597_Z_0 (.Z(FE_PHN3542_U597_Z_0), 
	.A(FE_PHN2148_U597_Z_0));
   BUF_X32 FE_PHC3541_U519_Z_0 (.Z(FE_PHN3541_U519_Z_0), 
	.A(FE_PHN2105_U519_Z_0));
   BUF_X32 FE_PHC3540_U235_Z_0 (.Z(FE_PHN3540_U235_Z_0), 
	.A(FE_PHN2109_U235_Z_0));
   BUF_X16 FE_PHC3539_U321_Z_0 (.Z(FE_PHN3539_U321_Z_0), 
	.A(FE_PHN2099_U321_Z_0));
   BUF_X32 FE_PHC3538_U632_Z_0 (.Z(FE_PHN3538_U632_Z_0), 
	.A(FE_PHN2093_U632_Z_0));
   BUF_X32 FE_PHC3537_U591_Z_0 (.Z(FE_PHN3537_U591_Z_0), 
	.A(FE_PHN5170_U591_Z_0));
   BUF_X32 FE_PHC3536_n4938 (.Z(FE_PHN3536_n4938), 
	.A(FE_PHN4783_n4938));
   BUF_X16 FE_PHC3535_U247_Z_0 (.Z(FE_PHN3535_U247_Z_0), 
	.A(FE_PHN5131_U247_Z_0));
   BUF_X32 FE_PHC3534_n4924 (.Z(FE_PHN3534_n4924), 
	.A(FE_PHN5010_n4924));
   BUF_X32 FE_PHC3533_U583_Z_0 (.Z(FE_PHN3533_U583_Z_0), 
	.A(FE_PHN5104_U583_Z_0));
   BUF_X16 FE_PHC3532_U528_Z_0 (.Z(FE_PHN3532_U528_Z_0), 
	.A(FE_PHN5119_U528_Z_0));
   BUF_X32 FE_PHC3531_U595_Z_0 (.Z(FE_PHN3531_U595_Z_0), 
	.A(FE_PHN5076_U595_Z_0));
   BUF_X32 FE_PHC3530_U589_Z_0 (.Z(FE_PHN3530_U589_Z_0), 
	.A(FE_PHN5077_U589_Z_0));
   BUF_X16 FE_PHC3529_U309_Z_0 (.Z(FE_PHN3529_U309_Z_0), 
	.A(FE_PHN5025_U309_Z_0));
   BUF_X32 FE_PHC3528_U557_Z_0 (.Z(FE_PHN3528_U557_Z_0), 
	.A(FE_PHN4983_U557_Z_0));
   BUF_X16 FE_PHC3527_U305_Z_0 (.Z(FE_PHN3527_U305_Z_0), 
	.A(FE_PHN4984_U305_Z_0));
   BUF_X16 FE_PHC3526_U566_Z_0 (.Z(FE_PHN3526_U566_Z_0), 
	.A(FE_PHN4943_U566_Z_0));
   BUF_X16 FE_PHC3525_U324_Z_0 (.Z(FE_PHN3525_U324_Z_0), 
	.A(FE_PHN4960_U324_Z_0));
   BUF_X32 FE_PHC3524_U563_Z_0 (.Z(FE_PHN3524_U563_Z_0), 
	.A(FE_PHN4930_U563_Z_0));
   BUF_X16 FE_PHC3523_U318_Z_0 (.Z(FE_PHN3523_U318_Z_0), 
	.A(FE_PHN4923_U318_Z_0));
   BUF_X16 FE_PHC3522_U323_Z_0 (.Z(FE_PHN3522_U323_Z_0), 
	.A(FE_PHN4944_U323_Z_0));
   BUF_X32 FE_PHC3521_n4937 (.Z(FE_PHN3521_n4937), 
	.A(FE_PHN4779_n4937));
   BUF_X32 FE_PHC3520_n4925 (.Z(FE_PHN3520_n4925), 
	.A(FE_PHN4749_n4925));
   BUF_X32 FE_PHC3519_n4935 (.Z(FE_PHN3519_n4935), 
	.A(FE_PHN4733_n4935));
   BUF_X32 FE_PHC3518_n4936 (.Z(FE_PHN3518_n4936), 
	.A(FE_PHN4731_n4936));
   BUF_X32 FE_PHC3517_n4926 (.Z(FE_PHN3517_n4926), 
	.A(FE_PHN4730_n4926));
   BUF_X32 FE_PHC3516_n4942 (.Z(FE_PHN3516_n4942), 
	.A(FE_PHN4729_n4942));
   CLKBUF_X1 FE_PHC3512_n5510 (.Z(FE_PHN3512_n5510), 
	.A(FE_PHN1748_n5510));
   CLKBUF_X1 FE_PHC3506_U795_Z_0 (.Z(FE_PHN3506_U795_Z_0), 
	.A(FE_PHN1644_U795_Z_0));
   CLKBUF_X1 FE_PHC3502_U755_Z_0 (.Z(FE_PHN3502_U755_Z_0), 
	.A(FE_PHN1649_U755_Z_0));
   CLKBUF_X1 FE_PHC3501_n5516 (.Z(FE_PHN3501_n5516), 
	.A(n5516));
   CLKBUF_X1 FE_PHC3500_n5099 (.Z(FE_PHN3500_n5099), 
	.A(n5099));
   CLKBUF_X1 FE_PHC3497_n5792 (.Z(FE_PHN3497_n5792), 
	.A(FE_PHN4985_n5792));
   CLKBUF_X1 FE_PHC3496_n262 (.Z(FE_PHN3496_n262), 
	.A(n262));
   BUF_X8 FE_PHC3482_n5711 (.Z(FE_PHN3482_n5711), 
	.A(FE_PHN2403_n5711));
   BUF_X16 FE_PHC3478_n5793 (.Z(FE_PHN3478_n5793), 
	.A(FE_PHN2379_n5793));
   BUF_X16 FE_PHC3477_n5790 (.Z(FE_PHN3477_n5790), 
	.A(FE_PHN2348_n5790));
   BUF_X32 FE_PHC3474_n5689 (.Z(FE_PHN3474_n5689), 
	.A(FE_PHN775_n5689));
   BUF_X32 FE_PHC3472_n5826 (.Z(FE_PHN3472_n5826), 
	.A(n5826));
   BUF_X32 FE_PHC3470_n5795 (.Z(FE_PHN3470_n5795), 
	.A(n5795));
   CLKBUF_X1 FE_PHC3466_n214 (.Z(FE_PHN3466_n214), 
	.A(n214));
   CLKBUF_X1 FE_PHC3437_n5783 (.Z(FE_PHN3437_n5783), 
	.A(FE_PHN1499_n5783));
   CLKBUF_X1 FE_PHC3421_n5684 (.Z(FE_PHN3421_n5684), 
	.A(FE_PHN1577_n5684));
   CLKBUF_X1 FE_PHC3414_n5679 (.Z(FE_PHN3414_n5679), 
	.A(FE_PHN991_n5679));
   CLKBUF_X1 FE_PHC3411_n222 (.Z(FE_PHN3411_n222), 
	.A(FE_PHN2049_n222));
   CLKBUF_X1 FE_PHC3405_n5677 (.Z(FE_PHN3405_n5677), 
	.A(FE_PHN946_n5677));
   CLKBUF_X1 FE_PHC3391_n5673 (.Z(FE_PHN3391_n5673), 
	.A(FE_PHN1004_n5673));
   CLKBUF_X1 FE_PHC3387_n5655 (.Z(FE_PHN3387_n5655), 
	.A(FE_PHN705_n5655));
   CLKBUF_X1 FE_PHC3377_n5682 (.Z(FE_PHN3377_n5682), 
	.A(FE_PHN1559_n5682));
   CLKBUF_X1 FE_PHC3375_n5676 (.Z(FE_PHN3375_n5676), 
	.A(FE_PHN1159_n5676));
   CLKBUF_X1 FE_PHC3353_n5675 (.Z(FE_PHN3353_n5675), 
	.A(FE_PHN1003_n5675));
   BUF_X8 FE_PHC3290_n4923 (.Z(FE_PHN3290_n4923), 
	.A(n4923));
   BUF_X32 FE_PHC3282_n5685 (.Z(FE_PHN3282_n5685), 
	.A(FE_PHN769_n5685));
   BUF_X32 FE_PHC3278_n4934 (.Z(FE_PHN3278_n4934), 
	.A(FE_PHN1389_n4934));
   BUF_X32 FE_PHC3277_n4939 (.Z(FE_PHN3277_n4939), 
	.A(FE_PHN4735_n4939));
   BUF_X32 FE_PHC3276_n4930 (.Z(FE_PHN3276_n4930), 
	.A(FE_PHN1391_n4930));
   BUF_X32 FE_PHC3275_n4928 (.Z(FE_PHN3275_n4928), 
	.A(FE_PHN1385_n4928));
   BUF_X32 FE_PHC3274_n4933 (.Z(FE_PHN3274_n4933), 
	.A(FE_PHN1175_n4933));
   BUF_X32 FE_PHC3273_n5800 (.Z(FE_PHN3273_n5800), 
	.A(n5800));
   BUF_X16 FE_PHC3217_n5736 (.Z(FE_PHN3217_n5736), 
	.A(FE_PHN1626_n5736));
   BUF_X32 FE_PHC3211_U229_Z_0 (.Z(FE_PHN3211_U229_Z_0), 
	.A(U229_Z_0));
   CLKBUF_X1 FE_PHC3209_n5791 (.Z(FE_PHN3209_n5791), 
	.A(n5791));
   BUF_X32 FE_PHC3206_n5712 (.Z(FE_PHN3206_n5712), 
	.A(FE_PHN4737_n5712));
   BUF_X32 FE_PHC3205_n5827 (.Z(FE_PHN3205_n5827), 
	.A(n5827));
   BUF_X32 FE_PHC3204_n13813 (.Z(FE_PHN3204_n13813), 
	.A(n13813));
   BUF_X32 FE_PHC3202_n13951 (.Z(FE_PHN3202_n13951), 
	.A(n13951));
   BUF_X32 FE_PHC3201_n13870 (.Z(FE_PHN3201_n13870), 
	.A(n13870));
   BUF_X32 FE_PHC3200_n5763 (.Z(FE_PHN3200_n5763), 
	.A(FE_PHN4706_n5763));
   BUF_X32 FE_PHC3199_n5756 (.Z(FE_PHN3199_n5756), 
	.A(FE_PHN4703_n5756));
   BUF_X32 FE_PHC3198_n5767 (.Z(FE_PHN3198_n5767), 
	.A(FE_PHN4661_n5767));
   CLKBUF_X1 FE_PHC3190_n4931 (.Z(FE_PHN3190_n4931), 
	.A(FE_PHN1909_n4931));
   BUF_X16 FE_PHC3153_n5668 (.Z(FE_PHN3153_n5668), 
	.A(FE_PHN1078_n5668));
   BUF_X32 FE_PHC3143_U227_Z_0 (.Z(FE_PHN3143_U227_Z_0), 
	.A(FE_PHN4711_U227_Z_0));
   BUF_X32 FE_PHC3142_n5765 (.Z(FE_PHN3142_n5765), 
	.A(FE_PHN4682_n5765));
   BUF_X32 FE_PHC3140_n4921 (.Z(FE_PHN3140_n4921), 
	.A(n4921));
   BUF_X32 FE_PHC3139_n5755 (.Z(FE_PHN3139_n5755), 
	.A(n5755));
   BUF_X32 FE_PHC3138_n5758 (.Z(FE_PHN3138_n5758), 
	.A(n5758));
   BUF_X32 FE_PHC3137_n4910 (.Z(FE_PHN3137_n4910), 
	.A(n4910));
   BUF_X32 FE_PHC3136_n4907 (.Z(FE_PHN3136_n4907), 
	.A(n4907));
   BUF_X32 FE_PHC3135_n4914 (.Z(FE_PHN3135_n4914), 
	.A(n4914));
   BUF_X32 FE_PHC3134_n5762 (.Z(FE_PHN3134_n5762), 
	.A(FE_PHN802_n5762));
   BUF_X32 FE_PHC3133_n14432 (.Z(FE_PHN3133_n14432), 
	.A(FE_PHN4694_n14432));
   BUF_X16 FE_PHC3103_n4847 (.Z(FE_PHN3103_n4847), 
	.A(n4847));
   BUF_X32 FE_PHC3102_n5237 (.Z(FE_PHN3102_n5237), 
	.A(n5237));
   BUF_X32 FE_PHC3101_n5235 (.Z(FE_PHN3101_n5235), 
	.A(n5235));
   BUF_X32 FE_PHC3100_n5573 (.Z(FE_PHN3100_n5573), 
	.A(n5573));
   BUF_X32 FE_PHC3099_n5601 (.Z(FE_PHN3099_n5601), 
	.A(n5601));
   BUF_X32 FE_PHC3098_n5238 (.Z(FE_PHN3098_n5238), 
	.A(n5238));
   BUF_X32 FE_PHC3097_n5236 (.Z(FE_PHN3097_n5236), 
	.A(n5236));
   BUF_X32 FE_PHC3094_n5761 (.Z(FE_PHN3094_n5761), 
	.A(FE_PHN4689_n5761));
   BUF_X32 FE_PHC3093_n4918 (.Z(FE_PHN3093_n4918), 
	.A(FE_PHN4690_n4918));
   BUF_X32 FE_PHC3092_n14001 (.Z(FE_PHN3092_n14001), 
	.A(n14001));
   BUF_X32 FE_PHC3091_n5768 (.Z(FE_PHN3091_n5768), 
	.A(FE_PHN4662_n5768));
   BUF_X32 FE_PHC3090_n5751 (.Z(FE_PHN3090_n5751), 
	.A(FE_PHN4710_n5751));
   BUF_X32 FE_PHC3089_n5754 (.Z(FE_PHN3089_n5754), 
	.A(FE_PHN4704_n5754));
   BUF_X32 FE_PHC3088_n5744 (.Z(FE_PHN3088_n5744), 
	.A(FE_PHN4686_n5744));
   CLKBUF_X1 FE_PHC3084_n5658 (.Z(FE_PHN3084_n5658), 
	.A(FE_PHN965_n5658));
   CLKBUF_X1 FE_PHC3078_n5729 (.Z(FE_PHN3078_n5729), 
	.A(FE_PHN1145_n5729));
   CLKBUF_X1 FE_PHC3076_U692_Z_0 (.Z(FE_PHN3076_U692_Z_0), 
	.A(U692_Z_0));
   BUF_X8 FE_PHC3074_n5798 (.Z(FE_PHN3074_n5798), 
	.A(n5798));
   BUF_X32 FE_PHC3073_n5782 (.Z(FE_PHN3073_n5782), 
	.A(FE_PHN1448_n5782));
   BUF_X16 FE_PHC3072_n5788 (.Z(FE_PHN3072_n5788), 
	.A(FE_PHN4937_n5788));
   BUF_X32 FE_PHC3071_n5717 (.Z(FE_PHN3071_n5717), 
	.A(FE_PHN1128_n5717));
   BUF_X32 FE_PHC3070_n4879 (.Z(FE_PHN3070_n4879), 
	.A(FE_PHN1377_n4879));
   BUF_X32 FE_PHC3069_n4945 (.Z(FE_PHN3069_n4945), 
	.A(n4945));
   BUF_X32 FE_PHC3068_n13795 (.Z(FE_PHN3068_n13795), 
	.A(n13795));
   BUF_X32 FE_PHC3067_n13989 (.Z(FE_PHN3067_n13989), 
	.A(n13989));
   BUF_X32 FE_PHC3066_n13963 (.Z(FE_PHN3066_n13963), 
	.A(n13963));
   BUF_X32 FE_PHC3065_n13932 (.Z(FE_PHN3065_n13932), 
	.A(n13932));
   BUF_X32 FE_PHC3064_n13835 (.Z(FE_PHN3064_n13835), 
	.A(n13835));
   BUF_X32 FE_PHC3063_n13919 (.Z(FE_PHN3063_n13919), 
	.A(n13919));
   BUF_X32 FE_PHC3061_n13894 (.Z(FE_PHN3061_n13894), 
	.A(n13894));
   BUF_X32 FE_PHC3060_n14956 (.Z(FE_PHN3060_n14956), 
	.A(n14956));
   BUF_X32 FE_PHC3059_n13907 (.Z(FE_PHN3059_n13907), 
	.A(n13907));
   BUF_X32 FE_PHC3058_n13758 (.Z(FE_PHN3058_n13758), 
	.A(n13758));
   BUF_X32 FE_PHC3057_n5769 (.Z(FE_PHN3057_n5769), 
	.A(FE_PHN4660_n5769));
   BUF_X32 FE_PHC3056_n5748 (.Z(FE_PHN3056_n5748), 
	.A(FE_PHN4657_n5748));
   CLKBUF_X1 FE_PHC3055_n166 (.Z(FE_PHN3055_n166), 
	.A(n166));
   BUF_X16 FE_PHC3050_n5713 (.Z(FE_PHN3050_n5713), 
	.A(FE_PHN1141_n5713));
   BUF_X32 FE_PHC3048_n11928 (.Z(FE_PHN3048_n11928), 
	.A(FE_PHN1502_n11928));
   BUF_X32 FE_PHC3018_IRQ_14_ (.Z(FE_PHN3018_IRQ_14_), 
	.A(FE_PHN1503_IRQ_14_));
   BUF_X32 FE_PHC3001_n4895 (.Z(FE_PHN3001_n4895), 
	.A(FE_PHN1367_n4895));
   BUF_X32 FE_PHC3000_n419 (.Z(FE_PHN3000_n419), 
	.A(FE_PHN4723_n419));
   BUF_X32 FE_PHC2995_IRQ_8_ (.Z(FE_PHN2995_IRQ_8_), 
	.A(FE_PHN1366_IRQ_8_));
   BUF_X32 FE_PHC2994_IRQ_11_ (.Z(FE_PHN2994_IRQ_11_), 
	.A(FE_PHN1351_IRQ_11_));
   BUF_X32 FE_PHC2993_IRQ_13_ (.Z(FE_PHN2993_IRQ_13_), 
	.A(FE_PHN1359_IRQ_13_));
   BUF_X32 FE_PHC2992_IRQ_2_ (.Z(FE_PHN2992_IRQ_2_), 
	.A(FE_PHN1349_IRQ_2_));
   BUF_X32 FE_PHC2991_IRQ_3_ (.Z(FE_PHN2991_IRQ_3_), 
	.A(FE_PHN1345_IRQ_3_));
   BUF_X32 FE_PHC2990_IRQ_7_ (.Z(FE_PHN2990_IRQ_7_), 
	.A(FE_PHN1361_IRQ_7_));
   BUF_X32 FE_PHC2989_IRQ_10_ (.Z(FE_PHN2989_IRQ_10_), 
	.A(FE_PHN1365_IRQ_10_));
   BUF_X32 FE_PHC2988_IRQ_9_ (.Z(FE_PHN2988_IRQ_9_), 
	.A(FE_PHN1346_IRQ_9_));
   BUF_X32 FE_PHC2987_IRQ_6_ (.Z(FE_PHN2987_IRQ_6_), 
	.A(FE_PHN1353_IRQ_6_));
   BUF_X32 FE_PHC2986_IRQ_4_ (.Z(FE_PHN2986_IRQ_4_), 
	.A(FE_PHN1363_IRQ_4_));
   BUF_X32 FE_PHC2985_IRQ_0_ (.Z(FE_PHN2985_IRQ_0_), 
	.A(FE_PHN1355_IRQ_0_));
   BUF_X32 FE_PHC2984_IRQ_5_ (.Z(FE_PHN2984_IRQ_5_), 
	.A(FE_PHN1357_IRQ_5_));
   BUF_X32 FE_PHC2983_IRQ_1_ (.Z(FE_PHN2983_IRQ_1_), 
	.A(FE_PHN1360_IRQ_1_));
   BUF_X32 FE_PHC2982_NMI (.Z(FE_PHN2982_NMI), 
	.A(FE_PHN1347_NMI));
   BUF_X32 FE_PHC2981_n5760 (.Z(FE_PHN2981_n5760), 
	.A(FE_PHN4726_n5760));
   BUF_X32 FE_PHC2980_IRQ_15_ (.Z(FE_PHN2980_IRQ_15_), 
	.A(FE_PHN1350_IRQ_15_));
   BUF_X32 FE_PHC2976_n5656 (.Z(FE_PHN2976_n5656), 
	.A(FE_PHN856_n5656));
   BUF_X32 FE_PHC2974_n5757 (.Z(FE_PHN2974_n5757), 
	.A(FE_PHN803_n5757));
   BUF_X32 FE_PHC2973_n4908 (.Z(FE_PHN2973_n4908), 
	.A(n4908));
   BUF_X32 FE_PHC2972_n5759 (.Z(FE_PHN2972_n5759), 
	.A(FE_PHN753_n5759));
   BUF_X32 FE_PHC2970_n1444 (.Z(FE_PHN2970_n1444), 
	.A(FE_PHN1164_n1444));
   BUF_X32 FE_PHC2969_n4917 (.Z(FE_PHN2969_n4917), 
	.A(FE_PHN4692_n4917));
   BUF_X32 FE_PHC2968_n4919 (.Z(FE_PHN2968_n4919), 
	.A(FE_PHN4691_n4919));
   BUF_X32 FE_PHC2967_n4920 (.Z(FE_PHN2967_n4920), 
	.A(FE_PHN4652_n4920));
   BUF_X32 FE_PHC2966_n5766 (.Z(FE_PHN2966_n5766), 
	.A(FE_PHN4684_n5766));
   BUF_X32 FE_PHC2965_n5750 (.Z(FE_PHN2965_n5750), 
	.A(FE_PHN4707_n5750));
   BUF_X32 FE_PHC2955_n5741 (.Z(FE_PHN2955_n5741), 
	.A(FE_PHN4687_n5741));
   BUF_X32 FE_PHC2954_n5753 (.Z(FE_PHN2954_n5753), 
	.A(FE_PHN4685_n5753));
   BUF_X32 FE_PHC2953_n5739 (.Z(FE_PHN2953_n5739), 
	.A(FE_PHN4683_n5739));
   BUF_X32 FE_PHC2952_n5740 (.Z(FE_PHN2952_n5740), 
	.A(FE_PHN4656_n5740));
   BUF_X32 FE_PHC2951_n4916 (.Z(FE_PHN2951_n4916), 
	.A(n4916));
   BUF_X32 FE_PHC2948_n5752 (.Z(FE_PHN2948_n5752), 
	.A(FE_PHN4709_n5752));
   BUF_X32 FE_PHC2947_n4911 (.Z(FE_PHN2947_n4911), 
	.A(n4911));
   BUF_X32 FE_PHC2946_n4913 (.Z(FE_PHN2946_n4913), 
	.A(n4913));
   BUF_X32 FE_PHC2945_n4906 (.Z(FE_PHN2945_n4906), 
	.A(n4906));
   BUF_X32 FE_PHC2944_n4909 (.Z(FE_PHN2944_n4909), 
	.A(FE_PHN4655_n4909));
   BUF_X32 FE_PHC2943_n4912 (.Z(FE_PHN2943_n4912), 
	.A(FE_PHN4654_n4912));
   BUF_X32 FE_PHC2939_n4915 (.Z(FE_PHN2939_n4915), 
	.A(FE_PHN4688_n4915));
   BUF_X32 FE_PHC2936_n5746 (.Z(FE_PHN2936_n5746), 
	.A(FE_PHN4708_n5746));
   BUF_X32 FE_PHC2935_n5745 (.Z(FE_PHN2935_n5745), 
	.A(FE_PHN4681_n5745));
   CLKBUF_X1 FE_PHC2928_n1145 (.Z(FE_PHN2928_n1145), 
	.A(FE_PHN756_n1145));
   CLKBUF_X1 FE_PHC2927_n5692 (.Z(FE_PHN2927_n5692), 
	.A(FE_PHN732_n5692));
   BUF_X32 FE_PHC2926_n5683 (.Z(FE_PHN2926_n5683), 
	.A(FE_PHN4813_n5683));
   BUF_X32 FE_PHC2922_n5747 (.Z(FE_PHN2922_n5747), 
	.A(FE_PHN4658_n5747));
   BUF_X32 FE_PHC2921_n5749 (.Z(FE_PHN2921_n5749), 
	.A(FE_PHN4680_n5749));
   BUF_X32 FE_PHC2920_n5743 (.Z(FE_PHN2920_n5743), 
	.A(FE_PHN4659_n5743));
   BUF_X32 FE_PHC2918_n5742 (.Z(FE_PHN2918_n5742), 
	.A(FE_PHN4679_n5742));
   BUF_X16 FE_PHC2916_n171 (.Z(FE_PHN2916_n171), 
	.A(FE_PHN702_n171));
   BUF_X32 FE_PHC2912_n17127 (.Z(FE_PHN2912_n17127), 
	.A(n17127));
   BUF_X32 FE_PHC2911_n17126 (.Z(FE_PHN2911_n17126), 
	.A(n17126));
   CLKBUF_X1 FE_PHC2903_n5707 (.Z(FE_PHN2903_n5707), 
	.A(n5707));
   CLKBUF_X1 FE_PHC2902_n5703 (.Z(FE_PHN2902_n5703), 
	.A(n5703));
   CLKBUF_X1 FE_PHC2901_n5706 (.Z(FE_PHN2901_n5706), 
	.A(n5706));
   CLKBUF_X1 FE_PHC2900_n5702 (.Z(FE_PHN2900_n5702), 
	.A(n5702));
   CLKBUF_X1 FE_PHC2899_n5799 (.Z(FE_PHN2899_n5799), 
	.A(n5799));
   BUF_X16 FE_PHC2898_n5710 (.Z(FE_PHN2898_n5710), 
	.A(n5710));
   BUF_X16 FE_PHC2897_U763_Z_0 (.Z(FE_PHN2897_U763_Z_0), 
	.A(U763_Z_0));
   BUF_X32 FE_PHC2896_U762_Z_0 (.Z(FE_PHN2896_U762_Z_0), 
	.A(FE_PHN4615_U762_Z_0));
   BUF_X16 FE_PHC2895_U774_Z_0 (.Z(FE_PHN2895_U774_Z_0), 
	.A(U774_Z_0));
   BUF_X32 FE_PHC2894_U781_Z_0 (.Z(FE_PHN2894_U781_Z_0), 
	.A(FE_PHN4596_U781_Z_0));
   BUF_X32 FE_PHC2893_U789_Z_0 (.Z(FE_PHN2893_U789_Z_0), 
	.A(FE_PHN4597_U789_Z_0));
   BUF_X32 FE_PHC2892_n5704 (.Z(FE_PHN2892_n5704), 
	.A(FE_PHN4588_n5704));
   BUF_X32 FE_PHC2891_n5651 (.Z(FE_PHN2891_n5651), 
	.A(FE_PHN4583_n5651));
   BUF_X32 FE_PHC2890_U791_Z_0 (.Z(FE_PHN2890_U791_Z_0), 
	.A(U791_Z_0));
   BUF_X32 FE_PHC2889_n4862 (.Z(FE_PHN2889_n4862), 
	.A(FE_PHN4575_n4862));
   BUF_X32 FE_PHC2888_n5705 (.Z(FE_PHN2888_n5705), 
	.A(FE_PHN4579_n5705));
   BUF_X32 FE_PHC2887_U771_Z_0 (.Z(FE_PHN2887_U771_Z_0), 
	.A(FE_PHN4566_U771_Z_0));
   BUF_X32 FE_PHC2886_U782_Z_0 (.Z(FE_PHN2886_U782_Z_0), 
	.A(FE_PHN4576_U782_Z_0));
   BUF_X32 FE_PHC2885_U783_Z_0 (.Z(FE_PHN2885_U783_Z_0), 
	.A(FE_PHN4572_U783_Z_0));
   BUF_X32 FE_PHC2884_U772_Z_0 (.Z(FE_PHN2884_U772_Z_0), 
	.A(FE_PHN4555_U772_Z_0));
   BUF_X16 FE_PHC2883_U353_Z_0 (.Z(FE_PHN2883_U353_Z_0), 
	.A(U353_Z_0));
   BUF_X32 FE_PHC2882_U775_Z_0 (.Z(FE_PHN2882_U775_Z_0), 
	.A(FE_PHN4478_U775_Z_0));
   BUF_X32 FE_PHC2881_U788_Z_0 (.Z(FE_PHN2881_U788_Z_0), 
	.A(FE_PHN4526_U788_Z_0));
   BUF_X16 FE_PHC2879_U441_Z_0 (.Z(FE_PHN2879_U441_Z_0), 
	.A(U441_Z_0));
   BUF_X32 FE_PHC2878_U787_Z_0 (.Z(FE_PHN2878_U787_Z_0), 
	.A(FE_PHN4479_U787_Z_0));
   BUF_X32 FE_PHC2877_U786_Z_0 (.Z(FE_PHN2877_U786_Z_0), 
	.A(FE_PHN4454_U786_Z_0));
   BUF_X32 FE_PHC2875_U770_Z_0 (.Z(FE_PHN2875_U770_Z_0), 
	.A(FE_PHN4512_U770_Z_0));
   BUF_X32 FE_PHC2874_U764_Z_0 (.Z(FE_PHN2874_U764_Z_0), 
	.A(U764_Z_0));
   BUF_X32 FE_PHC2873_U459_Z_0 (.Z(FE_PHN2873_U459_Z_0), 
	.A(FE_PHN4453_U459_Z_0));
   BUF_X32 FE_PHC2872_U261_Z_0 (.Z(FE_PHN2872_U261_Z_0), 
	.A(FE_PHN4297_U261_Z_0));
   BUF_X16 FE_PHC2871_U363_Z_0 (.Z(FE_PHN2871_U363_Z_0), 
	.A(U363_Z_0));
   BUF_X32 FE_PHC2870_U780_Z_0 (.Z(FE_PHN2870_U780_Z_0), 
	.A(FE_PHN4322_U780_Z_0));
   BUF_X16 FE_PHC2869_U279_Z_0 (.Z(FE_PHN2869_U279_Z_0), 
	.A(FE_PHN4326_U279_Z_0));
   BUF_X16 FE_PHC2868_U425_Z_0 (.Z(FE_PHN2868_U425_Z_0), 
	.A(U425_Z_0));
   BUF_X16 FE_PHC2867_U800_Z_0 (.Z(FE_PHN2867_U800_Z_0), 
	.A(U800_Z_0));
   BUF_X32 FE_PHC2866_U479_Z_0 (.Z(FE_PHN2866_U479_Z_0), 
	.A(FE_PHN4272_U479_Z_0));
   BUF_X32 FE_PHC2865_n4854 (.Z(FE_PHN2865_n4854), 
	.A(FE_PHN4289_n4854));
   BUF_X32 FE_PHC2864_U429_Z_0 (.Z(FE_PHN2864_U429_Z_0), 
	.A(FE_PHN4269_U429_Z_0));
   BUF_X32 FE_PHC2863_U606_Z_0 (.Z(FE_PHN2863_U606_Z_0), 
	.A(FE_PHN4982_U606_Z_0));
   BUF_X16 FE_PHC2862_U513_Z_0 (.Z(FE_PHN2862_U513_Z_0), 
	.A(U513_Z_0));
   BUF_X16 FE_PHC2861_U275_Z_0 (.Z(FE_PHN2861_U275_Z_0), 
	.A(FE_PHN5084_U275_Z_0));
   BUF_X16 FE_PHC2860_U667_Z_0 (.Z(FE_PHN2860_U667_Z_0), 
	.A(U667_Z_0));
   BUF_X32 FE_PHC2859_U726_Z_0 (.Z(FE_PHN2859_U726_Z_0), 
	.A(FE_PHN4920_U726_Z_0));
   BUF_X32 FE_PHC2858_U359_Z_0 (.Z(FE_PHN2858_U359_Z_0), 
	.A(FE_PHN5091_U359_Z_0));
   BUF_X32 FE_PHC2857_U766_Z_0 (.Z(FE_PHN2857_U766_Z_0), 
	.A(U766_Z_0));
   BUF_X16 FE_PHC2856_U395_Z_0 (.Z(FE_PHN2856_U395_Z_0), 
	.A(FE_PHN4927_U395_Z_0));
   BUF_X16 FE_PHC2855_U497_Z_0 (.Z(FE_PHN2855_U497_Z_0), 
	.A(U497_Z_0));
   BUF_X32 FE_PHC2854_U509_Z_0 (.Z(FE_PHN2854_U509_Z_0), 
	.A(FE_PHN4270_U509_Z_0));
   BUF_X32 FE_PHC2853_U506_Z_0 (.Z(FE_PHN2853_U506_Z_0), 
	.A(FE_PHN4932_U506_Z_0));
   BUF_X32 FE_PHC2852_U660_Z_0 (.Z(FE_PHN2852_U660_Z_0), 
	.A(FE_PHN4882_U660_Z_0));
   BUF_X32 FE_PHC2851_U448_Z_0 (.Z(FE_PHN2851_U448_Z_0), 
	.A(FE_PHN3989_U448_Z_0));
   BUF_X32 FE_PHC2849_U761_Z_0 (.Z(FE_PHN2849_U761_Z_0), 
	.A(FE_PHN5113_U761_Z_0));
   BUF_X32 FE_PHC2848_U411_Z_0 (.Z(FE_PHN2848_U411_Z_0), 
	.A(FE_PHN4958_U411_Z_0));
   BUF_X32 FE_PHC2847_U475_Z_0 (.Z(FE_PHN2847_U475_Z_0), 
	.A(FE_PHN4869_U475_Z_0));
   BUF_X16 FE_PHC2846_U407_Z_0 (.Z(FE_PHN2846_U407_Z_0), 
	.A(U407_Z_0));
   BUF_X32 FE_PHC2845_U673_Z_0 (.Z(FE_PHN2845_U673_Z_0), 
	.A(FE_PHN4921_U673_Z_0));
   BUF_X16 FE_PHC2844_U610_Z_0 (.Z(FE_PHN2844_U610_Z_0), 
	.A(U610_Z_0));
   BUF_X16 FE_PHC2843_U291_Z_0 (.Z(FE_PHN2843_U291_Z_0), 
	.A(FE_PHN4862_U291_Z_0));
   BUF_X16 FE_PHC2842_U463_Z_0 (.Z(FE_PHN2842_U463_Z_0), 
	.A(U463_Z_0));
   BUF_X32 FE_PHC2841_U777_Z_0 (.Z(FE_PHN2841_U777_Z_0), 
	.A(FE_PHN4264_U777_Z_0));
   BUF_X16 FE_PHC2839_U801_Z_0 (.Z(FE_PHN2839_U801_Z_0), 
	.A(U801_Z_0));
   BUF_X16 FE_PHC2838_U493_Z_0 (.Z(FE_PHN2838_U493_Z_0), 
	.A(U493_Z_0));
   BUF_X32 FE_PHC2837_U785_Z_0 (.Z(FE_PHN2837_U785_Z_0), 
	.A(FE_PHN4298_U785_Z_0));
   BUF_X32 FE_PHC2836_U257_Z_0 (.Z(FE_PHN2836_U257_Z_0), 
	.A(FE_PHN4047_U257_Z_0));
   BUF_X32 FE_PHC2835_U466_Z_0 (.Z(FE_PHN2835_U466_Z_0), 
	.A(FE_PHN4863_U466_Z_0));
   BUF_X16 FE_PHC2834_U712_Z_0 (.Z(FE_PHN2834_U712_Z_0), 
	.A(FE_PHN4844_U712_Z_0));
   BUF_X16 FE_PHC2833_U727_Z_0 (.Z(FE_PHN2833_U727_Z_0), 
	.A(U727_Z_0));
   BUF_X32 FE_PHC2832_U784_Z_0 (.Z(FE_PHN2832_U784_Z_0), 
	.A(FE_PHN5031_U784_Z_0));
   BUF_X32 FE_PHC2831_U644_Z_0 (.Z(FE_PHN2831_U644_Z_0), 
	.A(FE_PHN5089_U644_Z_0));
   BUF_X16 FE_PHC2830_U711_Z_0 (.Z(FE_PHN2830_U711_Z_0), 
	.A(FE_PHN5080_U711_Z_0));
   BUF_X16 FE_PHC2829_U295_Z_0 (.Z(FE_PHN2829_U295_Z_0), 
	.A(FE_PHN4138_U295_Z_0));
   BUF_X16 FE_PHC2828_U386_Z_0 (.Z(FE_PHN2828_U386_Z_0), 
	.A(FE_PHN3900_U386_Z_0));
   BUF_X32 FE_PHC2827_U503_Z_0 (.Z(FE_PHN2827_U503_Z_0), 
	.A(FE_PHN5166_U503_Z_0));
   BUF_X32 FE_PHC2826_n5097 (.Z(FE_PHN2826_n5097), 
	.A(FE_PHN4586_n5097));
   BUF_X32 FE_PHC2824_U428_Z_0 (.Z(FE_PHN2824_U428_Z_0), 
	.A(FE_PHN5096_U428_Z_0));
   BUF_X16 FE_PHC2823_U263_Z_0 (.Z(FE_PHN2823_U263_Z_0), 
	.A(FE_PHN4900_U263_Z_0));
   BUF_X32 FE_PHC2822_U504_Z_0 (.Z(FE_PHN2822_U504_Z_0), 
	.A(FE_PHN4884_U504_Z_0));
   BUF_X32 FE_PHC2821_U677_Z_0 (.Z(FE_PHN2821_U677_Z_0), 
	.A(FE_PHN5049_U677_Z_0));
   BUF_X32 FE_PHC2820_U646_Z_0 (.Z(FE_PHN2820_U646_Z_0), 
	.A(FE_PHN5097_U646_Z_0));
   BUF_X32 FE_PHC2819_U471_Z_0 (.Z(FE_PHN2819_U471_Z_0), 
	.A(FE_PHN4954_U471_Z_0));
   BUF_X32 FE_PHC2818_n5650 (.Z(FE_PHN2818_n5650), 
	.A(FE_PHN3902_n5650));
   BUF_X32 FE_PHC2817_U779_Z_0 (.Z(FE_PHN2817_U779_Z_0), 
	.A(FE_PHN4860_U779_Z_0));
   BUF_X16 FE_PHC2816_U721_Z_0 (.Z(FE_PHN2816_U721_Z_0), 
	.A(U721_Z_0));
   BUF_X32 FE_PHC2815_U490_Z_0 (.Z(FE_PHN2815_U490_Z_0), 
	.A(FE_PHN3802_U490_Z_0));
   BUF_X32 FE_PHC2814_U612_Z_0 (.Z(FE_PHN2814_U612_Z_0), 
	.A(FE_PHN3836_U612_Z_0));
   BUF_X16 FE_PHC2813_U391_Z_0 (.Z(FE_PHN2813_U391_Z_0), 
	.A(FE_PHN3797_U391_Z_0));
   BUF_X32 FE_PHC2812_U683_Z_0 (.Z(FE_PHN2812_U683_Z_0), 
	.A(FE_PHN4774_U683_Z_0));
   BUF_X16 FE_PHC2811_U728_Z_0 (.Z(FE_PHN2811_U728_Z_0), 
	.A(FE_PHN4781_U728_Z_0));
   BUF_X32 FE_PHC2810_U663_Z_0 (.Z(FE_PHN2810_U663_Z_0), 
	.A(FE_PHN4891_U663_Z_0));
   BUF_X32 FE_PHC2809_U445_Z_0 (.Z(FE_PHN2809_U445_Z_0), 
	.A(FE_PHN4814_U445_Z_0));
   BUF_X16 FE_PHC2808_U651_Z_0 (.Z(FE_PHN2808_U651_Z_0), 
	.A(FE_PHN4815_U651_Z_0));
   BUF_X16 FE_PHC2807_U745_Z_0 (.Z(FE_PHN2807_U745_Z_0), 
	.A(FE_PHN4895_U745_Z_0));
   BUF_X32 FE_PHC2806_U680_Z_0 (.Z(FE_PHN2806_U680_Z_0), 
	.A(FE_PHN3718_U680_Z_0));
   BUF_X32 FE_PHC2805_U454_Z_0 (.Z(FE_PHN2805_U454_Z_0), 
	.A(FE_PHN4835_U454_Z_0));
   BUF_X16 FE_PHC2804_U743_Z_0 (.Z(FE_PHN2804_U743_Z_0), 
	.A(FE_PHN4834_U743_Z_0));
   BUF_X32 FE_PHC2803_U769_Z_0 (.Z(FE_PHN2803_U769_Z_0), 
	.A(FE_PHN5145_U769_Z_0));
   BUF_X32 FE_PHC2802_U496_Z_0 (.Z(FE_PHN2802_U496_Z_0), 
	.A(FE_PHN4788_U496_Z_0));
   BUF_X32 FE_PHC2801_n5457 (.Z(FE_PHN2801_n5457), 
	.A(FE_PHN4559_n5457));
   BUF_X16 FE_PHC2800_U453_Z_0 (.Z(FE_PHN2800_U453_Z_0), 
	.A(U453_Z_0));
   BUF_X16 FE_PHC2799_U708_Z_0 (.Z(FE_PHN2799_U708_Z_0), 
	.A(FE_PHN4810_U708_Z_0));
   BUF_X16 FE_PHC2798_U748_Z_0 (.Z(FE_PHN2798_U748_Z_0), 
	.A(FE_PHN4830_U748_Z_0));
   BUF_X32 FE_PHC2796_n5267 (.Z(FE_PHN2796_n5267), 
	.A(FE_PHN4560_n5267));
   BUF_X32 FE_PHC2795_U481_Z_0 (.Z(FE_PHN2795_U481_Z_0), 
	.A(FE_PHN4890_U481_Z_0));
   BUF_X32 FE_PHC2794_U500_Z_0 (.Z(FE_PHN2794_U500_Z_0), 
	.A(FE_PHN4865_U500_Z_0));
   BUF_X32 FE_PHC2793_U656_Z_0 (.Z(FE_PHN2793_U656_Z_0), 
	.A(FE_PHN4743_U656_Z_0));
   BUF_X32 FE_PHC2792_U634_Z_0 (.Z(FE_PHN2792_U634_Z_0), 
	.A(FE_PHN4761_U634_Z_0));
   BUF_X32 FE_PHC2791_n5297 (.Z(FE_PHN2791_n5297), 
	.A(FE_PHN4540_n5297));
   BUF_X32 FE_PHC2790_n5284 (.Z(FE_PHN2790_n5284), 
	.A(FE_PHN4549_n5284));
   BUF_X32 FE_PHC2789_n5130 (.Z(FE_PHN2789_n5130), 
	.A(FE_PHN4573_n5130));
   BUF_X32 FE_PHC2788_n5062 (.Z(FE_PHN2788_n5062), 
	.A(FE_PHN4533_n5062));
   BUF_X32 FE_PHC2787_n5603 (.Z(FE_PHN2787_n5603), 
	.A(FE_PHN4536_n5603));
   BUF_X32 FE_PHC2786_n5072 (.Z(FE_PHN2786_n5072), 
	.A(FE_PHN4534_n5072));
   BUF_X32 FE_PHC2785_n5288 (.Z(FE_PHN2785_n5288), 
	.A(FE_PHN4516_n5288));
   BUF_X32 FE_PHC2784_n5568 (.Z(FE_PHN2784_n5568), 
	.A(FE_PHN4570_n5568));
   BUF_X32 FE_PHC2783_n5622 (.Z(FE_PHN2783_n5622), 
	.A(FE_PHN4509_n5622));
   BUF_X32 FE_PHC2782_n5487 (.Z(FE_PHN2782_n5487), 
	.A(FE_PHN4523_n5487));
   BUF_X32 FE_PHC2781_n5169 (.Z(FE_PHN2781_n5169), 
	.A(FE_PHN4505_n5169));
   BUF_X32 FE_PHC2780_n5612 (.Z(FE_PHN2780_n5612), 
	.A(FE_PHN4577_n5612));
   BUF_X32 FE_PHC2779_n5604 (.Z(FE_PHN2779_n5604), 
	.A(FE_PHN4553_n5604));
   BUF_X32 FE_PHC2778_n5075 (.Z(FE_PHN2778_n5075), 
	.A(FE_PHN4495_n5075));
   BUF_X32 FE_PHC2777_n5557 (.Z(FE_PHN2777_n5557), 
	.A(FE_PHN4493_n5557));
   BUF_X32 FE_PHC2776_n5141 (.Z(FE_PHN2776_n5141), 
	.A(FE_PHN4518_n5141));
   BUF_X32 FE_PHC2775_n5470 (.Z(FE_PHN2775_n5470), 
	.A(FE_PHN4506_n5470));
   BUF_X32 FE_PHC2774_n5083 (.Z(FE_PHN2774_n5083), 
	.A(FE_PHN4515_n5083));
   BUF_X32 FE_PHC2773_n5170 (.Z(FE_PHN2773_n5170), 
	.A(FE_PHN4511_n5170));
   BUF_X32 FE_PHC2772_n5172 (.Z(FE_PHN2772_n5172), 
	.A(FE_PHN4567_n5172));
   BUF_X32 FE_PHC2771_n5468 (.Z(FE_PHN2771_n5468), 
	.A(FE_PHN4514_n5468));
   BUF_X32 FE_PHC2770_n5178 (.Z(FE_PHN2770_n5178), 
	.A(FE_PHN4554_n5178));
   BUF_X32 FE_PHC2769_n5299 (.Z(FE_PHN2769_n5299), 
	.A(FE_PHN4557_n5299));
   BUF_X32 FE_PHC2768_n5478 (.Z(FE_PHN2768_n5478), 
	.A(FE_PHN4487_n5478));
   BUF_X32 FE_PHC2767_n5450 (.Z(FE_PHN2767_n5450), 
	.A(FE_PHN4563_n5450));
   BUF_X32 FE_PHC2766_n5186 (.Z(FE_PHN2766_n5186), 
	.A(FE_PHN4492_n5186));
   BUF_X32 FE_PHC2765_n5039 (.Z(FE_PHN2765_n5039), 
	.A(FE_PHN4500_n5039));
   BUF_X32 FE_PHC2764_n5173 (.Z(FE_PHN2764_n5173), 
	.A(FE_PHN4477_n5173));
   BUF_X32 FE_PHC2763_n5196 (.Z(FE_PHN2763_n5196), 
	.A(FE_PHN4485_n5196));
   BUF_X32 FE_PHC2762_n5174 (.Z(FE_PHN2762_n5174), 
	.A(FE_PHN4531_n5174));
   BUF_X32 FE_PHC2761_n5472 (.Z(FE_PHN2761_n5472), 
	.A(FE_PHN4494_n5472));
   BUF_X32 FE_PHC2760_n5455 (.Z(FE_PHN2760_n5455), 
	.A(FE_PHN4482_n5455));
   BUF_X32 FE_PHC2759_n5396 (.Z(FE_PHN2759_n5396), 
	.A(FE_PHN4556_n5396));
   BUF_X32 FE_PHC2758_n5296 (.Z(FE_PHN2758_n5296), 
	.A(FE_PHN4452_n5296));
   BUF_X32 FE_PHC2757_n5641 (.Z(FE_PHN2757_n5641), 
	.A(FE_PHN4535_n5641));
   BUF_X32 FE_PHC2756_n4985 (.Z(FE_PHN2756_n4985), 
	.A(FE_PHN4484_n4985));
   BUF_X32 FE_PHC2755_n5461 (.Z(FE_PHN2755_n5461), 
	.A(FE_PHN4496_n5461));
   BUF_X32 FE_PHC2754_n5633 (.Z(FE_PHN2754_n5633), 
	.A(FE_PHN4476_n5633));
   BUF_X32 FE_PHC2753_n5553 (.Z(FE_PHN2753_n5553), 
	.A(FE_PHN4467_n5553));
   BUF_X32 FE_PHC2752_n5187 (.Z(FE_PHN2752_n5187), 
	.A(FE_PHN4538_n5187));
   BUF_X32 FE_PHC2751_n4969 (.Z(FE_PHN2751_n4969), 
	.A(FE_PHN4486_n4969));
   BUF_X32 FE_PHC2750_n5015 (.Z(FE_PHN2750_n5015), 
	.A(FE_PHN4565_n5015));
   BUF_X32 FE_PHC2749_n5598 (.Z(FE_PHN2749_n5598), 
	.A(FE_PHN4451_n5598));
   BUF_X32 FE_PHC2748_n5312 (.Z(FE_PHN2748_n5312), 
	.A(FE_PHN4466_n5312));
   BUF_X32 FE_PHC2747_n5437 (.Z(FE_PHN2747_n5437), 
	.A(FE_PHN4458_n5437));
   BUF_X32 FE_PHC2746_n5428 (.Z(FE_PHN2746_n5428), 
	.A(FE_PHN4539_n5428));
   BUF_X32 FE_PHC2745_n5426 (.Z(FE_PHN2745_n5426), 
	.A(FE_PHN4468_n5426));
   BUF_X32 FE_PHC2744_n5486 (.Z(FE_PHN2744_n5486), 
	.A(FE_PHN4450_n5486));
   BUF_X32 FE_PHC2743_n5597 (.Z(FE_PHN2743_n5597), 
	.A(FE_PHN4475_n5597));
   BUF_X32 FE_PHC2742_n5121 (.Z(FE_PHN2742_n5121), 
	.A(FE_PHN4457_n5121));
   BUF_X32 FE_PHC2741_n5040 (.Z(FE_PHN2741_n5040), 
	.A(FE_PHN4510_n5040));
   BUF_X32 FE_PHC2740_n5420 (.Z(FE_PHN2740_n5420), 
	.A(FE_PHN4545_n5420));
   BUF_X32 FE_PHC2739_n5161 (.Z(FE_PHN2739_n5161), 
	.A(FE_PHN4463_n5161));
   BUF_X32 FE_PHC2738_n5469 (.Z(FE_PHN2738_n5469), 
	.A(FE_PHN4460_n5469));
   BUF_X32 FE_PHC2737_n5135 (.Z(FE_PHN2737_n5135), 
	.A(FE_PHN4532_n5135));
   BUF_X32 FE_PHC2736_n5103 (.Z(FE_PHN2736_n5103), 
	.A(FE_PHN4569_n5103));
   BUF_X32 FE_PHC2735_n5021 (.Z(FE_PHN2735_n5021), 
	.A(FE_PHN4449_n5021));
   BUF_X32 FE_PHC2734_n5464 (.Z(FE_PHN2734_n5464), 
	.A(FE_PHN4436_n5464));
   BUF_X32 FE_PHC2733_n5616 (.Z(FE_PHN2733_n5616), 
	.A(FE_PHN4440_n5616));
   BUF_X32 FE_PHC2732_n5636 (.Z(FE_PHN2732_n5636), 
	.A(FE_PHN4438_n5636));
   BUF_X32 FE_PHC2731_n5138 (.Z(FE_PHN2731_n5138), 
	.A(FE_PHN4499_n5138));
   BUF_X32 FE_PHC2730_n5046 (.Z(FE_PHN2730_n5046), 
	.A(FE_PHN4437_n5046));
   BUF_X32 FE_PHC2729_n5463 (.Z(FE_PHN2729_n5463), 
	.A(FE_PHN4508_n5463));
   BUF_X32 FE_PHC2728_n5115 (.Z(FE_PHN2728_n5115), 
	.A(FE_PHN4517_n5115));
   BUF_X32 FE_PHC2727_n5086 (.Z(FE_PHN2727_n5086), 
	.A(FE_PHN4432_n5086));
   BUF_X32 FE_PHC2726_n5022 (.Z(FE_PHN2726_n5022), 
	.A(FE_PHN4418_n5022));
   BUF_X32 FE_PHC2725_n5392 (.Z(FE_PHN2725_n5392), 
	.A(FE_PHN4422_n5392));
   BUF_X32 FE_PHC2724_n5477 (.Z(FE_PHN2724_n5477), 
	.A(FE_PHN4421_n5477));
   BUF_X32 FE_PHC2723_n5485 (.Z(FE_PHN2723_n5485), 
	.A(FE_PHN4430_n5485));
   BUF_X32 FE_PHC2722_n5012 (.Z(FE_PHN2722_n5012), 
	.A(FE_PHN4564_n5012));
   BUF_X32 FE_PHC2721_n5433 (.Z(FE_PHN2721_n5433), 
	.A(FE_PHN4525_n5433));
   BUF_X32 FE_PHC2720_n5020 (.Z(FE_PHN2720_n5020), 
	.A(FE_PHN4427_n5020));
   BUF_X32 FE_PHC2719_n5181 (.Z(FE_PHN2719_n5181), 
	.A(FE_PHN4504_n5181));
   BUF_X32 FE_PHC2718_n5300 (.Z(FE_PHN2718_n5300), 
	.A(FE_PHN4529_n5300));
   BUF_X32 FE_PHC2717_n5438 (.Z(FE_PHN2717_n5438), 
	.A(FE_PHN4403_n5438));
   BUF_X32 FE_PHC2716_n5366 (.Z(FE_PHN2716_n5366), 
	.A(FE_PHN4426_n5366));
   BUF_X32 FE_PHC2715_n5397 (.Z(FE_PHN2715_n5397), 
	.A(FE_PHN4400_n5397));
   BUF_X32 FE_PHC2714_n5442 (.Z(FE_PHN2714_n5442), 
	.A(FE_PHN4412_n5442));
   BUF_X32 FE_PHC2713_n5171 (.Z(FE_PHN2713_n5171), 
	.A(FE_PHN4404_n5171));
   BUF_X32 FE_PHC2712_n5287 (.Z(FE_PHN2712_n5287), 
	.A(FE_PHN4401_n5287));
   BUF_X32 FE_PHC2711_n5453 (.Z(FE_PHN2711_n5453), 
	.A(FE_PHN4490_n5453));
   BUF_X32 FE_PHC2710_n5427 (.Z(FE_PHN2710_n5427), 
	.A(FE_PHN4474_n5427));
   BUF_X32 FE_PHC2709_n5564 (.Z(FE_PHN2709_n5564), 
	.A(FE_PHN4462_n5564));
   BUF_X32 FE_PHC2708_n5452 (.Z(FE_PHN2708_n5452), 
	.A(FE_PHN4396_n5452));
   BUF_X32 FE_PHC2707_n5459 (.Z(FE_PHN2707_n5459), 
	.A(FE_PHN4481_n5459));
   BUF_X32 FE_PHC2706_n5575 (.Z(FE_PHN2706_n5575), 
	.A(FE_PHN4392_n5575));
   BUF_X32 FE_PHC2705_n5432 (.Z(FE_PHN2705_n5432), 
	.A(FE_PHN4406_n5432));
   BUF_X32 FE_PHC2703_n5197 (.Z(FE_PHN2703_n5197), 
	.A(FE_PHN4456_n5197));
   BUF_X32 FE_PHC2702_n5449 (.Z(FE_PHN2702_n5449), 
	.A(FE_PHN4548_n5449));
   BUF_X32 FE_PHC2701_n5430 (.Z(FE_PHN2701_n5430), 
	.A(FE_PHN4413_n5430));
   BUF_X32 FE_PHC2700_n5069 (.Z(FE_PHN2700_n5069), 
	.A(FE_PHN4387_n5069));
   BUF_X32 FE_PHC2699_n5462 (.Z(FE_PHN2699_n5462), 
	.A(FE_PHN4393_n5462));
   BUF_X32 FE_PHC2698_n5439 (.Z(FE_PHN2698_n5439), 
	.A(FE_PHN4386_n5439));
   BUF_X32 FE_PHC2697_n5184 (.Z(FE_PHN2697_n5184), 
	.A(FE_PHN4376_n5184));
   BUF_X32 FE_PHC2696_n5424 (.Z(FE_PHN2696_n5424), 
	.A(FE_PHN4382_n5424));
   BUF_X32 FE_PHC2695_n5401 (.Z(FE_PHN2695_n5401), 
	.A(FE_PHN4459_n5401));
   BUF_X32 FE_PHC2694_n5466 (.Z(FE_PHN2694_n5466), 
	.A(FE_PHN4375_n5466));
   BUF_X32 FE_PHC2693_n5190 (.Z(FE_PHN2693_n5190), 
	.A(FE_PHN4471_n5190));
   BUF_X32 FE_PHC2692_n5398 (.Z(FE_PHN2692_n5398), 
	.A(FE_PHN4417_n5398));
   BUF_X32 FE_PHC2691_n5550 (.Z(FE_PHN2691_n5550), 
	.A(FE_PHN4380_n5550));
   BUF_X32 FE_PHC2690_n5051 (.Z(FE_PHN2690_n5051), 
	.A(FE_PHN4351_n5051));
   BUF_X32 FE_PHC2689_n5043 (.Z(FE_PHN2689_n5043), 
	.A(FE_PHN4362_n5043));
   BUF_X32 FE_PHC2688_n5421 (.Z(FE_PHN2688_n5421), 
	.A(FE_PHN4377_n5421));
   BUF_X32 FE_PHC2687_n5175 (.Z(FE_PHN2687_n5175), 
	.A(FE_PHN4371_n5175));
   BUF_X32 FE_PHC2686_n5576 (.Z(FE_PHN2686_n5576), 
	.A(FE_PHN4448_n5576));
   BUF_X32 FE_PHC2685_n5030 (.Z(FE_PHN2685_n5030), 
	.A(FE_PHN4373_n5030));
   BUF_X32 FE_PHC2684_n5010 (.Z(FE_PHN2684_n5010), 
	.A(FE_PHN4372_n5010));
   BUF_X32 FE_PHC2683_n5191 (.Z(FE_PHN2683_n5191), 
	.A(FE_PHN4356_n5191));
   BUF_X32 FE_PHC2682_n5447 (.Z(FE_PHN2682_n5447), 
	.A(FE_PHN4444_n5447));
   BUF_X32 FE_PHC2681_n5108 (.Z(FE_PHN2681_n5108), 
	.A(FE_PHN4363_n5108));
   BUF_X32 FE_PHC2680_n5041 (.Z(FE_PHN2680_n5041), 
	.A(FE_PHN4369_n5041));
   BUF_X32 FE_PHC2679_n5123 (.Z(FE_PHN2679_n5123), 
	.A(FE_PHN4368_n5123));
   BUF_X32 FE_PHC2678_n5606 (.Z(FE_PHN2678_n5606), 
	.A(FE_PHN4399_n5606));
   BUF_X32 FE_PHC2676_n4987 (.Z(FE_PHN2676_n4987), 
	.A(FE_PHN4361_n4987));
   BUF_X32 FE_PHC2675_n5539 (.Z(FE_PHN2675_n5539), 
	.A(FE_PHN4420_n5539));
   BUF_X32 FE_PHC2674_n5476 (.Z(FE_PHN2674_n5476), 
	.A(FE_PHN4405_n5476));
   BUF_X32 FE_PHC2673_n5091 (.Z(FE_PHN2673_n5091), 
	.A(FE_PHN4350_n5091));
   BUF_X32 FE_PHC2672_n5538 (.Z(FE_PHN2672_n5538), 
	.A(FE_PHN5107_n5538));
   BUF_X32 FE_PHC2671_n5473 (.Z(FE_PHN2671_n5473), 
	.A(FE_PHN4352_n5473));
   BUF_X32 FE_PHC2670_n5192 (.Z(FE_PHN2670_n5192), 
	.A(FE_PHN4357_n5192));
   BUF_X32 FE_PHC2669_n5434 (.Z(FE_PHN2669_n5434), 
	.A(FE_PHN4411_n5434));
   BUF_X32 FE_PHC2668_n5444 (.Z(FE_PHN2668_n5444), 
	.A(FE_PHN4419_n5444));
   BUF_X32 FE_PHC2667_n5183 (.Z(FE_PHN2667_n5183), 
	.A(FE_PHN4327_n5183));
   BUF_X32 FE_PHC2666_n5106 (.Z(FE_PHN2666_n5106), 
	.A(FE_PHN4340_n5106));
   BUF_X32 FE_PHC2665_n5410 (.Z(FE_PHN2665_n5410), 
	.A(FE_PHN4348_n5410));
   BUF_X32 FE_PHC2664_n5093 (.Z(FE_PHN2664_n5093), 
	.A(FE_PHN4446_n5093));
   BUF_X32 FE_PHC2663_n5195 (.Z(FE_PHN2663_n5195), 
	.A(FE_PHN4311_n5195));
   BUF_X32 FE_PHC2662_n5132 (.Z(FE_PHN2662_n5132), 
	.A(FE_PHN4338_n5132));
   BUF_X32 FE_PHC2661_n5304 (.Z(FE_PHN2661_n5304), 
	.A(FE_PHN4336_n5304));
   BUF_X32 FE_PHC2660_n5567 (.Z(FE_PHN2660_n5567), 
	.A(FE_PHN4447_n5567));
   BUF_X32 FE_PHC2659_n5435 (.Z(FE_PHN2659_n5435), 
	.A(FE_PHN4330_n5435));
   BUF_X32 FE_PHC2658_n5448 (.Z(FE_PHN2658_n5448), 
	.A(FE_PHN4378_n5448));
   BUF_X32 FE_PHC2657_n5399 (.Z(FE_PHN2657_n5399), 
	.A(FE_PHN4331_n5399));
   BUF_X32 FE_PHC2655_n5393 (.Z(FE_PHN2655_n5393), 
	.A(FE_PHN4334_n5393));
   BUF_X32 FE_PHC2654_n5411 (.Z(FE_PHN2654_n5411), 
	.A(FE_PHN4367_n5411));
   BUF_X32 FE_PHC2653_n5451 (.Z(FE_PHN2653_n5451), 
	.A(FE_PHN4320_n5451));
   BUF_X32 FE_PHC2652_n5298 (.Z(FE_PHN2652_n5298), 
	.A(FE_PHN4374_n5298));
   BUF_X32 FE_PHC2651_n5412 (.Z(FE_PHN2651_n5412), 
	.A(FE_PHN4379_n5412));
   BUF_X32 FE_PHC2650_n5289 (.Z(FE_PHN2650_n5289), 
	.A(FE_PHN4317_n5289));
   BUF_X32 FE_PHC2649_n5182 (.Z(FE_PHN2649_n5182), 
	.A(FE_PHN4385_n5182));
   BUF_X32 FE_PHC2648_n4986 (.Z(FE_PHN2648_n4986), 
	.A(FE_PHN4325_n4986));
   BUF_X32 FE_PHC2647_n5189 (.Z(FE_PHN2647_n5189), 
	.A(FE_PHN4319_n5189));
   BUF_X32 FE_PHC2646_n5440 (.Z(FE_PHN2646_n5440), 
	.A(FE_PHN4302_n5440));
   BUF_X32 FE_PHC2645_n5301 (.Z(FE_PHN2645_n5301), 
	.A(FE_PHN4279_n5301));
   BUF_X32 FE_PHC2644_n5558 (.Z(FE_PHN2644_n5558), 
	.A(FE_PHN4425_n5558));
   BUF_X32 FE_PHC2643_n5180 (.Z(FE_PHN2643_n5180), 
	.A(FE_PHN4332_n5180));
   BUF_X32 FE_PHC2642_n5414 (.Z(FE_PHN2642_n5414), 
	.A(FE_PHN4366_n5414));
   BUF_X32 FE_PHC2641_n5441 (.Z(FE_PHN2641_n5441), 
	.A(FE_PHN4355_n5441));
   BUF_X32 FE_PHC2640_n5418 (.Z(FE_PHN2640_n5418), 
	.A(FE_PHN4282_n5418));
   BUF_X32 FE_PHC2639_n5643 (.Z(FE_PHN2639_n5643), 
	.A(FE_PHN5002_n5643));
   BUF_X32 FE_PHC2637_n5395 (.Z(FE_PHN2637_n5395), 
	.A(FE_PHN4333_n5395));
   BUF_X32 FE_PHC2636_n5363 (.Z(FE_PHN2636_n5363), 
	.A(FE_PHN4267_n5363));
   BUF_X32 FE_PHC2635_n5207 (.Z(FE_PHN2635_n5207), 
	.A(FE_PHN4291_n5207));
   BUF_X32 FE_PHC2634_n5028 (.Z(FE_PHN2634_n5028), 
	.A(FE_PHN4263_n5028));
   BUF_X32 FE_PHC2633_n5176 (.Z(FE_PHN2633_n5176), 
	.A(FE_PHN4274_n5176));
   BUF_X32 FE_PHC2632_n5419 (.Z(FE_PHN2632_n5419), 
	.A(FE_PHN4343_n5419));
   BUF_X32 FE_PHC2631_n5203 (.Z(FE_PHN2631_n5203), 
	.A(FE_PHN4248_n5203));
   BUF_X32 FE_PHC2630_n5629 (.Z(FE_PHN2630_n5629), 
	.A(FE_PHN4314_n5629));
   BUF_X32 FE_PHC2629_n5409 (.Z(FE_PHN2629_n5409), 
	.A(FE_PHN4301_n5409));
   BUF_X32 FE_PHC2628_n5348 (.Z(FE_PHN2628_n5348), 
	.A(FE_PHN4182_n5348));
   BUF_X32 FE_PHC2627_n5013 (.Z(FE_PHN2627_n5013), 
	.A(FE_PHN4262_n5013));
   BUF_X32 FE_PHC2626_n5360 (.Z(FE_PHN2626_n5360), 
	.A(FE_PHN5136_n5360));
   BUF_X32 FE_PHC2625_n5266 (.Z(FE_PHN2625_n5266), 
	.A(FE_PHN4193_n5266));
   BUF_X32 FE_PHC2624_n5415 (.Z(FE_PHN2624_n5415), 
	.A(FE_PHN4287_n5415));
   BUF_X32 FE_PHC2623_n5159 (.Z(FE_PHN2623_n5159), 
	.A(FE_PHN5146_n5159));
   BUF_X32 FE_PHC2622_n5483 (.Z(FE_PHN2622_n5483), 
	.A(FE_PHN5155_n5483));
   BUF_X32 FE_PHC2621_n5521 (.Z(FE_PHN2621_n5521), 
	.A(FE_PHN4318_n5521));
   BUF_X32 FE_PHC2620_n5367 (.Z(FE_PHN2620_n5367), 
	.A(FE_PHN5059_n5367));
   BUF_X32 FE_PHC2619_n5273 (.Z(FE_PHN2619_n5273), 
	.A(FE_PHN4931_n5273));
   BUF_X32 FE_PHC2618_n5596 (.Z(FE_PHN2618_n5596), 
	.A(FE_PHN4313_n5596));
   BUF_X32 FE_PHC2617_n5481 (.Z(FE_PHN2617_n5481), 
	.A(FE_PHN4261_n5481));
   BUF_X32 FE_PHC2616_n5205 (.Z(FE_PHN2616_n5205), 
	.A(FE_PHN4329_n5205));
   BUF_X32 FE_PHC2615_n5045 (.Z(FE_PHN2615_n5045), 
	.A(FE_PHN4260_n5045));
   BUF_X32 FE_PHC2614_n4979 (.Z(FE_PHN2614_n4979), 
	.A(FE_PHN5158_n4979));
   BUF_X32 FE_PHC2613_n5270 (.Z(FE_PHN2613_n5270), 
	.A(FE_PHN4247_n5270));
   BUF_X32 FE_PHC2612_n5199 (.Z(FE_PHN2612_n5199), 
	.A(FE_PHN4312_n5199));
   BUF_X32 FE_PHC2611_n5436 (.Z(FE_PHN2611_n5436), 
	.A(FE_PHN4295_n5436));
   BUF_X32 FE_PHC2610_n5308 (.Z(FE_PHN2610_n5308), 
	.A(FE_PHN5124_n5308));
   BUF_X32 FE_PHC2609_n5112 (.Z(FE_PHN2609_n5112), 
	.A(FE_PHN4200_n5112));
   BUF_X32 FE_PHC2608_n5624 (.Z(FE_PHN2608_n5624), 
	.A(FE_PHN4280_n5624));
   BUF_X32 FE_PHC2607_n5076 (.Z(FE_PHN2607_n5076), 
	.A(FE_PHN4237_n5076));
   BUF_X32 FE_PHC2606_n5364 (.Z(FE_PHN2606_n5364), 
	.A(FE_PHN5106_n5364));
   BUF_X32 FE_PHC2605_n5384 (.Z(FE_PHN2605_n5384), 
	.A(FE_PHN5027_n5384));
   BUF_X32 FE_PHC2604_n5309 (.Z(FE_PHN2604_n5309), 
	.A(FE_PHN4283_n5309));
   BUF_X32 FE_PHC2603_n5343 (.Z(FE_PHN2603_n5343), 
	.A(FE_PHN4833_n5343));
   BUF_X32 FE_PHC2602_n5386 (.Z(FE_PHN2602_n5386), 
	.A(FE_PHN4335_n5386));
   BUF_X32 FE_PHC2601_n5413 (.Z(FE_PHN2601_n5413), 
	.A(FE_PHN5134_n5413));
   BUF_X32 FE_PHC2600_n5362 (.Z(FE_PHN2600_n5362), 
	.A(FE_PHN5160_n5362));
   BUF_X32 FE_PHC2599_n5361 (.Z(FE_PHN2599_n5361), 
	.A(FE_PHN5156_n5361));
   BUF_X32 FE_PHC2598_n5224 (.Z(FE_PHN2598_n5224), 
	.A(FE_PHN4234_n5224));
   BUF_X32 FE_PHC2597_n5422 (.Z(FE_PHN2597_n5422), 
	.A(FE_PHN4305_n5422));
   BUF_X32 FE_PHC2596_n5261 (.Z(FE_PHN2596_n5261), 
	.A(FE_PHN4972_n5261));
   BUF_X32 FE_PHC2595_n5357 (.Z(FE_PHN2595_n5357), 
	.A(FE_PHN4947_n5357));
   BUF_X32 FE_PHC2594_n5443 (.Z(FE_PHN2594_n5443), 
	.A(FE_PHN5125_n5443));
   BUF_X32 FE_PHC2593_n5638 (.Z(FE_PHN2593_n5638), 
	.A(FE_PHN4215_n5638));
   BUF_X32 FE_PHC2592_n5219 (.Z(FE_PHN2592_n5219), 
	.A(FE_PHN4109_n5219));
   BUF_X32 FE_PHC2591_n5394 (.Z(FE_PHN2591_n5394), 
	.A(FE_PHN4967_n5394));
   BUF_X32 FE_PHC2590_n5554 (.Z(FE_PHN2590_n5554), 
	.A(FE_PHN4181_n5554));
   BUF_X32 FE_PHC2589_n5081 (.Z(FE_PHN2589_n5081), 
	.A(FE_PHN5167_n5081));
   BUF_X32 FE_PHC2588_n5225 (.Z(FE_PHN2588_n5225), 
	.A(FE_PHN4273_n5225));
   BUF_X32 FE_PHC2587_n5374 (.Z(FE_PHN2587_n5374), 
	.A(FE_PHN4904_n5374));
   BUF_X32 FE_PHC2586_n5049 (.Z(FE_PHN2586_n5049), 
	.A(FE_PHN4259_n5049));
   BUF_X32 FE_PHC2585_n4995 (.Z(FE_PHN2585_n4995), 
	.A(FE_PHN5028_n4995));
   BUF_X32 FE_PHC2584_n5202 (.Z(FE_PHN2584_n5202), 
	.A(FE_PHN5086_n5202));
   BUF_X32 FE_PHC2583_n5070 (.Z(FE_PHN2583_n5070), 
	.A(FE_PHN4178_n5070));
   BUF_X32 FE_PHC2582_n5403 (.Z(FE_PHN2582_n5403), 
	.A(FE_PHN4950_n5403));
   BUF_X32 FE_PHC2581_n5107 (.Z(FE_PHN2581_n5107), 
	.A(FE_PHN4161_n5107));
   BUF_X32 FE_PHC2580_n5271 (.Z(FE_PHN2580_n5271), 
	.A(FE_PHN5053_n5271));
   BUF_X32 FE_PHC2579_n5128 (.Z(FE_PHN2579_n5128), 
	.A(FE_PHN5151_n5128));
   BUF_X32 FE_PHC2578_n5125 (.Z(FE_PHN2578_n5125), 
	.A(FE_PHN4790_n5125));
   BUF_X32 FE_PHC2577_n5079 (.Z(FE_PHN2577_n5079), 
	.A(FE_PHN4217_n5079));
   BUF_X32 FE_PHC2576_n5201 (.Z(FE_PHN2576_n5201), 
	.A(FE_PHN5090_n5201));
   BUF_X32 FE_PHC2574_n5019 (.Z(FE_PHN2574_n5019), 
	.A(FE_PHN5008_n5019));
   BUF_X32 FE_PHC2573_n5405 (.Z(FE_PHN2573_n5405), 
	.A(FE_PHN4145_n5405));
   BUF_X32 FE_PHC2572_n5365 (.Z(FE_PHN2572_n5365), 
	.A(FE_PHN4970_n5365));
   BUF_X32 FE_PHC2571_n5355 (.Z(FE_PHN2571_n5355), 
	.A(FE_PHN5088_n5355));
   BUF_X32 FE_PHC2570_n5479 (.Z(FE_PHN2570_n5479), 
	.A(FE_PHN4902_n5479));
   BUF_X32 FE_PHC2569_n5136 (.Z(FE_PHN2569_n5136), 
	.A(FE_PHN5060_n5136));
   BUF_X32 FE_PHC2568_n5200 (.Z(FE_PHN2568_n5200), 
	.A(FE_PHN5045_n5200));
   BUF_X32 FE_PHC2566_n5336 (.Z(FE_PHN2566_n5336), 
	.A(FE_PHN4994_n5336));
   BUF_X32 FE_PHC2564_n5319 (.Z(FE_PHN2564_n5319), 
	.A(FE_PHN5139_n5319));
   BUF_X32 FE_PHC2563_n5372 (.Z(FE_PHN2563_n5372), 
	.A(FE_PHN4946_n5372));
   BUF_X32 FE_PHC2562_n5278 (.Z(FE_PHN2562_n5278), 
	.A(FE_PHN4861_n5278));
   BUF_X32 FE_PHC2561_n5139 (.Z(FE_PHN2561_n5139), 
	.A(FE_PHN4167_n5139));
   BUF_X32 FE_PHC2560_n5560 (.Z(FE_PHN2560_n5560), 
	.A(FE_PHN4149_n5560));
   BUF_X32 FE_PHC2559_n5368 (.Z(FE_PHN2559_n5368), 
	.A(FE_PHN4795_n5368));
   BUF_X32 FE_PHC2557_n5369 (.Z(FE_PHN2557_n5369), 
	.A(FE_PHN5130_n5369));
   BUF_X32 FE_PHC2556_n5640 (.Z(FE_PHN2556_n5640), 
	.A(FE_PHN5006_n5640));
   BUF_X32 FE_PHC2555_n5335 (.Z(FE_PHN2555_n5335), 
	.A(FE_PHN4912_n5335));
   BUF_X32 FE_PHC2554_n5316 (.Z(FE_PHN2554_n5316), 
	.A(FE_PHN4346_n5316));
   BUF_X32 FE_PHC2553_n5218 (.Z(FE_PHN2553_n5218), 
	.A(FE_PHN4988_n5218));
   BUF_X32 FE_PHC2552_n5562 (.Z(FE_PHN2552_n5562), 
	.A(FE_PHN4101_n5562));
   BUF_X32 FE_PHC2551_n5268 (.Z(FE_PHN2551_n5268), 
	.A(FE_PHN4230_n5268));
   BUF_X32 FE_PHC2550_n5131 (.Z(FE_PHN2550_n5131), 
	.A(FE_PHN4838_n5131));
   BUF_X32 FE_PHC2549_n5334 (.Z(FE_PHN2549_n5334), 
	.A(FE_PHN4870_n5334));
   BUF_X32 FE_PHC2548_n5213 (.Z(FE_PHN2548_n5213), 
	.A(FE_PHN4154_n5213));
   BUF_X32 FE_PHC2547_n5383 (.Z(FE_PHN2547_n5383), 
	.A(FE_PHN5052_n5383));
   BUF_X32 FE_PHC2546_n5018 (.Z(FE_PHN2546_n5018), 
	.A(FE_PHN5127_n5018));
   BUF_X32 FE_PHC2545_n5317 (.Z(FE_PHN2545_n5317), 
	.A(FE_PHN4227_n5317));
   BUF_X32 FE_PHC2544_n5621 (.Z(FE_PHN2544_n5621), 
	.A(FE_PHN4214_n5621));
   BUF_X32 FE_PHC2543_n5217 (.Z(FE_PHN2543_n5217), 
	.A(FE_PHN4140_n5217));
   BUF_X32 FE_PHC2542_n5491 (.Z(FE_PHN2542_n5491), 
	.A(FE_PHN5129_n5491));
   BUF_X32 FE_PHC2541_n5356 (.Z(FE_PHN2541_n5356), 
	.A(FE_PHN4963_n5356));
   BUF_X32 FE_PHC2540_n5063 (.Z(FE_PHN2540_n5063), 
	.A(FE_PHN4853_n5063));
   BUF_X32 FE_PHC2539_n5347 (.Z(FE_PHN2539_n5347), 
	.A(FE_PHN5149_n5347));
   BUF_X32 FE_PHC2538_n5109 (.Z(FE_PHN2538_n5109), 
	.A(FE_PHN4995_n5109));
   BUF_X32 FE_PHC2537_n5211 (.Z(FE_PHN2537_n5211), 
	.A(FE_PHN4004_n5211));
   BUF_X32 FE_PHC2536_n5209 (.Z(FE_PHN2536_n5209), 
	.A(FE_PHN5055_n5209));
   BUF_X32 FE_PHC2535_n5339 (.Z(FE_PHN2535_n5339), 
	.A(FE_PHN5044_n5339));
   BUF_X32 FE_PHC2534_n5630 (.Z(FE_PHN2534_n5630), 
	.A(FE_PHN4874_n5630));
   BUF_X32 FE_PHC2533_n5349 (.Z(FE_PHN2533_n5349), 
	.A(FE_PHN5169_n5349));
   BUF_X32 FE_PHC2532_n5376 (.Z(FE_PHN2532_n5376), 
	.A(FE_PHN5001_n5376));
   BUF_X32 FE_PHC2531_n5566 (.Z(FE_PHN2531_n5566), 
	.A(FE_PHN4873_n5566));
   BUF_X32 FE_PHC2530_n5133 (.Z(FE_PHN2530_n5133), 
	.A(FE_PHN5108_n5133));
   BUF_X32 FE_PHC2529_n5634 (.Z(FE_PHN2529_n5634), 
	.A(FE_PHN4974_n5634));
   BUF_X32 FE_PHC2528_n5283 (.Z(FE_PHN2528_n5283), 
	.A(FE_PHN4980_n5283));
   BUF_X32 FE_PHC2527_n5279 (.Z(FE_PHN2527_n5279), 
	.A(FE_PHN5114_n5279));
   BUF_X32 FE_PHC2526_n5044 (.Z(FE_PHN2526_n5044), 
	.A(FE_PHN4076_n5044));
   BUF_X32 FE_PHC2525_n5381 (.Z(FE_PHN2525_n5381), 
	.A(FE_PHN5023_n5381));
   BUF_X32 FE_PHC2524_n5292 (.Z(FE_PHN2524_n5292), 
	.A(FE_PHN4067_n5292));
   BUF_X32 FE_PHC2523_n5563 (.Z(FE_PHN2523_n5563), 
	.A(FE_PHN4859_n5563));
   BUF_X32 FE_PHC2522_n5378 (.Z(FE_PHN2522_n5378), 
	.A(FE_PHN5150_n5378));
   BUF_X32 FE_PHC2521_n5263 (.Z(FE_PHN2521_n5263), 
	.A(FE_PHN4802_n5263));
   BUF_X32 FE_PHC2520_n5212 (.Z(FE_PHN2520_n5212), 
	.A(FE_PHN3912_n5212));
   BUF_X32 FE_PHC2519_n5221 (.Z(FE_PHN2519_n5221), 
	.A(FE_PHN5017_n5221));
   BUF_X32 FE_PHC2518_n5543 (.Z(FE_PHN2518_n5543), 
	.A(FE_PHN4801_n5543));
   BUF_X32 FE_PHC2517_n5220 (.Z(FE_PHN2517_n5220), 
	.A(FE_PHN5093_n5220));
   BUF_X32 FE_PHC2516_n5542 (.Z(FE_PHN2516_n5542), 
	.A(FE_PHN4233_n5542));
   BUF_X32 FE_PHC2515_n5617 (.Z(FE_PHN2515_n5617), 
	.A(FE_PHN5120_n5617));
   BUF_X32 FE_PHC2514_n5610 (.Z(FE_PHN2514_n5610), 
	.A(FE_PHN5137_n5610));
   BUF_X32 FE_PHC2513_n5280 (.Z(FE_PHN2513_n5280), 
	.A(FE_PHN5126_n5280));
   BUF_X32 FE_PHC2512_n5391 (.Z(FE_PHN2512_n5391), 
	.A(FE_PHN5135_n5391));
   BUF_X32 FE_PHC2511_n5104 (.Z(FE_PHN2511_n5104), 
	.A(FE_PHN5034_n5104));
   BUF_X32 FE_PHC2510_n5599 (.Z(FE_PHN2510_n5599), 
	.A(FE_PHN4976_n5599));
   BUF_X32 FE_PHC2509_n5124 (.Z(FE_PHN2509_n5124), 
	.A(FE_PHN4123_n5124));
   BUF_X32 FE_PHC2508_n5264 (.Z(FE_PHN2508_n5264), 
	.A(FE_PHN4809_n5264));
   BUF_X32 FE_PHC2507_n5084 (.Z(FE_PHN2507_n5084), 
	.A(FE_PHN5029_n5084));
   BUF_X32 FE_PHC2506_n5480 (.Z(FE_PHN2506_n5480), 
	.A(FE_PHN4876_n5480));
   BUF_X32 FE_PHC2505_n5385 (.Z(FE_PHN2505_n5385), 
	.A(FE_PHN3975_n5385));
   BUF_X32 FE_PHC2504_n5337 (.Z(FE_PHN2504_n5337), 
	.A(FE_PHN5085_n5337));
   BUF_X32 FE_PHC2503_n5497 (.Z(FE_PHN2503_n5497), 
	.A(FE_PHN4910_n5497));
   BUF_X32 FE_PHC2502_n5037 (.Z(FE_PHN2502_n5037), 
	.A(FE_PHN4866_n5037));
   BUF_X32 FE_PHC2501_n4984 (.Z(FE_PHN2501_n4984), 
	.A(FE_PHN4000_n4984));
   BUF_X32 FE_PHC2500_n5216 (.Z(FE_PHN2500_n5216), 
	.A(FE_PHN4886_n5216));
   BUF_X32 FE_PHC2499_n5142 (.Z(FE_PHN2499_n5142), 
	.A(FE_PHN5094_n5142));
   BUF_X32 FE_PHC2498_n5350 (.Z(FE_PHN2498_n5350), 
	.A(FE_PHN4959_n5350));
   BUF_X32 FE_PHC2497_n5602 (.Z(FE_PHN2497_n5602), 
	.A(FE_PHN5035_n5602));
   BUF_X32 FE_PHC2496_n5052 (.Z(FE_PHN2496_n5052), 
	.A(FE_PHN5122_n5052));
   BUF_X32 FE_PHC2495_n5042 (.Z(FE_PHN2495_n5042), 
	.A(FE_PHN5061_n5042));
   BUF_X32 FE_PHC2494_n5489 (.Z(FE_PHN2494_n5489), 
	.A(FE_PHN5015_n5489));
   BUF_X32 FE_PHC2493_n5198 (.Z(FE_PHN2493_n5198), 
	.A(FE_PHN4969_n5198));
   BUF_X32 FE_PHC2492_n5611 (.Z(FE_PHN2492_n5611), 
	.A(FE_PHN5099_n5611));
   BUF_X32 FE_PHC2491_n5066 (.Z(FE_PHN2491_n5066), 
	.A(FE_PHN4953_n5066));
   BUF_X32 FE_PHC2490_n5294 (.Z(FE_PHN2490_n5294), 
	.A(FE_PHN5014_n5294));
   BUF_X32 FE_PHC2489_n5087 (.Z(FE_PHN2489_n5087), 
	.A(FE_PHN4827_n5087));
   BUF_X32 FE_PHC2488_n4998 (.Z(FE_PHN2488_n4998), 
	.A(FE_PHN4888_n4998));
   BUF_X32 FE_PHC2487_n5607 (.Z(FE_PHN2487_n5607), 
	.A(FE_PHN4821_n5607));
   BUF_X32 FE_PHC2486_n5276 (.Z(FE_PHN2486_n5276), 
	.A(FE_PHN4854_n5276));
   BUF_X32 FE_PHC2485_n5379 (.Z(FE_PHN2485_n5379), 
	.A(FE_PHN4940_n5379));
   BUF_X32 FE_PHC2484_n5574 (.Z(FE_PHN2484_n5574), 
	.A(FE_PHN4828_n5574));
   BUF_X32 FE_PHC2483_n5226 (.Z(FE_PHN2483_n5226), 
	.A(FE_PHN4933_n5226));
   BUF_X32 FE_PHC2482_n5352 (.Z(FE_PHN2482_n5352), 
	.A(FE_PHN5168_n5352));
   BUF_X32 FE_PHC2481_n5277 (.Z(FE_PHN2481_n5277), 
	.A(FE_PHN4909_n5277));
   BUF_X32 FE_PHC2480_n5494 (.Z(FE_PHN2480_n5494), 
	.A(FE_PHN4919_n5494));
   BUF_X32 FE_PHC2479_n5116 (.Z(FE_PHN2479_n5116), 
	.A(FE_PHN3927_n5116));
   BUF_X32 FE_PHC2478_n5631 (.Z(FE_PHN2478_n5631), 
	.A(FE_PHN4823_n5631));
   BUF_X32 FE_PHC2477_n5380 (.Z(FE_PHN2477_n5380), 
	.A(FE_PHN4971_n5380));
   BUF_X32 FE_PHC2476_n5548 (.Z(FE_PHN2476_n5548), 
	.A(FE_PHN4782_n5548));
   BUF_X32 FE_PHC2475_n5215 (.Z(FE_PHN2475_n5215), 
	.A(FE_PHN4794_n5215));
   BUF_X32 FE_PHC2474_n5214 (.Z(FE_PHN2474_n5214), 
	.A(FE_PHN4955_n5214));
   BUF_X32 FE_PHC2473_n5092 (.Z(FE_PHN2473_n5092), 
	.A(FE_PHN4990_n5092));
   BUF_X32 FE_PHC2472_n5122 (.Z(FE_PHN2472_n5122), 
	.A(FE_PHN4796_n5122));
   BUF_X32 FE_PHC2471_n5089 (.Z(FE_PHN2471_n5089), 
	.A(FE_PHN5121_n5089));
   BUF_X32 FE_PHC2470_n5382 (.Z(FE_PHN2470_n5382), 
	.A(FE_PHN4847_n5382));
   BUF_X32 FE_PHC2469_n5351 (.Z(FE_PHN2469_n5351), 
	.A(FE_PHN3923_n5351));
   BUF_X32 FE_PHC2468_n5260 (.Z(FE_PHN2468_n5260), 
	.A(FE_PHN5074_n5260));
   BUF_X32 FE_PHC2467_n5492 (.Z(FE_PHN2467_n5492), 
	.A(FE_PHN5019_n5492));
   BUF_X32 FE_PHC2466_n5493 (.Z(FE_PHN2466_n5493), 
	.A(FE_PHN5018_n5493));
   BUF_X32 FE_PHC2465_n5559 (.Z(FE_PHN2465_n5559), 
	.A(FE_PHN4885_n5559));
   BUF_X32 FE_PHC2464_n5318 (.Z(FE_PHN2464_n5318), 
	.A(FE_PHN4257_n5318));
   BUF_X32 FE_PHC2463_n5354 (.Z(FE_PHN2463_n5354), 
	.A(FE_PHN4883_n5354));
   BUF_X32 FE_PHC2462_n5627 (.Z(FE_PHN2462_n5627), 
	.A(FE_PHN4784_n5627));
   BUF_X32 FE_PHC2461_n5490 (.Z(FE_PHN2461_n5490), 
	.A(FE_PHN4997_n5490));
   BUF_X32 FE_PHC2460_n5286 (.Z(FE_PHN2460_n5286), 
	.A(FE_PHN4924_n5286));
   BUF_X32 FE_PHC2459_n5608 (.Z(FE_PHN2459_n5608), 
	.A(FE_PHN4868_n5608));
   BUF_X32 FE_PHC2458_n5353 (.Z(FE_PHN2458_n5353), 
	.A(FE_PHN4977_n5353));
   BUF_X32 FE_PHC2457_n5635 (.Z(FE_PHN2457_n5635), 
	.A(FE_PHN4050_n5635));
   BUF_X32 FE_PHC2456_n5496 (.Z(FE_PHN2456_n5496), 
	.A(FE_PHN4989_n5496));
   BUF_X32 FE_PHC2454_n5345 (.Z(FE_PHN2454_n5345), 
	.A(FE_PHN4808_n5345));
   BUF_X32 FE_PHC2453_n5541 (.Z(FE_PHN2453_n5541), 
	.A(FE_PHN4906_n5541));
   BUF_X32 FE_PHC2452_n5569 (.Z(FE_PHN2452_n5569), 
	.A(FE_PHN4839_n5569));
   BUF_X32 FE_PHC2451_n4963 (.Z(FE_PHN2451_n4963), 
	.A(FE_PHN5046_n4963));
   BUF_X32 FE_PHC2450_n5341 (.Z(FE_PHN2450_n5341), 
	.A(FE_PHN4887_n5341));
   BUF_X32 FE_PHC2449_n5370 (.Z(FE_PHN2449_n5370), 
	.A(FE_PHN3910_n5370));
   BUF_X32 FE_PHC2448_n5614 (.Z(FE_PHN2448_n5614), 
	.A(FE_PHN4778_n5614));
   BUF_X32 FE_PHC2447_n5275 (.Z(FE_PHN2447_n5275), 
	.A(FE_PHN4941_n5275));
   BUF_X32 FE_PHC2446_n5262 (.Z(FE_PHN2446_n5262), 
	.A(FE_PHN5163_n5262));
   BUF_X32 FE_PHC2445_n5016 (.Z(FE_PHN2445_n5016), 
	.A(FE_PHN3906_n5016));
   BUF_X32 FE_PHC2444_n5390 (.Z(FE_PHN2444_n5390), 
	.A(FE_PHN4935_n5390));
   BUF_X32 FE_PHC2443_n5389 (.Z(FE_PHN2443_n5389), 
	.A(FE_PHN4822_n5389));
   BUF_X32 FE_PHC2442_n5495 (.Z(FE_PHN2442_n5495), 
	.A(FE_PHN4898_n5495));
   BUF_X32 FE_PHC2441_n5210 (.Z(FE_PHN2441_n5210), 
	.A(FE_PHN4911_n5210));
   BUF_X32 FE_PHC2440_n5307 (.Z(FE_PHN2440_n5307), 
	.A(FE_PHN5013_n5307));
   BUF_X32 FE_PHC2439_n5340 (.Z(FE_PHN2439_n5340), 
	.A(FE_PHN4807_n5340));
   BUF_X32 FE_PHC2438_n5073 (.Z(FE_PHN2438_n5073), 
	.A(FE_PHN4956_n5073));
   BUF_X32 FE_PHC2437_n5204 (.Z(FE_PHN2437_n5204), 
	.A(FE_PHN5105_n5204));
   BUF_X32 FE_PHC2436_n5577 (.Z(FE_PHN2436_n5577), 
	.A(FE_PHN4840_n5577));
   BUF_X32 FE_PHC2435_n5265 (.Z(FE_PHN2435_n5265), 
	.A(FE_PHN4767_n5265));
   BUF_X32 FE_PHC2430_n5520 (.Z(FE_PHN2430_n5520), 
	.A(n5520));
   BUF_X32 FE_PHC2429_n5505 (.Z(FE_PHN2429_n5505), 
	.A(n5505));
   BUF_X32 FE_PHC2428_n5507 (.Z(FE_PHN2428_n5507), 
	.A(n5507));
   BUF_X32 FE_PHC2426_n5581 (.Z(FE_PHN2426_n5581), 
	.A(n5581));
   BUF_X32 FE_PHC2420_n5652 (.Z(FE_PHN2420_n5652), 
	.A(FE_PHN4607_n5652));
   BUF_X8 FE_PHC2415_n5792 (.Z(FE_PHN2415_n5792), 
	.A(n5792));
   BUF_X32 FE_PHC2412_n5512 (.Z(FE_PHN2412_n5512), 
	.A(n5512));
   CLKBUF_X1 FE_PHC2403_n5711 (.Z(FE_PHN2403_n5711), 
	.A(n5711));
   BUF_X32 FE_PHC2385_n5625 (.Z(FE_PHN2385_n5625), 
	.A(n5625));
   BUF_X8 FE_PHC2379_n5793 (.Z(FE_PHN2379_n5793), 
	.A(n5793));
   BUF_X32 FE_PHC2378_n5618 (.Z(FE_PHN2378_n5618), 
	.A(n5618));
   BUF_X32 FE_PHC2376_n5571 (.Z(FE_PHN2376_n5571), 
	.A(n5571));
   BUF_X32 FE_PHC2364_n5639 (.Z(FE_PHN2364_n5639), 
	.A(n5639));
   BUF_X16 FE_PHC2355_U594_Z_0 (.Z(FE_PHN2355_U594_Z_0), 
	.A(U594_Z_0));
   BUF_X8 FE_PHC2348_n5790 (.Z(FE_PHN2348_n5790), 
	.A(n5790));
   BUF_X32 FE_PHC2347_n5513 (.Z(FE_PHN2347_n5513), 
	.A(n5513));
   BUF_X32 FE_PHC2346_U243_Z_0 (.Z(FE_PHN2346_U243_Z_0), 
	.A(FE_PHN4174_U243_Z_0));
   BUF_X32 FE_PHC2333_n5600 (.Z(FE_PHN2333_n5600), 
	.A(FE_PHN4439_n5600));
   BUF_X32 FE_PHC2330_n5579 (.Z(FE_PHN2330_n5579), 
	.A(FE_PHN4433_n5579));
   BUF_X32 FE_PHC2302_n5509 (.Z(FE_PHN2302_n5509), 
	.A(FE_PHN4337_n5509));
   BUF_X32 FE_PHC2300_U239_Z_0 (.Z(FE_PHN2300_U239_Z_0), 
	.A(FE_PHN3885_U239_Z_0));
   BUF_X16 FE_PHC2294_U325_Z_0 (.Z(FE_PHN2294_U325_Z_0), 
	.A(FE_PHN4797_U325_Z_0));
   BUF_X16 FE_PHC2286_U329_Z_0 (.Z(FE_PHN2286_U329_Z_0), 
	.A(FE_PHN3925_U329_Z_0));
   BUF_X32 FE_PHC2270_n5067 (.Z(FE_PHN2270_n5067), 
	.A(FE_PHN4416_n5067));
   BUF_X32 FE_PHC2254_n5074 (.Z(FE_PHN2254_n5074), 
	.A(FE_PHN4364_n5074));
   BUF_X32 FE_PHC2245_n5033 (.Z(FE_PHN2245_n5033), 
	.A(FE_PHN4402_n5033));
   BUF_X32 FE_PHC2241_U234_Z_0 (.Z(FE_PHN2241_U234_Z_0), 
	.A(FE_PHN4991_U234_Z_0));
   BUF_X32 FE_PHC2240_n5514 (.Z(FE_PHN2240_n5514), 
	.A(FE_PHN4216_n5514));
   BUF_X32 FE_PHC2233_U624_Z_0 (.Z(FE_PHN2233_U624_Z_0), 
	.A(FE_PHN3904_U624_Z_0));
   BUF_X32 FE_PHC2232_n5511 (.Z(FE_PHN2232_n5511), 
	.A(FE_PHN5050_n5511));
   BUF_X32 FE_PHC2225_U619_Z_0 (.Z(FE_PHN2225_U619_Z_0), 
	.A(FE_PHN4907_U619_Z_0));
   BUF_X32 FE_PHC2224_U628_Z_0 (.Z(FE_PHN2224_U628_Z_0), 
	.A(FE_PHN4772_U628_Z_0));
   BUF_X32 FE_PHC2223_n5508 (.Z(FE_PHN2223_n5508), 
	.A(FE_PHN5000_n5508));
   BUF_X32 FE_PHC2219_U585_Z_0 (.Z(FE_PHN2219_U585_Z_0), 
	.A(FE_PHN4864_U585_Z_0));
   BUF_X32 FE_PHC2215_U242_Z_0 (.Z(FE_PHN2215_U242_Z_0), 
	.A(FE_PHN4820_U242_Z_0));
   BUF_X32 FE_PHC2212_U233_Z_0 (.Z(FE_PHN2212_U233_Z_0), 
	.A(FE_PHN3763_U233_Z_0));
   BUF_X16 FE_PHC2210_U320_Z_0 (.Z(FE_PHN2210_U320_Z_0), 
	.A(U320_Z_0));
   BUF_X32 FE_PHC2200_U593_Z_0 (.Z(FE_PHN2200_U593_Z_0), 
	.A(U593_Z_0));
   BUF_X32 FE_PHC2196_U245_Z_0 (.Z(FE_PHN2196_U245_Z_0), 
	.A(U245_Z_0));
   BUF_X32 FE_PHC2189_U620_Z_0 (.Z(FE_PHN2189_U620_Z_0), 
	.A(U620_Z_0));
   BUF_X32 FE_PHC2187_U618_Z_0 (.Z(FE_PHN2187_U618_Z_0), 
	.A(U618_Z_0));
   BUF_X32 FE_PHC2181_U584_Z_0 (.Z(FE_PHN2181_U584_Z_0), 
	.A(U584_Z_0));
   BUF_X32 FE_PHC2180_n5517 (.Z(FE_PHN2180_n5517), 
	.A(FE_PHN4132_n5517));
   BUF_X16 FE_PHC2179_U627_Z_0 (.Z(FE_PHN2179_U627_Z_0), 
	.A(U627_Z_0));
   BUF_X32 FE_PHC2166_U596_Z_0 (.Z(FE_PHN2166_U596_Z_0), 
	.A(U596_Z_0));
   BUF_X32 FE_PHC2164_n4863 (.Z(FE_PHN2164_n4863), 
	.A(n4863));
   BUF_X32 FE_PHC2163_U332_Z_0 (.Z(FE_PHN2163_U332_Z_0), 
	.A(U332_Z_0));
   BUF_X32 FE_PHC2157_U328_Z_0 (.Z(FE_PHN2157_U328_Z_0), 
	.A(U328_Z_0));
   BUF_X32 FE_PHC2156_U311_Z_0 (.Z(FE_PHN2156_U311_Z_0), 
	.A(U311_Z_0));
   BUF_X32 FE_PHC2154_U302_Z_0 (.Z(FE_PHN2154_U302_Z_0), 
	.A(U302_Z_0));
   BUF_X32 FE_PHC2150_U310_Z_0 (.Z(FE_PHN2150_U310_Z_0), 
	.A(U310_Z_0));
   BUF_X32 FE_PHC2149_U621_Z_0 (.Z(FE_PHN2149_U621_Z_0), 
	.A(U621_Z_0));
   BUF_X16 FE_PHC2148_U597_Z_0 (.Z(FE_PHN2148_U597_Z_0), 
	.A(U597_Z_0));
   BUF_X32 FE_PHC2145_U303_Z_0 (.Z(FE_PHN2145_U303_Z_0), 
	.A(U303_Z_0));
   BUF_X32 FE_PHC2143_U631_Z_0 (.Z(FE_PHN2143_U631_Z_0), 
	.A(U631_Z_0));
   BUF_X32 FE_PHC2141_U301_Z_0 (.Z(FE_PHN2141_U301_Z_0), 
	.A(U301_Z_0));
   BUF_X32 FE_PHC2140_n5515 (.Z(FE_PHN2140_n5515), 
	.A(FE_PHN4949_n5515));
   BUF_X32 FE_PHC2125_U236_Z_0 (.Z(FE_PHN2125_U236_Z_0), 
	.A(U236_Z_0));
   BUF_X32 FE_PHC2120_U322_Z_0 (.Z(FE_PHN2120_U322_Z_0), 
	.A(U322_Z_0));
   BUF_X16 FE_PHC2114_U586_Z_0 (.Z(FE_PHN2114_U586_Z_0), 
	.A(U586_Z_0));
   BUF_X16 FE_PHC2109_U235_Z_0 (.Z(FE_PHN2109_U235_Z_0), 
	.A(U235_Z_0));
   BUF_X32 FE_PHC2107_U300_Z_0 (.Z(FE_PHN2107_U300_Z_0), 
	.A(U300_Z_0));
   BUF_X32 FE_PHC2106_n5506 (.Z(FE_PHN2106_n5506), 
	.A(FE_PHN4867_n5506));
   BUF_X16 FE_PHC2105_U519_Z_0 (.Z(FE_PHN2105_U519_Z_0), 
	.A(U519_Z_0));
   BUF_X32 FE_PHC2104_U524_Z_0 (.Z(FE_PHN2104_U524_Z_0), 
	.A(U524_Z_0));
   BUF_X32 FE_PHC2103_U314_Z_0 (.Z(FE_PHN2103_U314_Z_0), 
	.A(U314_Z_0));
   BUF_X32 FE_PHC2102_U331_Z_0 (.Z(FE_PHN2102_U331_Z_0), 
	.A(U331_Z_0));
   BUF_X16 FE_PHC2101_U246_Z_0 (.Z(FE_PHN2101_U246_Z_0), 
	.A(U246_Z_0));
   BUF_X32 FE_PHC2100_U592_Z_0 (.Z(FE_PHN2100_U592_Z_0), 
	.A(U592_Z_0));
   BUF_X16 FE_PHC2099_U321_Z_0 (.Z(FE_PHN2099_U321_Z_0), 
	.A(U321_Z_0));
   BUF_X32 FE_PHC2098_U587_Z_0 (.Z(FE_PHN2098_U587_Z_0), 
	.A(U587_Z_0));
   BUF_X32 FE_PHC2097_U626_Z_0 (.Z(FE_PHN2097_U626_Z_0), 
	.A(U626_Z_0));
   BUF_X32 FE_PHC2096_U326_Z_0 (.Z(FE_PHN2096_U326_Z_0), 
	.A(U326_Z_0));
   BUF_X32 FE_PHC2095_U629_Z_0 (.Z(FE_PHN2095_U629_Z_0), 
	.A(U629_Z_0));
   BUF_X32 FE_PHC2094_U306_Z_0 (.Z(FE_PHN2094_U306_Z_0), 
	.A(U306_Z_0));
   BUF_X16 FE_PHC2093_U632_Z_0 (.Z(FE_PHN2093_U632_Z_0), 
	.A(U632_Z_0));
   BUF_X32 FE_PHC2092_U534_Z_0 (.Z(FE_PHN2092_U534_Z_0), 
	.A(U534_Z_0));
   BUF_X32 FE_PHC2091_U232_Z_0 (.Z(FE_PHN2091_U232_Z_0), 
	.A(U232_Z_0));
   BUF_X32 FE_PHC2090_U307_Z_0 (.Z(FE_PHN2090_U307_Z_0), 
	.A(U307_Z_0));
   BUF_X32 FE_PHC2089_U565_Z_0 (.Z(FE_PHN2089_U565_Z_0), 
	.A(U565_Z_0));
   BUF_X16 FE_PHC2088_U583_Z_0 (.Z(FE_PHN2088_U583_Z_0), 
	.A(U583_Z_0));
   BUF_X32 FE_PHC2087_U617_Z_0 (.Z(FE_PHN2087_U617_Z_0), 
	.A(U617_Z_0));
   BUF_X32 FE_PHC2086_n4882 (.Z(FE_PHN2086_n4882), 
	.A(n4882));
   BUF_X16 FE_PHC2085_U591_Z_0 (.Z(FE_PHN2085_U591_Z_0), 
	.A(U591_Z_0));
   BUF_X32 FE_PHC2084_U238_Z_0 (.Z(FE_PHN2084_U238_Z_0), 
	.A(U238_Z_0));
   BUF_X32 FE_PHC2083_U327_Z_0 (.Z(FE_PHN2083_U327_Z_0), 
	.A(U327_Z_0));
   BUF_X32 FE_PHC2082_U532_Z_0 (.Z(FE_PHN2082_U532_Z_0), 
	.A(U532_Z_0));
   BUF_X32 FE_PHC2081_U623_Z_0 (.Z(FE_PHN2081_U623_Z_0), 
	.A(U623_Z_0));
   BUF_X32 FE_PHC2080_U622_Z_0 (.Z(FE_PHN2080_U622_Z_0), 
	.A(U622_Z_0));
   BUF_X32 FE_PHC2079_U523_Z_0 (.Z(FE_PHN2079_U523_Z_0), 
	.A(U523_Z_0));
   BUF_X32 FE_PHC2078_U312_Z_0 (.Z(FE_PHN2078_U312_Z_0), 
	.A(U312_Z_0));
   BUF_X32 FE_PHC2077_U555_Z_0 (.Z(FE_PHN2077_U555_Z_0), 
	.A(U555_Z_0));
   BUF_X32 FE_PHC2076_U564_Z_0 (.Z(FE_PHN2076_U564_Z_0), 
	.A(U564_Z_0));
   BUF_X32 FE_PHC2075_U333_Z_0 (.Z(FE_PHN2075_U333_Z_0), 
	.A(U333_Z_0));
   BUF_X16 FE_PHC2074_U557_Z_0 (.Z(FE_PHN2074_U557_Z_0), 
	.A(U557_Z_0));
   BUF_X32 FE_PHC2073_U240_Z_0 (.Z(FE_PHN2073_U240_Z_0), 
	.A(U240_Z_0));
   BUF_X16 FE_PHC2072_U324_Z_0 (.Z(FE_PHN2072_U324_Z_0), 
	.A(U324_Z_0));
   BUF_X32 FE_PHC2071_U237_Z_0 (.Z(FE_PHN2071_U237_Z_0), 
	.A(U237_Z_0));
   BUF_X32 FE_PHC2070_U625_Z_0 (.Z(FE_PHN2070_U625_Z_0), 
	.A(U625_Z_0));
   BUF_X16 FE_PHC2069_U589_Z_0 (.Z(FE_PHN2069_U589_Z_0), 
	.A(U589_Z_0));
   BUF_X32 FE_PHC2068_U330_Z_0 (.Z(FE_PHN2068_U330_Z_0), 
	.A(U330_Z_0));
   BUF_X32 FE_PHC2067_U588_Z_0 (.Z(FE_PHN2067_U588_Z_0), 
	.A(U588_Z_0));
   BUF_X16 FE_PHC2066_U305_Z_0 (.Z(FE_PHN2066_U305_Z_0), 
	.A(U305_Z_0));
   BUF_X32 FE_PHC2065_U556_Z_0 (.Z(FE_PHN2065_U556_Z_0), 
	.A(U556_Z_0));
   BUF_X32 FE_PHC2064_U308_Z_0 (.Z(FE_PHN2064_U308_Z_0), 
	.A(U308_Z_0));
   BUF_X32 FE_PHC2063_U598_Z_0 (.Z(FE_PHN2063_U598_Z_0), 
	.A(U598_Z_0));
   BUF_X16 FE_PHC2062_U595_Z_0 (.Z(FE_PHN2062_U595_Z_0), 
	.A(U595_Z_0));
   BUF_X32 FE_PHC2061_U304_Z_0 (.Z(FE_PHN2061_U304_Z_0), 
	.A(U304_Z_0));
   BUF_X16 FE_PHC2060_U318_Z_0 (.Z(FE_PHN2060_U318_Z_0), 
	.A(U318_Z_0));
   BUF_X16 FE_PHC2059_U563_Z_0 (.Z(FE_PHN2059_U563_Z_0), 
	.A(U563_Z_0));
   BUF_X16 FE_PHC2058_U309_Z_0 (.Z(FE_PHN2058_U309_Z_0), 
	.A(U309_Z_0));
   BUF_X16 FE_PHC2057_U528_Z_0 (.Z(FE_PHN2057_U528_Z_0), 
	.A(U528_Z_0));
   BUF_X16 FE_PHC2056_U323_Z_0 (.Z(FE_PHN2056_U323_Z_0), 
	.A(U323_Z_0));
   BUF_X32 FE_PHC2055_U241_Z_0 (.Z(FE_PHN2055_U241_Z_0), 
	.A(U241_Z_0));
   BUF_X32 FE_PHC2054_U533_Z_0 (.Z(FE_PHN2054_U533_Z_0), 
	.A(U533_Z_0));
   BUF_X32 FE_PHC2053_U315_Z_0 (.Z(FE_PHN2053_U315_Z_0), 
	.A(U315_Z_0));
   BUF_X32 FE_PHC2052_U244_Z_0 (.Z(FE_PHN2052_U244_Z_0), 
	.A(U244_Z_0));
   CLKBUF_X1 FE_PHC2050_n5694 (.Z(FE_PHN2050_n5694), 
	.A(n5694));
   CLKBUF_X1 FE_PHC2049_n222 (.Z(FE_PHN2049_n222), 
	.A(n222));
   BUF_X16 FE_PHC2048_n227 (.Z(FE_PHN2048_n227), 
	.A(n227));
   BUF_X16 FE_PHC2047_n216 (.Z(FE_PHN2047_n216), 
	.A(n216));
   BUF_X16 FE_PHC2046_n5699 (.Z(FE_PHN2046_n5699), 
	.A(n5699));
   BUF_X32 FE_PHC2045_n1000 (.Z(FE_PHN2045_n1000), 
	.A(n1000));
   BUF_X32 FE_PHC2043_n230 (.Z(FE_PHN2043_n230), 
	.A(n230));
   BUF_X32 FE_PHC2042_n1051 (.Z(FE_PHN2042_n1051), 
	.A(n1051));
   BUF_X32 FE_PHC2041_n220 (.Z(FE_PHN2041_n220), 
	.A(n220));
   BUF_X16 FE_PHC2039_U144_Z_0 (.Z(FE_PHN2039_U144_Z_0), 
	.A(U144_Z_0));
   BUF_X32 FE_PHC2035_n214 (.Z(FE_PHN2035_n214), 
	.A(FE_PHN3466_n214));
   BUF_X8 FE_PHC2028_n5776 (.Z(FE_PHN2028_n5776), 
	.A(n5776));
   BUF_X32 FE_PHC1983_n4923 (.Z(FE_PHN1983_n4923), 
	.A(FE_PHN4712_n4923));
   BUF_X4 FE_PHC1978_n4938 (.Z(FE_PHN1978_n4938), 
	.A(n4938));
   BUF_X32 FE_PHC1970_U754_Z_0 (.Z(FE_PHN1970_U754_Z_0), 
	.A(FE_PHN3796_U754_Z_0));
   BUF_X32 FE_PHC1967_U122_Z_0 (.Z(FE_PHN1967_U122_Z_0), 
	.A(U122_Z_0));
   CLKBUF_X1 FE_PHC1934_n4924 (.Z(FE_PHN1934_n4924), 
	.A(n4924));
   BUF_X4 FE_PHC1920_n4935 (.Z(FE_PHN1920_n4935), 
	.A(n4935));
   CLKBUF_X1 FE_PHC1919_n5712 (.Z(FE_PHN1919_n5712), 
	.A(n5712));
   BUF_X4 FE_PHC1915_n4936 (.Z(FE_PHN1915_n4936), 
	.A(n4936));
   BUF_X4 FE_PHC1914_n4942 (.Z(FE_PHN1914_n4942), 
	.A(n4942));
   BUF_X4 FE_PHC1912_n4926 (.Z(FE_PHN1912_n4926), 
	.A(n4926));
   CLKBUF_X1 FE_PHC1910_n4937 (.Z(FE_PHN1910_n4937), 
	.A(n4937));
   CLKBUF_X1 FE_PHC1909_n4931 (.Z(FE_PHN1909_n4931), 
	.A(n4931));
   CLKBUF_X1 FE_PHC1908_n4925 (.Z(FE_PHN1908_n4925), 
	.A(n4925));
   BUF_X32 FE_PHC1906_n5800 (.Z(FE_PHN1906_n5800), 
	.A(FE_PHN3273_n5800));
   BUF_X16 FE_PHC1905_n5828 (.Z(FE_PHN1905_n5828), 
	.A(n5828));
   BUF_X32 FE_PHC1903_n5795 (.Z(FE_PHN1903_n5795), 
	.A(FE_PHN3470_n5795));
   BUF_X32 FE_PHC1902_n4903 (.Z(FE_PHN1902_n4903), 
	.A(FE_PHN4671_n4903));
   BUF_X32 FE_PHC1901_n4902 (.Z(FE_PHN1901_n4902), 
	.A(FE_PHN4675_n4902));
   BUF_X32 FE_PHC1900_n4324 (.Z(FE_PHN1900_n4324), 
	.A(FE_PHN4669_n4324));
   BUF_X32 FE_PHC1899_n4326 (.Z(FE_PHN1899_n4326), 
	.A(n4326));
   CLKBUF_X1 FE_PHC1898_U317_Z_0 (.Z(FE_PHN1898_U317_Z_0), 
	.A(U317_Z_0));
   CLKBUF_X1 FE_PHC1894_n5149 (.Z(FE_PHN1894_n5149), 
	.A(n5149));
   BUF_X16 FE_PHC1875_n5653 (.Z(FE_PHN1875_n5653), 
	.A(n5653));
   BUF_X32 FE_PHC1846_U590_Z_0 (.Z(FE_PHN1846_U590_Z_0), 
	.A(FE_PHN4212_U590_Z_0));
   BUF_X32 FE_PHC1809_n4874 (.Z(FE_PHN1809_n4874), 
	.A(FE_PHN5161_n4874));
   BUF_X16 FE_PHC1759_U630_Z_0 (.Z(FE_PHN1759_U630_Z_0), 
	.A(U630_Z_0));
   BUF_X16 FE_PHC1751_U319_Z_0 (.Z(FE_PHN1751_U319_Z_0), 
	.A(U319_Z_0));
   BUF_X32 FE_PHC1748_n5510 (.Z(FE_PHN1748_n5510), 
	.A(n5510));
   BUF_X32 FE_PHC1744_U531_Z_0 (.Z(FE_PHN1744_U531_Z_0), 
	.A(U531_Z_0));
   BUF_X32 FE_PHC1743_U313_Z_0 (.Z(FE_PHN1743_U313_Z_0), 
	.A(U313_Z_0));
   BUF_X16 FE_PHC1742_U566_Z_0 (.Z(FE_PHN1742_U566_Z_0), 
	.A(U566_Z_0));
   BUF_X16 FE_PHC1741_U247_Z_0 (.Z(FE_PHN1741_U247_Z_0), 
	.A(U247_Z_0));
   BUF_X32 FE_PHC1717_n5114 (.Z(FE_PHN1717_n5114), 
	.A(n5114));
   BUF_X32 FE_PHC1682_n16735 (.Z(FE_PHN1682_n16735), 
	.A(n16735));
   BUF_X32 FE_PHC1674_n13951 (.Z(FE_PHN1674_n13951), 
	.A(FE_PHN3202_n13951));
   BUF_X32 FE_PHC1673_n14956 (.Z(FE_PHN1673_n14956), 
	.A(FE_PHN3060_n14956));
   BUF_X32 FE_PHC1672_n13963 (.Z(FE_PHN1672_n13963), 
	.A(FE_PHN3066_n13963));
   BUF_X32 FE_PHC1671_n13870 (.Z(FE_PHN1671_n13870), 
	.A(FE_PHN3201_n13870));
   BUF_X32 FE_PHC1670_n13932 (.Z(FE_PHN1670_n13932), 
	.A(FE_PHN3065_n13932));
   BUF_X32 FE_PHC1669_n13894 (.Z(FE_PHN1669_n13894), 
	.A(FE_PHN3061_n13894));
   BUF_X32 FE_PHC1668_n4389 (.Z(FE_PHN1668_n4389), 
	.A(FE_PHN5193_n4389));
   BUF_X32 FE_PHC1667_n13989 (.Z(FE_PHN1667_n13989), 
	.A(FE_PHN3067_n13989));
   BUF_X32 FE_PHC1666_n13919 (.Z(FE_PHN1666_n13919), 
	.A(FE_PHN3063_n13919));
   BUF_X32 FE_PHC1665_n1127 (.Z(FE_PHN1665_n1127), 
	.A(n1127));
   BUF_X32 FE_PHC1664_n13747 (.Z(FE_PHN1664_n13747), 
	.A(n13747));
   BUF_X16 FE_PHC1657_n5779 (.Z(FE_PHN1657_n5779), 
	.A(n5779));
   BUF_X32 FE_PHC1655_n4860 (.Z(FE_PHN1655_n4860), 
	.A(n4860));
   BUF_X16 FE_PHC1654_U105_Z_0 (.Z(FE_PHN1654_U105_Z_0), 
	.A(U105_Z_0));
   BUF_X32 FE_PHC1653_U802_Z_0 (.Z(FE_PHN1653_U802_Z_0), 
	.A(FE_PHN4608_U802_Z_0));
   BUF_X16 FE_PHC1652_U134_Z_0 (.Z(FE_PHN1652_U134_Z_0), 
	.A(U134_Z_0));
   BUF_X16 FE_PHC1651_U121_Z_0 (.Z(FE_PHN1651_U121_Z_0), 
	.A(U121_Z_0));
   CLKBUF_X1 FE_PHC1649_U755_Z_0 (.Z(FE_PHN1649_U755_Z_0), 
	.A(U755_Z_0));
   CLKBUF_X1 FE_PHC1648_U811_Z_0 (.Z(FE_PHN1648_U811_Z_0), 
	.A(U811_Z_0));
   BUF_X32 FE_PHC1646_U518_Z_0 (.Z(FE_PHN1646_U518_Z_0), 
	.A(FE_PHN4590_U518_Z_0));
   BUF_X8 FE_PHC1644_U795_Z_0 (.Z(FE_PHN1644_U795_Z_0), 
	.A(U795_Z_0));
   BUF_X32 FE_PHC1636_n4878 (.Z(FE_PHN1636_n4878), 
	.A(FE_PHN5043_n4878));
   BUF_X16 FE_PHC1633_U98_Z_0 (.Z(FE_PHN1633_U98_Z_0), 
	.A(U98_Z_0));
   BUF_X16 FE_PHC1632_U97_Z_0 (.Z(FE_PHN1632_U97_Z_0), 
	.A(U97_Z_0));
   BUF_X32 FE_PHC1631_n4943 (.Z(FE_PHN1631_n4943), 
	.A(n4943));
   BUF_X32 FE_PHC1629_n5784 (.Z(FE_PHN1629_n5784), 
	.A(FE_PHN3608_n5784));
   BUF_X32 FE_PHC1627_n5786 (.Z(FE_PHN1627_n5786), 
	.A(n5786));
   BUF_X4 FE_PHC1626_n5736 (.Z(FE_PHN1626_n5736), 
	.A(n5736));
   BUF_X32 FE_PHC1625_n4864 (.Z(FE_PHN1625_n4864), 
	.A(n4864));
   BUF_X32 FE_PHC1624_n4881 (.Z(FE_PHN1624_n4881), 
	.A(n4881));
   BUF_X32 FE_PHC1615_n5827 (.Z(FE_PHN1615_n5827), 
	.A(FE_PHN3205_n5827));
   BUF_X32 FE_PHC1614_U665_Z_0 (.Z(FE_PHN1614_U665_Z_0), 
	.A(U665_Z_0));
   BUF_X32 FE_PHC1613_n5777 (.Z(FE_PHN1613_n5777), 
	.A(n5777));
   BUF_X32 FE_PHC1612_n5781 (.Z(FE_PHN1612_n5781), 
	.A(n5781));
   BUF_X32 FE_PHC1610_n4886 (.Z(FE_PHN1610_n4886), 
	.A(n4886));
   BUF_X32 FE_PHC1606_n13795 (.Z(FE_PHN1606_n13795), 
	.A(FE_PHN3068_n13795));
   BUF_X32 FE_PHC1603_n13813 (.Z(FE_PHN1603_n13813), 
	.A(FE_PHN3204_n13813));
   BUF_X32 FE_PHC1602_n13835 (.Z(FE_PHN1602_n13835), 
	.A(FE_PHN3064_n13835));
   BUF_X32 FE_PHC1601_n13758 (.Z(FE_PHN1601_n13758), 
	.A(FE_PHN3058_n13758));
   BUF_X32 FE_PHC1600_n13907 (.Z(FE_PHN1600_n13907), 
	.A(FE_PHN3059_n13907));
   BUF_X32 FE_PHC1599_n1431 (.Z(FE_PHN1599_n1431), 
	.A(n1431));
   BUF_X32 FE_PHC1598_n4328 (.Z(FE_PHN1598_n4328), 
	.A(n4328));
   CLKBUF_X1 FE_PHC1588_n5737 (.Z(FE_PHN1588_n5737), 
	.A(n5737));
   BUF_X32 FE_PHC1586_n5256 (.Z(FE_PHN1586_n5256), 
	.A(n5256));
   BUF_X4 FE_PHC1577_n5684 (.Z(FE_PHN1577_n5684), 
	.A(n5684));
   BUF_X16 FE_PHC1571_n5771 (.Z(FE_PHN1571_n5771), 
	.A(n5771));
   BUF_X16 FE_PHC1566_n8706 (.Z(FE_PHN1566_n8706), 
	.A(n8706));
   BUF_X16 FE_PHC1565_n8698 (.Z(FE_PHN1565_n8698), 
	.A(n8698));
   BUF_X4 FE_PHC1559_n5682 (.Z(FE_PHN1559_n5682), 
	.A(n5682));
   BUF_X32 FE_PHC1551_n1319 (.Z(FE_PHN1551_n1319), 
	.A(FE_PHN4288_n1319));
   BUF_X32 FE_PHC1538_n5772 (.Z(FE_PHN1538_n5772), 
	.A(n5772));
   BUF_X32 FE_PHC1512_n4331 (.Z(FE_PHN1512_n4331), 
	.A(n4331));
   CLKBUF_X1 FE_PHC1508_n10553 (.Z(FE_PHN1508_n10553), 
	.A(n10553));
   BUF_X32 FE_PHC1503_IRQ_14_ (.Z(FE_PHN1503_IRQ_14_), 
	.A(irq_i[14]));
   BUF_X32 FE_PHC1502_n11928 (.Z(FE_PHN1502_n11928), 
	.A(n11928));
   CLKBUF_X1 FE_PHC1501_n779 (.Z(FE_PHN1501_n779), 
	.A(n779));
   CLKBUF_X1 FE_PHC1500_n5785 (.Z(FE_PHN1500_n5785), 
	.A(n5785));
   CLKBUF_X1 FE_PHC1499_n5783 (.Z(FE_PHN1499_n5783), 
	.A(n5783));
   CLKBUF_X1 FE_PHC1490_n5787 (.Z(FE_PHN1490_n5787), 
	.A(n5787));
   BUF_X32 FE_PHC1488_U691_Z_0 (.Z(FE_PHN1488_U691_Z_0), 
	.A(FE_PHN4524_U691_Z_0));
   BUF_X4 FE_PHC1472_n5738 (.Z(FE_PHN1472_n5738), 
	.A(n5738));
   BUF_X32 FE_PHC1469_n4875 (.Z(FE_PHN1469_n4875), 
	.A(FE_PHN5141_n4875));
   BUF_X16 FE_PHC1468_n5662 (.Z(FE_PHN1468_n5662), 
	.A(n5662));
   BUF_X16 FE_PHC1463_n5665 (.Z(FE_PHN1463_n5665), 
	.A(n5665));
   BUF_X16 FE_PHC1462_n5660 (.Z(FE_PHN1462_n5660), 
	.A(n5660));
   BUF_X32 FE_PHC1461_n4944 (.Z(FE_PHN1461_n4944), 
	.A(n4944));
   BUF_X32 FE_PHC1457_n5654 (.Z(FE_PHN1457_n5654), 
	.A(n5654));
   CLKBUF_X1 FE_PHC1450_n5788 (.Z(FE_PHN1450_n5788), 
	.A(n5788));
   BUF_X4 FE_PHC1448_n5782 (.Z(FE_PHN1448_n5782), 
	.A(n5782));
   BUF_X32 FE_PHC1433_n5824 (.Z(FE_PHN1433_n5824), 
	.A(n5824));
   BUF_X32 FE_PHC1431_n5775 (.Z(FE_PHN1431_n5775), 
	.A(n5775));
   BUF_X32 FE_PHC1429_n4945 (.Z(FE_PHN1429_n4945), 
	.A(FE_PHN3069_n4945));
   CLKBUF_X1 FE_PHC1428_n5789 (.Z(FE_PHN1428_n5789), 
	.A(n5789));
   BUF_X32 FE_PHC1426_U227_Z_0 (.Z(FE_PHN1426_U227_Z_0), 
	.A(FE_PHN3143_U227_Z_0));
   BUF_X32 FE_PHC1425_n14001 (.Z(FE_PHN1425_n14001), 
	.A(FE_PHN3092_n14001));
   BUF_X32 FE_PHC1399_n5723 (.Z(FE_PHN1399_n5723), 
	.A(n5723));
   BUF_X32 FE_PHC1398_n5727 (.Z(FE_PHN1398_n5727), 
	.A(n5727));
   BUF_X32 FE_PHC1397_n5725 (.Z(FE_PHN1397_n5725), 
	.A(FE_PHN3610_n5725));
   BUF_X32 FE_PHC1396_n5730 (.Z(FE_PHN1396_n5730), 
	.A(FE_PHN3604_n5730));
   BUF_X32 FE_PHC1395_n5719 (.Z(FE_PHN1395_n5719), 
	.A(n5719));
   BUF_X32 FE_PHC1394_n5721 (.Z(FE_PHN1394_n5721), 
	.A(n5721));
   BUF_X32 FE_PHC1393_n5724 (.Z(FE_PHN1393_n5724), 
	.A(n5724));
   CLKBUF_X1 FE_PHC1392_n4932 (.Z(FE_PHN1392_n4932), 
	.A(n4932));
   CLKBUF_X1 FE_PHC1391_n4930 (.Z(FE_PHN1391_n4930), 
	.A(n4930));
   BUF_X32 FE_PHC1390_n4876 (.Z(FE_PHN1390_n4876), 
	.A(n4876));
   CLKBUF_X1 FE_PHC1389_n4934 (.Z(FE_PHN1389_n4934), 
	.A(n4934));
   CLKBUF_X1 FE_PHC1385_n4928 (.Z(FE_PHN1385_n4928), 
	.A(n4928));
   BUF_X32 FE_PHC1379_n5798 (.Z(FE_PHN1379_n5798), 
	.A(FE_PHN3074_n5798));
   BUF_X16 FE_PHC1377_n4879 (.Z(FE_PHN1377_n4879), 
	.A(n4879));
   CLKBUF_X1 FE_PHC1367_n4895 (.Z(FE_PHN1367_n4895), 
	.A(n4895));
   BUF_X32 FE_PHC1366_IRQ_8_ (.Z(FE_PHN1366_IRQ_8_), 
	.A(irq_i[8]));
   CLKBUF_X1 FE_PHC1365_IRQ_10_ (.Z(FE_PHN1365_IRQ_10_), 
	.A(irq_i[10]));
   BUF_X32 FE_PHC1364_n4896 (.Z(FE_PHN1364_n4896), 
	.A(n4896));
   CLKBUF_X1 FE_PHC1363_IRQ_4_ (.Z(FE_PHN1363_IRQ_4_), 
	.A(irq_i[4]));
   BUF_X32 FE_PHC1362_n4397 (.Z(FE_PHN1362_n4397), 
	.A(FE_PHN4667_n4397));
   CLKBUF_X1 FE_PHC1361_IRQ_7_ (.Z(FE_PHN1361_IRQ_7_), 
	.A(irq_i[7]));
   CLKBUF_X1 FE_PHC1360_IRQ_1_ (.Z(FE_PHN1360_IRQ_1_), 
	.A(irq_i[1]));
   CLKBUF_X1 FE_PHC1359_IRQ_13_ (.Z(FE_PHN1359_IRQ_13_), 
	.A(irq_i[13]));
   BUF_X32 FE_PHC1358_n4394 (.Z(FE_PHN1358_n4394), 
	.A(FE_PHN4674_n4394));
   CLKBUF_X1 FE_PHC1357_IRQ_5_ (.Z(FE_PHN1357_IRQ_5_), 
	.A(irq_i[5]));
   BUF_X32 FE_PHC1356_n4336 (.Z(FE_PHN1356_n4336), 
	.A(n4336));
   BUF_X2 FE_PHC1355_IRQ_0_ (.Z(FE_PHN1355_IRQ_0_), 
	.A(irq_i[0]));
   BUF_X32 FE_PHC1354_n4190 (.Z(FE_PHN1354_n4190), 
	.A(FE_PHN4666_n4190));
   CLKBUF_X1 FE_PHC1353_IRQ_6_ (.Z(FE_PHN1353_IRQ_6_), 
	.A(irq_i[6]));
   BUF_X32 FE_PHC1352_n4391 (.Z(FE_PHN1352_n4391), 
	.A(FE_PHN4668_n4391));
   CLKBUF_X1 FE_PHC1351_IRQ_11_ (.Z(FE_PHN1351_IRQ_11_), 
	.A(irq_i[11]));
   BUF_X2 FE_PHC1350_IRQ_15_ (.Z(FE_PHN1350_IRQ_15_), 
	.A(irq_i[15]));
   CLKBUF_X1 FE_PHC1349_IRQ_2_ (.Z(FE_PHN1349_IRQ_2_), 
	.A(irq_i[2]));
   BUF_X32 FE_PHC1348_n4300 (.Z(FE_PHN1348_n4300), 
	.A(FE_PHN4672_n4300));
   BUF_X2 FE_PHC1347_NMI (.Z(FE_PHN1347_NMI), 
	.A(nmi_i));
   CLKBUF_X1 FE_PHC1346_IRQ_9_ (.Z(FE_PHN1346_IRQ_9_), 
	.A(irq_i[9]));
   CLKBUF_X1 FE_PHC1345_IRQ_3_ (.Z(FE_PHN1345_IRQ_3_), 
	.A(irq_i[3]));
   BUF_X32 FE_PHC1344_n4193 (.Z(FE_PHN1344_n4193), 
	.A(FE_PHN4670_n4193));
   BUF_X32 FE_PHC1341_SYNOPSYS_UNCONNECTED_531 (.Z(FE_PHN1341_SYNOPSYS_UNCONNECTED_531), 
	.A(vis_pc_o[14]));
   BUF_X32 FE_PHC1339_SYNOPSYS_UNCONNECTED_540 (.Z(FE_PHN1339_SYNOPSYS_UNCONNECTED_540), 
	.A(vis_pc_o[5]));
   BUF_X32 FE_PHC1331_SYNOPSYS_UNCONNECTED_522 (.Z(FE_PHN1331_SYNOPSYS_UNCONNECTED_522), 
	.A(vis_pc_o[23]));
   BUF_X32 FE_PHC1320_SYNOPSYS_UNCONNECTED_518 (.Z(FE_PHN1320_SYNOPSYS_UNCONNECTED_518), 
	.A(vis_pc_o[27]));
   BUF_X16 FE_PHC1283_n5770 (.Z(FE_PHN1283_n5770), 
	.A(n5770));
   BUF_X16 FE_PHC1255_n5735 (.Z(FE_PHN1255_n5735), 
	.A(n5735));
   BUF_X32 FE_PHC1241_U229_Z_0 (.Z(FE_PHN1241_U229_Z_0), 
	.A(FE_PHN3211_U229_Z_0));
   BUF_X32 FE_PHC1237_U809_Z_0 (.Z(FE_PHN1237_U809_Z_0), 
	.A(U809_Z_0));
   BUF_X16 FE_PHC1196_n5664 (.Z(FE_PHN1196_n5664), 
	.A(n5664));
   BUF_X16 FE_PHC1195_n5663 (.Z(FE_PHN1195_n5663), 
	.A(n5663));
   BUF_X16 FE_PHC1183_n5659 (.Z(FE_PHN1183_n5659), 
	.A(n5659));
   CLKBUF_X1 FE_PHC1177_n4929 (.Z(FE_PHN1177_n4929), 
	.A(n4929));
   CLKBUF_X1 FE_PHC1175_n4933 (.Z(FE_PHN1175_n4933), 
	.A(n4933));
   CLKBUF_X1 FE_PHC1174_n4939 (.Z(FE_PHN1174_n4939), 
	.A(n4939));
   BUF_X32 FE_PHC1172_n5826 (.Z(FE_PHN1172_n5826), 
	.A(FE_PHN3472_n5826));
   BUF_X32 FE_PHC1164_n1444 (.Z(FE_PHN1164_n1444), 
	.A(n1444));
   BUF_X8 FE_PHC1159_n5676 (.Z(FE_PHN1159_n5676), 
	.A(n5676));
   BUF_X16 FE_PHC1157_n5823 (.Z(FE_PHN1157_n5823), 
	.A(n5823));
   BUF_X16 FE_PHC1145_n5729 (.Z(FE_PHN1145_n5729), 
	.A(n5729));
   BUF_X16 FE_PHC1142_n5733 (.Z(FE_PHN1142_n5733), 
	.A(n5733));
   BUF_X16 FE_PHC1141_n5713 (.Z(FE_PHN1141_n5713), 
	.A(n5713));
   BUF_X16 FE_PHC1139_n5734 (.Z(FE_PHN1139_n5734), 
	.A(n5734));
   BUF_X32 FE_PHC1138_n5715 (.Z(FE_PHN1138_n5715), 
	.A(n5715));
   BUF_X32 FE_PHC1137_n5732 (.Z(FE_PHN1137_n5732), 
	.A(FE_PHN3625_n5732));
   BUF_X32 FE_PHC1136_n5731 (.Z(FE_PHN1136_n5731), 
	.A(FE_PHN3612_n5731));
   BUF_X32 FE_PHC1135_n5722 (.Z(FE_PHN1135_n5722), 
	.A(n5722));
   BUF_X16 FE_PHC1134_n5716 (.Z(FE_PHN1134_n5716), 
	.A(n5716));
   BUF_X16 FE_PHC1133_n5728 (.Z(FE_PHN1133_n5728), 
	.A(n5728));
   BUF_X32 FE_PHC1131_n5718 (.Z(FE_PHN1131_n5718), 
	.A(n5718));
   BUF_X32 FE_PHC1130_n5726 (.Z(FE_PHN1130_n5726), 
	.A(FE_PHN3591_n5726));
   BUF_X32 FE_PHC1129_n5714 (.Z(FE_PHN1129_n5714), 
	.A(FE_PHN3592_n5714));
   BUF_X16 FE_PHC1128_n5717 (.Z(FE_PHN1128_n5717), 
	.A(n5717));
   BUF_X32 FE_PHC1126_U692_Z_0 (.Z(FE_PHN1126_U692_Z_0), 
	.A(FE_PHN4905_U692_Z_0));
   BUF_X16 FE_PHC1086_n5661 (.Z(FE_PHN1086_n5661), 
	.A(n5661));
   BUF_X32 FE_PHC1085_n5720 (.Z(FE_PHN1085_n5720), 
	.A(FE_PHN3595_n5720));
   BUF_X32 FE_PHC1078_n5668 (.Z(FE_PHN1078_n5668), 
	.A(n5668));
   CLKBUF_X1 FE_PHC1063_n5667 (.Z(FE_PHN1063_n5667), 
	.A(n5667));
   BUF_X16 FE_PHC1038_n5761 (.Z(FE_PHN1038_n5761), 
	.A(n5761));
   CLKBUF_X1 FE_PHC1037_n5007 (.Z(FE_PHN1037_n5007), 
	.A(n5007));
   BUF_X32 FE_PHC1025_n3063 (.Z(FE_PHN1025_n3063), 
	.A(n3063));
   BUF_X4 FE_PHC1024_n5690 (.Z(FE_PHN1024_n5690), 
	.A(n5690));
   BUF_X4 FE_PHC1010_n5766 (.Z(FE_PHN1010_n5766), 
	.A(n5766));
   BUF_X4 FE_PHC1009_n5765 (.Z(FE_PHN1009_n5765), 
	.A(n5765));
   BUF_X4 FE_PHC1008_n5767 (.Z(FE_PHN1008_n5767), 
	.A(n5767));
   BUF_X4 FE_PHC1007_n5768 (.Z(FE_PHN1007_n5768), 
	.A(n5768));
   BUF_X4 FE_PHC1006_n5769 (.Z(FE_PHN1006_n5769), 
	.A(n5769));
   BUF_X32 FE_PHC1005_n5764 (.Z(FE_PHN1005_n5764), 
	.A(n5764));
   BUF_X4 FE_PHC1004_n5673 (.Z(FE_PHN1004_n5673), 
	.A(n5673));
   BUF_X4 FE_PHC1003_n5675 (.Z(FE_PHN1003_n5675), 
	.A(n5675));
   BUF_X8 FE_PHC991_n5679 (.Z(FE_PHN991_n5679), 
	.A(n5679));
   BUF_X32 FE_PHC972_n5755 (.Z(FE_PHN972_n5755), 
	.A(FE_PHN3139_n5755));
   CLKBUF_X1 FE_PHC965_n5658 (.Z(FE_PHN965_n5658), 
	.A(n5658));
   BUF_X16 FE_PHC963_n5671 (.Z(FE_PHN963_n5671), 
	.A(n5671));
   BUF_X8 FE_PHC946_n5677 (.Z(FE_PHN946_n5677), 
	.A(n5677));
   BUF_X16 FE_PHC941_n5674 (.Z(FE_PHN941_n5674), 
	.A(n5674));
   CLKBUF_X1 FE_PHC939_n5680 (.Z(FE_PHN939_n5680), 
	.A(n5680));
   CLKBUF_X1 FE_PHC936_n5683 (.Z(FE_PHN936_n5683), 
	.A(n5683));
   BUF_X32 FE_PHC935_n2982 (.Z(FE_PHN935_n2982), 
	.A(n2982));
   BUF_X16 FE_PHC928_n14432 (.Z(FE_PHN928_n14432), 
	.A(n14432));
   CLKBUF_X1 FE_PHC904_n393 (.Z(FE_PHN904_n393), 
	.A(n393));
   BUF_X16 FE_PHC892_n14928 (.Z(FE_PHN892_n14928), 
	.A(n14928));
   CLKBUF_X1 FE_PHC875_n423 (.Z(FE_PHN875_n423), 
	.A(n423));
   CLKBUF_X1 FE_PHC870_n420 (.Z(FE_PHN870_n420), 
	.A(n420));
   BUF_X32 FE_PHC869_n427 (.Z(FE_PHN869_n427), 
	.A(n427));
   BUF_X32 FE_PHC859_n2624 (.Z(FE_PHN859_n2624), 
	.A(n2624));
   BUF_X16 FE_PHC856_n5656 (.Z(FE_PHN856_n5656), 
	.A(n5656));
   BUF_X16 FE_PHC852_n5763 (.Z(FE_PHN852_n5763), 
	.A(n5763));
   BUF_X32 FE_PHC851_n4920 (.Z(FE_PHN851_n4920), 
	.A(FE_PHN2967_n4920));
   BUF_X32 FE_PHC849_n4918 (.Z(FE_PHN849_n4918), 
	.A(FE_PHN3093_n4918));
   BUF_X32 FE_PHC847_n4917 (.Z(FE_PHN847_n4917), 
	.A(FE_PHN2969_n4917));
   BUF_X16 FE_PHC846_n4915 (.Z(FE_PHN846_n4915), 
	.A(n4915));
   BUF_X32 FE_PHC845_n4919 (.Z(FE_PHN845_n4919), 
	.A(FE_PHN2968_n4919));
   CLKBUF_X1 FE_PHC844_n425 (.Z(FE_PHN844_n425), 
	.A(n425));
   BUF_X32 FE_PHC839_n5678 (.Z(FE_PHN839_n5678), 
	.A(n5678));
   BUF_X16 FE_PHC830_n5760 (.Z(FE_PHN830_n5760), 
	.A(n5760));
   BUF_X16 FE_PHC829_n5756 (.Z(FE_PHN829_n5756), 
	.A(n5756));
   BUF_X32 FE_PHC826_n4921 (.Z(FE_PHN826_n4921), 
	.A(FE_PHN3140_n4921));
   BUF_X32 FE_PHC825_n4913 (.Z(FE_PHN825_n4913), 
	.A(FE_PHN2946_n4913));
   BUF_X32 FE_PHC824_n4908 (.Z(FE_PHN824_n4908), 
	.A(FE_PHN2973_n4908));
   BUF_X32 FE_PHC823_n4914 (.Z(FE_PHN823_n4914), 
	.A(FE_PHN3135_n4914));
   BUF_X32 FE_PHC822_n4910 (.Z(FE_PHN822_n4910), 
	.A(FE_PHN3137_n4910));
   BUF_X32 FE_PHC821_n4911 (.Z(FE_PHN821_n4911), 
	.A(FE_PHN2947_n4911));
   BUF_X32 FE_PHC820_n4916 (.Z(FE_PHN820_n4916), 
	.A(FE_PHN2951_n4916));
   BUF_X16 FE_PHC819_n4909 (.Z(FE_PHN819_n4909), 
	.A(n4909));
   BUF_X16 FE_PHC818_n4912 (.Z(FE_PHN818_n4912), 
	.A(n4912));
   BUF_X16 FE_PHC813_n5670 (.Z(FE_PHN813_n5670), 
	.A(n5670));
   CLKBUF_X1 FE_PHC806_n1143 (.Z(FE_PHN806_n1143), 
	.A(n1143));
   CLKBUF_X1 FE_PHC804_n429 (.Z(FE_PHN804_n429), 
	.A(n429));
   BUF_X32 FE_PHC803_n5757 (.Z(FE_PHN803_n5757), 
	.A(n5757));
   BUF_X16 FE_PHC802_n5762 (.Z(FE_PHN802_n5762), 
	.A(n5762));
   BUF_X32 FE_PHC801_n5758 (.Z(FE_PHN801_n5758), 
	.A(FE_PHN3138_n5758));
   BUF_X32 FE_PHC793_n4907 (.Z(FE_PHN793_n4907), 
	.A(FE_PHN3136_n4907));
   BUF_X4 FE_PHC783_n152 (.Z(FE_PHN783_n152), 
	.A(n152));
   BUF_X32 FE_PHC780_n2892 (.Z(FE_PHN780_n2892), 
	.A(n2892));
   BUF_X16 FE_PHC779_n5669 (.Z(FE_PHN779_n5669), 
	.A(n5669));
   CLKBUF_X1 FE_PHC778_n160 (.Z(FE_PHN778_n160), 
	.A(n160));
   BUF_X32 FE_PHC776_n1108 (.Z(FE_PHN776_n1108), 
	.A(n1108));
   CLKBUF_X1 FE_PHC775_n5689 (.Z(FE_PHN775_n5689), 
	.A(n5689));
   BUF_X4 FE_PHC774_n14825 (.Z(FE_PHN774_n14825), 
	.A(n14825));
   BUF_X4 FE_PHC770_n140 (.Z(FE_PHN770_n140), 
	.A(n140));
   CLKBUF_X1 FE_PHC769_n5685 (.Z(FE_PHN769_n5685), 
	.A(n5685));
   BUF_X16 FE_PHC768_n72 (.Z(FE_PHN768_n72), 
	.A(n72));
   BUF_X32 FE_PHC765_n1144 (.Z(FE_PHN765_n1144), 
	.A(n1144));
   BUF_X32 FE_PHC763_n1140 (.Z(FE_PHN763_n1140), 
	.A(n1140));
   BUF_X32 FE_PHC762_n4906 (.Z(FE_PHN762_n4906), 
	.A(FE_PHN2945_n4906));
   BUF_X32 FE_PHC760_n5666 (.Z(FE_PHN760_n5666), 
	.A(n5666));
   CLKBUF_X1 FE_PHC756_n1145 (.Z(FE_PHN756_n1145), 
	.A(n1145));
   BUF_X32 FE_PHC755_n1142 (.Z(FE_PHN755_n1142), 
	.A(n1142));
   BUF_X16 FE_PHC753_n5759 (.Z(FE_PHN753_n5759), 
	.A(n5759));
   BUF_X32 FE_PHC752_n1337 (.Z(FE_PHN752_n1337), 
	.A(n1337));
   BUF_X16 FE_PHC749_n5657 (.Z(FE_PHN749_n5657), 
	.A(n5657));
   BUF_X32 FE_PHC748_n2415 (.Z(FE_PHN748_n2415), 
	.A(n2415));
   BUF_X32 FE_PHC743_n3096 (.Z(FE_PHN743_n3096), 
	.A(n3096));
   BUF_X16 FE_PHC741_n5681 (.Z(FE_PHN741_n5681), 
	.A(n5681));
   BUF_X32 FE_PHC739_n5751 (.Z(FE_PHN739_n5751), 
	.A(n5751));
   BUF_X16 FE_PHC738_n5745 (.Z(FE_PHN738_n5745), 
	.A(n5745));
   BUF_X32 FE_PHC737_n5744 (.Z(FE_PHN737_n5744), 
	.A(n5744));
   BUF_X32 FE_PHC735_n100 (.Z(FE_PHN735_n100), 
	.A(n100));
   BUF_X16 FE_PHC733_n5748 (.Z(FE_PHN733_n5748), 
	.A(n5748));
   CLKBUF_X1 FE_PHC732_n5692 (.Z(FE_PHN732_n5692), 
	.A(n5692));
   BUF_X8 FE_PHC731_n5691 (.Z(FE_PHN731_n5691), 
	.A(n5691));
   BUF_X32 FE_PHC730_n5750 (.Z(FE_PHN730_n5750), 
	.A(n5750));
   BUF_X32 FE_PHC729_n5746 (.Z(FE_PHN729_n5746), 
	.A(FE_PHN2936_n5746));
   BUF_X32 FE_PHC728_n2421 (.Z(FE_PHN728_n2421), 
	.A(n2421));
   BUF_X32 FE_PHC727_n3344 (.Z(FE_PHN727_n3344), 
	.A(n3344));
   BUF_X32 FE_PHC723_n5741 (.Z(FE_PHN723_n5741), 
	.A(n5741));
   BUF_X16 FE_PHC722_n5740 (.Z(FE_PHN722_n5740), 
	.A(n5740));
   BUF_X8 FE_PHC721_n5749 (.Z(FE_PHN721_n5749), 
	.A(n5749));
   BUF_X32 FE_PHC720_n5739 (.Z(FE_PHN720_n5739), 
	.A(n5739));
   BUF_X32 FE_PHC719_n190 (.Z(FE_PHN719_n190), 
	.A(n190));
   BUF_X16 FE_PHC717_n5743 (.Z(FE_PHN717_n5743), 
	.A(n5743));
   BUF_X32 FE_PHC716_n5753 (.Z(FE_PHN716_n5753), 
	.A(n5753));
   BUF_X32 FE_PHC715_n5754 (.Z(FE_PHN715_n5754), 
	.A(n5754));
   CLKBUF_X1 FE_PHC712_n5687 (.Z(FE_PHN712_n5687), 
	.A(n5687));
   BUF_X16 FE_PHC711_n28 (.Z(FE_PHN711_n28), 
	.A(n28));
   BUF_X16 FE_PHC707_n5747 (.Z(FE_PHN707_n5747), 
	.A(n5747));
   BUF_X16 FE_PHC705_n5655 (.Z(FE_PHN705_n5655), 
	.A(n5655));
   BUF_X32 FE_PHC704_n5752 (.Z(FE_PHN704_n5752), 
	.A(n5752));
   BUF_X16 FE_PHC703_n44 (.Z(FE_PHN703_n44), 
	.A(n44));
   CLKBUF_X1 FE_PHC702_n171 (.Z(FE_PHN702_n171), 
	.A(n171));
   BUF_X8 FE_PHC701_n5742 (.Z(FE_PHN701_n5742), 
	.A(n5742));
   BUF_X4 FE_PHC693_n166 (.Z(FE_PHN693_n166), 
	.A(FE_PHN3055_n166));
   BUF_X32 FE_PHC685_n2516 (.Z(FE_PHN685_n2516), 
	.A(n2516));
   BUF_X32 FE_PHC679_n2465 (.Z(FE_PHN679_n2465), 
	.A(n2465));
   CLKBUF_X3 FE_PHC675_n17126 (.Z(FE_PHN675_n17126), 
	.A(FE_PHN4624_n17126));
   BUF_X2 FE_PHC674_n17127 (.Z(FE_PHN674_n17127), 
	.A(FE_PHN4629_n17127));
   BUF_X4 FE_OFC667_n17122 (.Z(FE_OFN667_n17122), 
	.A(n17122));
   BUF_X4 FE_OFC666_n17077 (.Z(FE_OFN666_n17077), 
	.A(n17077));
   BUF_X4 FE_OFC665_n17074 (.Z(FE_OFN665_n17074), 
	.A(n17074));
   BUF_X4 FE_OFC663_n17058 (.Z(FE_OFN663_n17058), 
	.A(n17058));
   BUF_X4 FE_OFC661_n17057 (.Z(FE_OFN661_n17057), 
	.A(n17057));
   BUF_X4 FE_OFC659_n17053 (.Z(FE_OFN659_n17053), 
	.A(n17053));
   BUF_X4 FE_OFC656_n17048 (.Z(FE_OFN656_n17048), 
	.A(n17048));
   BUF_X4 FE_OFC654_n17038 (.Z(FE_OFN654_n17038), 
	.A(n17038));
   BUF_X4 FE_OFC652_n17033 (.Z(FE_OFN652_n17033), 
	.A(n17033));
   BUF_X4 FE_OFC651_n17027 (.Z(FE_OFN651_n17027), 
	.A(n17027));
   BUF_X4 FE_OFC648_n17017 (.Z(FE_OFN648_n17017), 
	.A(n17017));
   BUF_X4 FE_OFC646_n16977 (.Z(FE_OFN646_n16977), 
	.A(n16977));
   BUF_X4 FE_OFC645_n16939 (.Z(FE_OFN645_n16939), 
	.A(n16939));
   BUF_X4 FE_OFC644_n16936 (.Z(FE_OFN644_n16936), 
	.A(n16936));
   BUF_X2 FE_OFC643_n16916 (.Z(FE_OFN643_n16916), 
	.A(n16916));
   BUF_X2 FE_OFC642_n16913 (.Z(FE_OFN642_n16913), 
	.A(n16913));
   BUF_X4 FE_OFC641_n16902 (.Z(FE_OFN641_n16902), 
	.A(n16902));
   BUF_X4 FE_OFC639_n16897 (.Z(FE_OFN639_n16897), 
	.A(n16897));
   BUF_X4 FE_OFC638_n16891 (.Z(FE_OFN638_n16891), 
	.A(n16891));
   BUF_X4 FE_OFC636_n16886 (.Z(FE_OFN636_n16886), 
	.A(n16886));
   BUF_X4 FE_OFC635_n16877 (.Z(FE_OFN635_n16877), 
	.A(n16877));
   BUF_X32 FE_OFC634_n16871 (.Z(FE_OFN634_n16871), 
	.A(n16871));
   BUF_X4 FE_OFC633_n16868 (.Z(FE_OFN633_n16868), 
	.A(n16868));
   BUF_X4 FE_OFC632_n16859 (.Z(FE_OFN632_n16859), 
	.A(n16859));
   BUF_X32 FE_OFC631_n16851 (.Z(FE_OFN631_n16851), 
	.A(n16851));
   BUF_X32 FE_OFC629_n16850 (.Z(FE_OFN629_n16850), 
	.A(n16850));
   BUF_X4 FE_OFC628_n16833 (.Z(FE_OFN628_n16833), 
	.A(n16833));
   BUF_X4 FE_OFC627_n16828 (.Z(FE_OFN627_n16828), 
	.A(n16828));
   BUF_X4 FE_OFC626_n16820 (.Z(FE_OFN626_n16820), 
	.A(n16820));
   BUF_X4 FE_OFC625_n16814 (.Z(FE_OFN625_n16814), 
	.A(n16814));
   BUF_X4 FE_OFC610_n16690 (.Z(FE_OFN610_n16690), 
	.A(n16690));
   BUF_X4 FE_OFC608_n16686 (.Z(FE_OFN608_n16686), 
	.A(n16686));
   BUF_X4 FE_OFC602_n16656 (.Z(FE_OFN602_n16656), 
	.A(n16656));
   BUF_X4 FE_OFC598_n5805 (.Z(FE_OFN598_n5805), 
	.A(n5805));
   BUF_X4 FE_OFC587_n5162 (.Z(FE_OFN587_n5162), 
	.A(n5162));
   BUF_X2 FE_OFC583_n5036 (.Z(FE_OFN583_n5036), 
	.A(n5036));
   BUF_X4 FE_OFC573_n4905 (.Z(FE_OFN573_n4905), 
	.A(n4905));
   BUF_X4 FE_OFC568_n4401 (.Z(FE_OFN568_n4401), 
	.A(n4401));
   BUF_X4 FE_OFC567_n4069 (.Z(FE_OFN567_n4069), 
	.A(n4069));
   BUF_X4 FE_OFC566_n4065 (.Z(FE_OFN566_n4065), 
	.A(n4065));
   BUF_X4 FE_OFC565_n4058 (.Z(FE_OFN565_n4058), 
	.A(n4058));
   BUF_X4 FE_OFC560_n3199 (.Z(FE_OFN560_n3199), 
	.A(n3199));
   BUF_X4 FE_OFC559_n3180 (.Z(FE_OFN559_n3180), 
	.A(n3180));
   BUF_X4 FE_OFC549_n2774 (.Z(FE_OFN549_n2774), 
	.A(n2774));
   BUF_X4 FE_OFC544_n2612 (.Z(FE_OFN544_n2612), 
	.A(n2612));
   BUF_X4 FE_OFC543_n2585 (.Z(FE_OFN543_n2585), 
	.A(n2585));
   BUF_X4 FE_OFC542_n2562 (.Z(FE_OFN542_n2562), 
	.A(n2562));
   BUF_X4 FE_OFC541_n2556 (.Z(FE_OFN541_n2556), 
	.A(n2556));
   BUF_X4 FE_OFC539_n2519 (.Z(FE_OFN539_n2519), 
	.A(n2519));
   BUF_X4 FE_OFC538_n2501 (.Z(FE_OFN538_n2501), 
	.A(n2501));
   BUF_X4 FE_OFC537_n2496 (.Z(FE_OFN537_n2496), 
	.A(n2496));
   BUF_X4 FE_OFC534_n2388 (.Z(FE_OFN534_n2388), 
	.A(n2388));
   BUF_X4 FE_OFC533_n2357 (.Z(FE_OFN533_n2357), 
	.A(n2357));
   BUF_X4 FE_OFC530_n2350 (.Z(FE_OFN530_n2350), 
	.A(n2350));
   BUF_X4 FE_OFC529_n2338 (.Z(FE_OFN529_n2338), 
	.A(n2338));
   BUF_X4 FE_OFC527_n2336 (.Z(FE_OFN527_n2336), 
	.A(n2336));
   BUF_X4 FE_OFC525_n2332 (.Z(FE_OFN525_n2332), 
	.A(n2332));
   BUF_X4 FE_OFC523_n2329 (.Z(FE_OFN523_n2329), 
	.A(n2329));
   BUF_X4 FE_OFC519_n2257 (.Z(FE_OFN519_n2257), 
	.A(n2257));
   BUF_X4 FE_OFC516_n2196 (.Z(FE_OFN516_n2196), 
	.A(n2196));
   BUF_X4 FE_OFC514_n2062 (.Z(FE_OFN514_n2062), 
	.A(n2062));
   BUF_X4 FE_OFC512_n2058 (.Z(FE_OFN512_n2058), 
	.A(n2058));
   BUF_X4 FE_OFC511_n2057 (.Z(FE_OFN511_n2057), 
	.A(FE_PSN5239_n2057));
   BUF_X4 FE_OFC510_n2028 (.Z(FE_OFN510_n2028), 
	.A(n2028));
   BUF_X4 FE_OFC509_n2012 (.Z(FE_OFN509_n2012), 
	.A(n2012));
   BUF_X4 FE_OFC506_n1834 (.Z(FE_OFN506_n1834), 
	.A(n1834));
   BUF_X4 FE_OFC504_n1832 (.Z(FE_OFN504_n1832), 
	.A(n1832));
   BUF_X4 FE_OFC495_n1670 (.Z(FE_OFN495_n1670), 
	.A(n1670));
   BUF_X4 FE_OFC493_n1632 (.Z(FE_OFN493_n1632), 
	.A(n1632));
   BUF_X4 FE_OFC490_n1622 (.Z(FE_OFN490_n1622), 
	.A(n1622));
   BUF_X4 FE_OFC486_n1579 (.Z(FE_OFN486_n1579), 
	.A(n1579));
   BUF_X4 FE_OFC485_n1519 (.Z(FE_OFN485_n1519), 
	.A(n1519));
   BUF_X4 FE_OFC484_n1354 (.Z(FE_OFN484_n1354), 
	.A(n1354));
   BUF_X4 FE_OFC483_n1233 (.Z(FE_OFN483_n1233), 
	.A(n1233));
   BUF_X4 FE_OFC479_n1148 (.Z(FE_OFN479_n1148), 
	.A(n1148));
   BUF_X32 FE_OFC469_n1034 (.Z(FE_OFN469_n1034), 
	.A(n1034));
   BUF_X4 FE_OFC466_n998 (.Z(FE_OFN466_n998), 
	.A(n998));
   BUF_X4 FE_OFC465_n945 (.Z(FE_OFN465_n945), 
	.A(n945));
   BUF_X4 FE_OFC461_n890 (.Z(FE_OFN461_n890), 
	.A(n890));
   BUF_X4 FE_OFC458_n860 (.Z(FE_OFN458_n860), 
	.A(n860));
   BUF_X4 FE_OFC456_n822 (.Z(FE_OFN456_n822), 
	.A(n822));
   BUF_X4 FE_OFC450_n808 (.Z(FE_OFN450_n808), 
	.A(n808));
   BUF_X4 FE_OFC429_n673 (.Z(FE_OFN429_n673), 
	.A(n673));
   BUF_X4 FE_OFC426_n659 (.Z(FE_OFN426_n659), 
	.A(n659));
   BUF_X4 FE_OFC425_n650 (.Z(FE_OFN425_n650), 
	.A(n650));
   BUF_X4 FE_OFC422_n641 (.Z(FE_OFN422_n641), 
	.A(n641));
   BUF_X4 FE_OFC419_n628 (.Z(FE_OFN419_n628), 
	.A(n628));
   BUF_X4 FE_OFC414_n556 (.Z(FE_OFN414_n556), 
	.A(n556));
   BUF_X4 FE_OFC411_n499 (.Z(FE_OFN411_n499), 
	.A(n499));
   BUF_X4 FE_OFC384_n118 (.Z(FE_OFN384_n118), 
	.A(n118));
   BUF_X4 FE_OFC383_n71 (.Z(FE_OFN383_n71), 
	.A(n71));
   BUF_X4 FE_OFC382_n64 (.Z(FE_OFN382_n64), 
	.A(n64));
   BUF_X4 FE_OFC208_n2015 (.Z(FE_OFN208_n2015), 
	.A(FE_OFN2_n2015));
   BUF_X4 FE_OFC195_HRESETn (.Z(FE_OFN195_HRESETn), 
	.A(FE_OFN29_HRESETn));
   BUF_X4 FE_OFC194_HRESETn (.Z(FE_OFN194_HRESETn), 
	.A(FE_OFN29_HRESETn));
   BUF_X4 FE_OFC192_HRESETn (.Z(FE_OFN192_HRESETn), 
	.A(FE_OFN30_HRESETn));
   BUF_X4 FE_OFC190_HRESETn (.Z(FE_OFN190_HRESETn), 
	.A(FE_OFN33_HRESETn));
   BUF_X4 FE_OFC185_HRESETn (.Z(FE_OFN185_HRESETn), 
	.A(FE_OFN38_HRESETn));
   BUF_X4 FE_OFC184_HRESETn (.Z(FE_OFN184_HRESETn), 
	.A(FE_OFN38_HRESETn));
   BUF_X4 FE_OFC182_HRESETn (.Z(FE_OFN182_HRESETn), 
	.A(FE_OFN40_HRESETn));
   BUF_X4 FE_OFC181_HRESETn (.Z(FE_OFN181_HRESETn), 
	.A(FE_OFN40_HRESETn));
   BUF_X4 FE_OFC180_HRESETn (.Z(FE_OFN180_HRESETn), 
	.A(FE_OFN41_HRESETn));
   BUF_X4 FE_OFC179_HRESETn (.Z(FE_OFN179_HRESETn), 
	.A(FE_OFN41_HRESETn));
   BUF_X4 FE_OFC178_HRESETn (.Z(FE_OFN178_HRESETn), 
	.A(FE_OFN41_HRESETn));
   BUF_X4 FE_OFC177_HRESETn (.Z(FE_OFN177_HRESETn), 
	.A(FE_OFN41_HRESETn));
   BUF_X4 FE_OFC175_HRESETn (.Z(FE_OFN175_HRESETn), 
	.A(FE_OFN43_HRESETn));
   BUF_X4 FE_OFC174_HRESETn (.Z(FE_OFN174_HRESETn), 
	.A(FE_OFN43_HRESETn));
   BUF_X4 FE_OFC167_HRESETn (.Z(FE_OFN167_HRESETn), 
	.A(FE_OFN48_HRESETn));
   BUF_X4 FE_OFC166_HRESETn (.Z(FE_OFN166_HRESETn), 
	.A(FE_OFN48_HRESETn));
   BUF_X4 FE_OFC165_HRESETn (.Z(FE_OFN165_HRESETn), 
	.A(FE_OFN48_HRESETn));
   BUF_X4 FE_OFC164_HRESETn (.Z(FE_OFN164_HRESETn), 
	.A(FE_OFN49_HRESETn));
   BUF_X4 FE_OFC163_HRESETn (.Z(FE_OFN163_HRESETn), 
	.A(FE_OFN49_HRESETn));
   BUF_X4 FE_OFC159_HRESETn (.Z(FE_OFN159_HRESETn), 
	.A(FE_OFN52_HRESETn));
   BUF_X4 FE_OFC152_HRESETn (.Z(FE_OFN152_HRESETn), 
	.A(FE_OFN56_HRESETn));
   BUF_X4 FE_OFC145_HRESETn (.Z(FE_OFN145_HRESETn), 
	.A(FE_OFN60_HRESETn));
   BUF_X4 FE_OFC144_HRESETn (.Z(FE_OFN144_HRESETn), 
	.A(FE_OFN61_HRESETn));
   BUF_X4 FE_OFC139_HRESETn (.Z(FE_OFN139_HRESETn), 
	.A(FE_OFN65_HRESETn));
   BUF_X4 FE_OFC138_HRESETn (.Z(FE_OFN138_HRESETn), 
	.A(FE_OFN66_HRESETn));
   BUF_X4 FE_OFC135_HRESETn (.Z(FE_OFN135_HRESETn), 
	.A(FE_OFN68_HRESETn));
   INV_X4 FE_OFC132_n2391 (.ZN(FE_OFN132_n2391), 
	.A(FE_OFN131_n2391));
   INV_X4 FE_OFC131_n2391 (.ZN(FE_OFN131_n2391), 
	.A(n2391));
   INV_X4 FE_OFC130_n1750 (.ZN(FE_OFN130_n1750), 
	.A(FE_OFN129_n1750));
   INV_X4 FE_OFC129_n1750 (.ZN(FE_OFN129_n1750), 
	.A(n1750));
   INV_X4 FE_OFC128_n1809 (.ZN(FE_OFN128_n1809), 
	.A(FE_OFN127_n1809));
   INV_X4 FE_OFC127_n1809 (.ZN(FE_OFN127_n1809), 
	.A(n1809));
   INV_X4 FE_OFC126_n2416 (.ZN(FE_OFN126_n2416), 
	.A(FE_OFN125_n2416));
   INV_X4 FE_OFC125_n2416 (.ZN(FE_OFN125_n2416), 
	.A(n2416));
   INV_X4 FE_OFC124_n2079 (.ZN(FE_OFN124_n2079), 
	.A(FE_OFN123_n2079));
   INV_X4 FE_OFC123_n2079 (.ZN(FE_OFN123_n2079), 
	.A(n2079));
   INV_X4 FE_OFC118_HADDR_31_ (.ZN(haddr_o[31]), 
	.A(FE_OFN117_HADDR_31_));
   BUF_X2 FE_OFC117_HADDR_31_ (.Z(FE_OFN118_HADDR_31_), 
	.A(FE_OFN117_HADDR_31_));
   BUF_X2 FE_OFC114_HADDR_29_ (.Z(FE_OFN115_HADDR_29_), 
	.A(FE_OFN113_HADDR_29_));
   INV_X4 FE_OFC113_HADDR_29_ (.ZN(haddr_o[29]), 
	.A(FE_OFN113_HADDR_29_));
   INV_X4 FE_OFC112_HADDR_30_ (.ZN(haddr_o[30]), 
	.A(FE_OFN111_HADDR_30_));
   BUF_X2 FE_OFC111_HADDR_30_ (.Z(FE_OFN112_HADDR_30_), 
	.A(FE_OFN110_HADDR_30_));
   INV_X4 FE_OFC110_HADDR_30_ (.ZN(FE_OFN111_HADDR_30_), 
	.A(FE_OFN110_HADDR_30_));
   INV_X4 FE_OFC109_n16964 (.ZN(FE_OFN109_n16964), 
	.A(FE_OFN108_n16964));
   INV_X1 FE_OFC108_n16964 (.ZN(FE_OFN108_n16964), 
	.A(n16964));
   INV_X4 FE_OFC107_n585 (.ZN(FE_OFN107_n585), 
	.A(FE_OFN105_n585));
   INV_X4 FE_OFC106_n585 (.ZN(FE_OFN106_n585), 
	.A(FE_OFN105_n585));
   INV_X4 FE_OFC105_n585 (.ZN(FE_OFN105_n585), 
	.A(n585));
   INV_X4 FE_OFC104_n715 (.ZN(FE_OFN104_n715), 
	.A(FE_OFN102_n715));
   INV_X4 FE_OFC103_n715 (.ZN(FE_OFN103_n715), 
	.A(FE_OFN102_n715));
   INV_X4 FE_OFC102_n715 (.ZN(FE_OFN102_n715), 
	.A(n715));
   INV_X4 FE_OFC100_n1086 (.ZN(FE_OFN100_n1086), 
	.A(FE_OFN99_n1086));
   INV_X4 FE_OFC99_n1086 (.ZN(FE_OFN99_n1086), 
	.A(n1086));
   BUF_X2 FE_OFC98_n1104 (.Z(FE_OFN98_n1104), 
	.A(n1104));
   INV_X4 FE_OFC95_n16864 (.ZN(FE_OFN95_n16864), 
	.A(FE_OFN93_n16864));
   INV_X4 FE_OFC93_n16864 (.ZN(FE_OFN93_n16864), 
	.A(n16864));
   BUF_X2 FE_OFC91_n16864 (.Z(FE_OFN91_n16864), 
	.A(n16864));
   INV_X4 FE_OFC90_n16849 (.ZN(FE_OFN90_n16849), 
	.A(FE_OFN88_n16849));
   INV_X1 FE_OFC89_n16849 (.ZN(FE_OFN89_n16849), 
	.A(FE_OFN88_n16849));
   INV_X4 FE_OFC88_n16849 (.ZN(FE_OFN88_n16849), 
	.A(n16849));
   INV_X4 FE_OFC87_n16848 (.ZN(FE_OFN87_n16848), 
	.A(FE_OFN86_n16848));
   INV_X4 FE_OFC86_n16848 (.ZN(FE_OFN86_n16848), 
	.A(n16848));
   INV_X4 FE_OFC85_n16839 (.ZN(FE_OFN85_n16839), 
	.A(FE_OFN83_n16839));
   INV_X1 FE_OFC84_n16839 (.ZN(FE_OFN84_n16839), 
	.A(FE_OFN83_n16839));
   INV_X4 FE_OFC83_n16839 (.ZN(FE_OFN83_n16839), 
	.A(n16839));
   INV_X4 FE_OFC82_n16856 (.ZN(FE_OFN82_n16856), 
	.A(FE_OFN80_n16856));
   INV_X4 FE_OFC81_n16856 (.ZN(FE_OFN81_n16856), 
	.A(FE_OFN80_n16856));
   INV_X4 FE_OFC80_n16856 (.ZN(FE_OFN80_n16856), 
	.A(n16856));
   INV_X4 FE_OFC79_n16834 (.ZN(FE_OFN79_n16834), 
	.A(FE_OFN77_n16834));
   INV_X4 FE_OFC78_n16834 (.ZN(FE_OFN78_n16834), 
	.A(FE_OFN77_n16834));
   INV_X4 FE_OFC77_n16834 (.ZN(FE_OFN77_n16834), 
	.A(n16834));
   BUF_X2 FE_OFC75_n16806 (.Z(FE_OFN75_n16806), 
	.A(FE_OFN73_n16806));
   BUF_X4 FE_OFC73_n16806 (.Z(FE_OFN73_n16806), 
	.A(n16806));
   INV_X4 FE_OFC72_n16867 (.ZN(FE_OFN72_n16867), 
	.A(FE_OFN70_n16867));
   INV_X4 FE_OFC70_n16867 (.ZN(FE_OFN70_n16867), 
	.A(n16867));
   BUF_X4 FE_OFC68_HRESETn (.Z(FE_OFN68_HRESETn), 
	.A(FE_OFN163_HRESETn));
   BUF_X4 FE_OFC66_HRESETn (.Z(FE_OFN66_HRESETn), 
	.A(FE_OFN41_HRESETn));
   BUF_X4 FE_OFC65_HRESETn (.Z(FE_OFN65_HRESETn), 
	.A(FE_OFN40_HRESETn));
   BUF_X4 FE_OFC61_HRESETn (.Z(FE_OFN61_HRESETn), 
	.A(FE_OFN38_HRESETn));
   BUF_X4 FE_OFC60_HRESETn (.Z(FE_OFN60_HRESETn), 
	.A(FE_OFN33_HRESETn));
   BUF_X8 FE_OFC56_HRESETn (.Z(FE_OFN56_HRESETn), 
	.A(FE_OFN34_HRESETn));
   BUF_X8 FE_OFC52_HRESETn (.Z(FE_OFN52_HRESETn), 
	.A(FE_OFN192_HRESETn));
   BUF_X8 FE_OFC49_HRESETn (.Z(FE_OFN49_HRESETn), 
	.A(FE_OFN29_HRESETn));
   BUF_X8 FE_OFC48_HRESETn (.Z(FE_OFN48_HRESETn), 
	.A(FE_OFN29_HRESETn));
   INV_X8 FE_OFC41_HRESETn (.ZN(FE_OFN41_HRESETn), 
	.A(hreset_n));
   INV_X8 FE_OFC40_HRESETn (.ZN(FE_OFN40_HRESETn), 
	.A(hreset_n));
   INV_X8 FE_OFC38_HRESETn (.ZN(FE_OFN38_HRESETn), 
	.A(hreset_n));
   INV_X8 FE_OFC33_HRESETn (.ZN(FE_OFN33_HRESETn), 
	.A(hreset_n));
   CLKBUF_X3 FE_OFC21_n503 (.Z(FE_OFN21_n503), 
	.A(n503));
   CLKBUF_X3 FE_OFC19_n1063 (.Z(FE_OFN19_n1063), 
	.A(n1063));
   CLKBUF_X3 FE_OFC17_n16805 (.Z(FE_OFN17_n16805), 
	.A(n16805));
   CLKBUF_X3 FE_OFC15_n16671 (.Z(FE_OFN15_n16671), 
	.A(n16671));
   CLKBUF_X3 FE_OFC10_n1697 (.Z(FE_OFN10_n1697), 
	.A(n1697));
   CLKBUF_X3 FE_OFC2_n2015 (.Z(FE_OFN2_n2015), 
	.A(n2015));
   XNOR2_X2 sub_2068_U1_A_1 (.ZN(sub_2068_SUM_1_), 
	.B(sub_2068_A_0_), 
	.A(sub_2068_A_1_));
   OR2_X1 sub_2068_U1_B_1 (.ZN(sub_2068_carry_2_), 
	.A2(sub_2068_A_0_), 
	.A1(sub_2068_A_1_));
   XNOR2_X2 sub_2068_U1_A_2 (.ZN(sub_2068_SUM_2_), 
	.B(sub_2068_carry_2_), 
	.A(sub_2068_A_2_));
   OR2_X1 sub_2068_U1_B_2 (.ZN(sub_2068_carry_3_), 
	.A2(sub_2068_carry_2_), 
	.A1(sub_2068_A_2_));
   XNOR2_X2 sub_2068_U1_A_3 (.ZN(sub_2068_SUM_3_), 
	.B(sub_2068_carry_3_), 
	.A(sub_2068_A_3_));
   OR2_X1 sub_2068_U1_B_3 (.ZN(sub_2068_carry_4_), 
	.A2(sub_2068_carry_3_), 
	.A1(sub_2068_A_3_));
   XNOR2_X2 sub_2068_U1_A_4 (.ZN(sub_2068_SUM_4_), 
	.B(sub_2068_carry_4_), 
	.A(sub_2068_A_4_));
   OR2_X1 sub_2068_U1_B_4 (.ZN(sub_2068_carry_5_), 
	.A2(sub_2068_carry_4_), 
	.A1(sub_2068_A_4_));
   XNOR2_X2 sub_2068_U1_A_5 (.ZN(sub_2068_SUM_5_), 
	.B(sub_2068_carry_5_), 
	.A(sub_2068_A_5_));
   OR2_X1 sub_2068_U1_B_5 (.ZN(sub_2068_carry_6_), 
	.A2(sub_2068_carry_5_), 
	.A1(sub_2068_A_5_));
   XNOR2_X2 sub_2068_U1_A_6 (.ZN(sub_2068_SUM_6_), 
	.B(sub_2068_carry_6_), 
	.A(sub_2068_A_6_));
   OR2_X1 sub_2068_U1_B_6 (.ZN(sub_2068_carry_7_), 
	.A2(sub_2068_carry_6_), 
	.A1(sub_2068_A_6_));
   XNOR2_X2 sub_2068_U1_A_7 (.ZN(sub_2068_SUM_7_), 
	.B(sub_2068_carry_7_), 
	.A(sub_2068_A_7_));
   OR2_X1 sub_2068_U1_B_7 (.ZN(sub_2068_carry_8_), 
	.A2(sub_2068_carry_7_), 
	.A1(sub_2068_A_7_));
   XNOR2_X2 sub_2068_U1_A_8 (.ZN(sub_2068_SUM_8_), 
	.B(sub_2068_carry_8_), 
	.A(sub_2068_A_8_));
   OR2_X1 sub_2068_U1_B_8 (.ZN(sub_2068_carry_9_), 
	.A2(sub_2068_carry_8_), 
	.A1(sub_2068_A_8_));
   XNOR2_X2 sub_2068_U1_A_9 (.ZN(sub_2068_SUM_9_), 
	.B(sub_2068_carry_9_), 
	.A(sub_2068_A_9_));
   OR2_X1 sub_2068_U1_B_9 (.ZN(sub_2068_carry_10_), 
	.A2(sub_2068_carry_9_), 
	.A1(sub_2068_A_9_));
   XNOR2_X2 sub_2068_U1_A_10 (.ZN(sub_2068_SUM_10_), 
	.B(sub_2068_carry_10_), 
	.A(sub_2068_A_10_));
   OR2_X1 sub_2068_U1_B_10 (.ZN(sub_2068_carry_11_), 
	.A2(sub_2068_carry_10_), 
	.A1(sub_2068_A_10_));
   XNOR2_X2 sub_2068_U1_A_11 (.ZN(sub_2068_SUM_11_), 
	.B(sub_2068_carry_11_), 
	.A(sub_2068_A_11_));
   OR2_X1 sub_2068_U1_B_11 (.ZN(sub_2068_carry_12_), 
	.A2(sub_2068_carry_11_), 
	.A1(sub_2068_A_11_));
   XNOR2_X2 sub_2068_U1_A_12 (.ZN(sub_2068_SUM_12_), 
	.B(sub_2068_carry_12_), 
	.A(sub_2068_A_12_));
   OR2_X1 sub_2068_U1_B_12 (.ZN(sub_2068_carry_13_), 
	.A2(sub_2068_carry_12_), 
	.A1(sub_2068_A_12_));
   XNOR2_X2 sub_2068_U1_A_13 (.ZN(sub_2068_SUM_13_), 
	.B(sub_2068_carry_13_), 
	.A(sub_2068_A_13_));
   OR2_X1 sub_2068_U1_B_13 (.ZN(sub_2068_carry_14_), 
	.A2(sub_2068_carry_13_), 
	.A1(sub_2068_A_13_));
   XNOR2_X2 sub_2068_U1_A_14 (.ZN(sub_2068_SUM_14_), 
	.B(sub_2068_carry_14_), 
	.A(sub_2068_A_14_));
   OR2_X1 sub_2068_U1_B_14 (.ZN(sub_2068_carry_15_), 
	.A2(sub_2068_carry_14_), 
	.A1(sub_2068_A_14_));
   XNOR2_X2 sub_2068_U1_A_15 (.ZN(sub_2068_SUM_15_), 
	.B(sub_2068_carry_15_), 
	.A(sub_2068_A_15_));
   OR2_X1 sub_2068_U1_B_15 (.ZN(sub_2068_carry_16_), 
	.A2(sub_2068_carry_15_), 
	.A1(sub_2068_A_15_));
   XNOR2_X2 sub_2068_U1_A_16 (.ZN(sub_2068_SUM_16_), 
	.B(sub_2068_carry_16_), 
	.A(sub_2068_A_16_));
   OR2_X1 sub_2068_U1_B_16 (.ZN(sub_2068_carry_17_), 
	.A2(sub_2068_carry_16_), 
	.A1(sub_2068_A_16_));
   XNOR2_X2 sub_2068_U1_A_17 (.ZN(sub_2068_SUM_17_), 
	.B(sub_2068_carry_17_), 
	.A(sub_2068_A_17_));
   OR2_X1 sub_2068_U1_B_17 (.ZN(sub_2068_carry_18_), 
	.A2(sub_2068_carry_17_), 
	.A1(sub_2068_A_17_));
   XNOR2_X2 sub_2068_U1_A_18 (.ZN(sub_2068_SUM_18_), 
	.B(sub_2068_carry_18_), 
	.A(sub_2068_A_18_));
   OR2_X1 sub_2068_U1_B_18 (.ZN(sub_2068_carry_19_), 
	.A2(sub_2068_carry_18_), 
	.A1(sub_2068_A_18_));
   XNOR2_X2 sub_2068_U1_A_19 (.ZN(sub_2068_SUM_19_), 
	.B(sub_2068_carry_19_), 
	.A(sub_2068_A_19_));
   OR2_X1 sub_2068_U1_B_19 (.ZN(sub_2068_carry_20_), 
	.A2(sub_2068_carry_19_), 
	.A1(sub_2068_A_19_));
   XNOR2_X2 sub_2068_U1_A_20 (.ZN(sub_2068_SUM_20_), 
	.B(sub_2068_carry_20_), 
	.A(sub_2068_A_20_));
   OR2_X1 sub_2068_U1_B_20 (.ZN(sub_2068_carry_21_), 
	.A2(sub_2068_carry_20_), 
	.A1(sub_2068_A_20_));
   XNOR2_X2 sub_2068_U1_A_21 (.ZN(sub_2068_SUM_21_), 
	.B(sub_2068_carry_21_), 
	.A(sub_2068_A_21_));
   OR2_X1 sub_2068_U1_B_21 (.ZN(sub_2068_carry_22_), 
	.A2(sub_2068_carry_21_), 
	.A1(sub_2068_A_21_));
   XNOR2_X2 sub_2068_U1_A_22 (.ZN(sub_2068_SUM_22_), 
	.B(sub_2068_carry_22_), 
	.A(sub_2068_A_22_));
   OR2_X1 sub_2068_U1_B_22 (.ZN(sub_2068_carry_23_), 
	.A2(sub_2068_carry_22_), 
	.A1(sub_2068_A_22_));
   XNOR2_X2 sub_2069_U1_A_1 (.ZN(sub_2069_SUM_1_), 
	.B(n5829), 
	.A(sub_2069_A_1_));
   OR2_X1 sub_2069_U1_B_1 (.ZN(sub_2069_carry_2_), 
	.A2(n5829), 
	.A1(sub_2069_A_1_));
   XNOR2_X2 sub_2069_U1_A_2 (.ZN(sub_2069_SUM_2_), 
	.B(sub_2069_carry_2_), 
	.A(sub_2069_A_2_));
   OR2_X1 sub_2069_U1_B_2 (.ZN(sub_2069_carry_3_), 
	.A2(sub_2069_carry_2_), 
	.A1(sub_2069_A_2_));
   XNOR2_X2 sub_2069_U1_A_3 (.ZN(sub_2069_SUM_3_), 
	.B(sub_2069_carry_3_), 
	.A(sub_2069_A_3_));
   OR2_X1 sub_2069_U1_B_3 (.ZN(sub_2069_carry_4_), 
	.A2(sub_2069_carry_3_), 
	.A1(sub_2069_A_3_));
   XNOR2_X2 sub_2069_U1_A_4 (.ZN(sub_2069_SUM_4_), 
	.B(sub_2069_carry_4_), 
	.A(sub_2069_A_4_));
   OR2_X1 sub_2069_U1_B_4 (.ZN(sub_2069_carry_5_), 
	.A2(sub_2069_carry_4_), 
	.A1(sub_2069_A_4_));
   XNOR2_X2 sub_2069_U1_A_5 (.ZN(sub_2069_SUM_5_), 
	.B(sub_2069_carry_5_), 
	.A(sub_2069_A_5_));
   OR2_X1 sub_2069_U1_B_5 (.ZN(sub_2069_carry_6_), 
	.A2(sub_2069_carry_5_), 
	.A1(sub_2069_A_5_));
   XNOR2_X2 sub_2069_U1_A_6 (.ZN(sub_2069_SUM_6_), 
	.B(sub_2069_carry_6_), 
	.A(sub_2069_A_6_));
   OR2_X1 sub_2069_U1_B_6 (.ZN(sub_2069_carry_7_), 
	.A2(sub_2069_carry_6_), 
	.A1(sub_2069_A_6_));
   XNOR2_X2 sub_2069_U1_A_7 (.ZN(sub_2069_SUM_7_), 
	.B(sub_2069_carry_7_), 
	.A(sub_2069_A_7_));
   OR2_X1 sub_2069_U1_B_7 (.ZN(sub_2069_carry_8_), 
	.A2(sub_2069_carry_7_), 
	.A1(sub_2069_A_7_));
   XNOR2_X2 sub_2069_U1_A_8 (.ZN(sub_2069_SUM_8_), 
	.B(sub_2069_carry_8_), 
	.A(sub_2069_A_8_));
   HA_X1 add_2071_U1_1_1 (.S(add_2071_SUM_1_), 
	.CO(add_2071_carry[2]), 
	.B(vis_pc_o[0]), 
	.A(vis_pc_o[1]));
   HA_X1 add_2071_U1_1_2 (.S(add_2071_SUM_2_), 
	.CO(add_2071_carry[3]), 
	.B(add_2071_carry[2]), 
	.A(vis_pc_o[2]));
   HA_X1 add_2071_U1_1_3 (.S(add_2071_SUM_3_), 
	.CO(add_2071_carry[4]), 
	.B(add_2071_carry[3]), 
	.A(vis_pc_o[3]));
   HA_X1 add_2071_U1_1_4 (.S(add_2071_SUM_4_), 
	.CO(add_2071_carry[5]), 
	.B(add_2071_carry[4]), 
	.A(vis_pc_o[4]));
   HA_X1 add_2071_U1_1_5 (.S(add_2071_SUM_5_), 
	.CO(add_2071_carry[6]), 
	.B(add_2071_carry[5]), 
	.A(FE_PHN1339_SYNOPSYS_UNCONNECTED_540));
   HA_X1 add_2071_U1_1_6 (.S(add_2071_SUM_6_), 
	.CO(add_2071_carry[7]), 
	.B(add_2071_carry[6]), 
	.A(vis_pc_o[6]));
   HA_X1 add_2071_U1_1_7 (.S(add_2071_SUM_7_), 
	.CO(add_2071_carry[8]), 
	.B(add_2071_carry[7]), 
	.A(vis_pc_o[7]));
   HA_X1 add_2071_U1_1_8 (.S(add_2071_SUM_8_), 
	.CO(add_2071_carry[9]), 
	.B(add_2071_carry[8]), 
	.A(vis_pc_o[8]));
   HA_X1 add_2071_U1_1_9 (.S(add_2071_SUM_9_), 
	.CO(add_2071_carry[10]), 
	.B(add_2071_carry[9]), 
	.A(vis_pc_o[9]));
   HA_X1 add_2071_U1_1_10 (.S(add_2071_SUM_10_), 
	.CO(add_2071_carry[11]), 
	.B(add_2071_carry[10]), 
	.A(vis_pc_o[10]));
   HA_X1 add_2071_U1_1_11 (.S(add_2071_SUM_11_), 
	.CO(add_2071_carry[12]), 
	.B(add_2071_carry[11]), 
	.A(vis_pc_o[11]));
   HA_X1 add_2071_U1_1_12 (.S(add_2071_SUM_12_), 
	.CO(add_2071_carry[13]), 
	.B(add_2071_carry[12]), 
	.A(vis_pc_o[12]));
   HA_X1 add_2071_U1_1_13 (.S(add_2071_SUM_13_), 
	.CO(add_2071_carry[14]), 
	.B(add_2071_carry[13]), 
	.A(vis_pc_o[13]));
   HA_X1 add_2071_U1_1_14 (.S(add_2071_SUM_14_), 
	.CO(add_2071_carry[15]), 
	.B(add_2071_carry[14]), 
	.A(FE_PHN1341_SYNOPSYS_UNCONNECTED_531));
   HA_X1 add_2071_U1_1_15 (.S(add_2071_SUM_15_), 
	.CO(add_2071_carry[16]), 
	.B(add_2071_carry[15]), 
	.A(vis_pc_o[15]));
   HA_X1 add_2071_U1_1_16 (.S(add_2071_SUM_16_), 
	.CO(add_2071_carry[17]), 
	.B(add_2071_carry[16]), 
	.A(vis_pc_o[16]));
   HA_X1 add_2071_U1_1_17 (.S(add_2071_SUM_17_), 
	.CO(add_2071_carry[18]), 
	.B(add_2071_carry[17]), 
	.A(vis_pc_o[17]));
   HA_X1 add_2071_U1_1_18 (.S(add_2071_SUM_18_), 
	.CO(add_2071_carry[19]), 
	.B(add_2071_carry[18]), 
	.A(vis_pc_o[18]));
   HA_X1 add_2071_U1_1_19 (.S(add_2071_SUM_19_), 
	.CO(add_2071_carry[20]), 
	.B(add_2071_carry[19]), 
	.A(vis_pc_o[19]));
   HA_X1 add_2071_U1_1_20 (.S(add_2071_SUM_20_), 
	.CO(add_2071_carry[21]), 
	.B(add_2071_carry[20]), 
	.A(vis_pc_o[20]));
   HA_X1 add_2071_U1_1_21 (.S(add_2071_SUM_21_), 
	.CO(add_2071_carry[22]), 
	.B(add_2071_carry[21]), 
	.A(vis_pc_o[21]));
   HA_X1 add_2071_U1_1_22 (.S(add_2071_SUM_22_), 
	.CO(add_2071_carry[23]), 
	.B(add_2071_carry[22]), 
	.A(vis_pc_o[22]));
   HA_X1 add_2071_U1_1_23 (.S(add_2071_SUM_23_), 
	.CO(add_2071_carry[24]), 
	.B(add_2071_carry[23]), 
	.A(FE_PHN1331_SYNOPSYS_UNCONNECTED_522));
   HA_X1 add_2071_U1_1_24 (.S(add_2071_SUM_24_), 
	.CO(add_2071_carry[25]), 
	.B(add_2071_carry[24]), 
	.A(vis_pc_o[24]));
   HA_X1 add_2071_U1_1_25 (.S(add_2071_SUM_25_), 
	.CO(add_2071_carry[26]), 
	.B(add_2071_carry[25]), 
	.A(vis_pc_o[25]));
   HA_X1 add_2071_U1_1_26 (.S(add_2071_SUM_26_), 
	.CO(add_2071_carry[27]), 
	.B(add_2071_carry[26]), 
	.A(vis_pc_o[26]));
   HA_X1 add_2071_U1_1_27 (.S(add_2071_SUM_27_), 
	.CO(add_2071_carry[28]), 
	.B(add_2071_carry[27]), 
	.A(FE_PHN1320_SYNOPSYS_UNCONNECTED_518));
   HA_X1 add_2071_U1_1_28 (.S(add_2071_SUM_28_), 
	.CO(add_2071_carry[29]), 
	.B(add_2071_carry[28]), 
	.A(vis_pc_o[28]));
   HA_X1 add_2071_U1_1_29 (.S(add_2071_SUM_29_), 
	.CO(add_2071_carry[30]), 
	.B(add_2071_carry[29]), 
	.A(vis_pc_o[29]));
   HA_X1 add_2072_U1_1_1 (.S(add_2072_SUM_1_), 
	.CO(add_2072_carry[2]), 
	.B(n5797), 
	.A(vis_pc_o[2]));
   HA_X1 add_2072_U1_1_2 (.S(add_2072_SUM_2_), 
	.CO(add_2072_carry[3]), 
	.B(add_2072_carry[2]), 
	.A(vis_pc_o[3]));
   HA_X1 add_2072_U1_1_3 (.S(add_2072_SUM_3_), 
	.CO(add_2072_carry[4]), 
	.B(add_2072_carry[3]), 
	.A(vis_pc_o[4]));
   HA_X1 add_2072_U1_1_4 (.S(add_2072_SUM_4_), 
	.CO(add_2072_carry[5]), 
	.B(add_2072_carry[4]), 
	.A(FE_PHN1339_SYNOPSYS_UNCONNECTED_540));
   HA_X1 add_2072_U1_1_5 (.S(add_2072_SUM_5_), 
	.CO(add_2072_carry[6]), 
	.B(add_2072_carry[5]), 
	.A(vis_pc_o[6]));
   HA_X1 add_2072_U1_1_6 (.S(add_2072_SUM_6_), 
	.CO(add_2072_carry[7]), 
	.B(add_2072_carry[6]), 
	.A(vis_pc_o[7]));
   HA_X1 add_2072_U1_1_7 (.S(add_2072_SUM_7_), 
	.CO(add_2072_carry[8]), 
	.B(add_2072_carry[7]), 
	.A(vis_pc_o[8]));
   HA_X1 add_2072_U1_1_8 (.S(add_2072_SUM_8_), 
	.CO(add_2072_carry[9]), 
	.B(add_2072_carry[8]), 
	.A(vis_pc_o[9]));
   HA_X1 add_2072_U1_1_9 (.S(add_2072_SUM_9_), 
	.CO(add_2072_carry[10]), 
	.B(add_2072_carry[9]), 
	.A(vis_pc_o[10]));
   HA_X1 add_2072_U1_1_10 (.S(add_2072_SUM_10_), 
	.CO(add_2072_carry[11]), 
	.B(add_2072_carry[10]), 
	.A(vis_pc_o[11]));
   HA_X1 add_2072_U1_1_11 (.S(add_2072_SUM_11_), 
	.CO(add_2072_carry[12]), 
	.B(add_2072_carry[11]), 
	.A(vis_pc_o[12]));
   HA_X1 add_2072_U1_1_12 (.S(add_2072_SUM_12_), 
	.CO(add_2072_carry[13]), 
	.B(add_2072_carry[12]), 
	.A(vis_pc_o[13]));
   HA_X1 add_2072_U1_1_13 (.S(add_2072_SUM_13_), 
	.CO(add_2072_carry[14]), 
	.B(add_2072_carry[13]), 
	.A(FE_PHN1341_SYNOPSYS_UNCONNECTED_531));
   HA_X1 add_2072_U1_1_14 (.S(add_2072_SUM_14_), 
	.CO(add_2072_carry[15]), 
	.B(add_2072_carry[14]), 
	.A(vis_pc_o[15]));
   HA_X1 add_2072_U1_1_15 (.S(add_2072_SUM_15_), 
	.CO(add_2072_carry[16]), 
	.B(add_2072_carry[15]), 
	.A(vis_pc_o[16]));
   HA_X1 add_2072_U1_1_16 (.S(add_2072_SUM_16_), 
	.CO(add_2072_carry[17]), 
	.B(add_2072_carry[16]), 
	.A(vis_pc_o[17]));
   HA_X1 add_2072_U1_1_17 (.S(add_2072_SUM_17_), 
	.CO(add_2072_carry[18]), 
	.B(add_2072_carry[17]), 
	.A(vis_pc_o[18]));
   HA_X1 add_2072_U1_1_18 (.S(add_2072_SUM_18_), 
	.CO(add_2072_carry[19]), 
	.B(add_2072_carry[18]), 
	.A(vis_pc_o[19]));
   HA_X1 add_2072_U1_1_19 (.S(add_2072_SUM_19_), 
	.CO(add_2072_carry[20]), 
	.B(add_2072_carry[19]), 
	.A(vis_pc_o[20]));
   HA_X1 add_2072_U1_1_20 (.S(add_2072_SUM_20_), 
	.CO(add_2072_carry[21]), 
	.B(add_2072_carry[20]), 
	.A(vis_pc_o[21]));
   HA_X1 add_2072_U1_1_21 (.S(add_2072_SUM_21_), 
	.CO(add_2072_carry[22]), 
	.B(add_2072_carry[21]), 
	.A(vis_pc_o[22]));
   HA_X1 add_2072_U1_1_22 (.S(add_2072_SUM_22_), 
	.CO(add_2072_carry[23]), 
	.B(add_2072_carry[22]), 
	.A(vis_pc_o[23]));
   HA_X1 add_2072_U1_1_23 (.S(add_2072_SUM_23_), 
	.CO(add_2072_carry[24]), 
	.B(add_2072_carry[23]), 
	.A(vis_pc_o[24]));
   HA_X1 add_2072_U1_1_24 (.S(add_2072_SUM_24_), 
	.CO(add_2072_carry[25]), 
	.B(add_2072_carry[24]), 
	.A(vis_pc_o[25]));
   HA_X1 add_2072_U1_1_25 (.S(add_2072_SUM_25_), 
	.CO(add_2072_carry[26]), 
	.B(add_2072_carry[25]), 
	.A(vis_pc_o[26]));
   HA_X1 add_2072_U1_1_26 (.S(add_2072_SUM_26_), 
	.CO(add_2072_carry[27]), 
	.B(add_2072_carry[26]), 
	.A(FE_PHN1320_SYNOPSYS_UNCONNECTED_518));
   HA_X1 add_2072_U1_1_27 (.S(add_2072_SUM_27_), 
	.CO(add_2072_carry[28]), 
	.B(add_2072_carry[27]), 
	.A(vis_pc_o[28]));
   HA_X1 add_2072_U1_1_28 (.S(add_2072_SUM_28_), 
	.CO(add_2072_carry[29]), 
	.B(add_2072_carry[28]), 
	.A(vis_pc_o[29]));
   FA_X1 add_2082_U1_2 (.S(add_2073_A_2_), 
	.CO(add_2082_carry[3]), 
	.CI(n16691), 
	.B(n5822), 
	.A(add_2082_A_2_));
   FA_X1 add_2082_U1_3 (.S(add_2073_A_3_), 
	.CO(add_2082_carry[4]), 
	.CI(add_2082_carry[3]), 
	.B(n5806), 
	.A(add_2082_A_3_));
   FA_X1 add_2082_U1_4 (.S(add_2073_A_4_), 
	.CO(add_2082_carry[5]), 
	.CI(add_2082_carry[4]), 
	.B(add_2082_B_4_), 
	.A(add_2082_A_4_));
   FA_X1 add_2082_U1_5 (.S(add_2073_A_5_), 
	.CO(add_2082_carry[6]), 
	.CI(add_2082_carry[5]), 
	.B(n5801), 
	.A(add_2082_A_5_));
   FA_X1 add_2082_U1_6 (.S(add_2073_A_6_), 
	.CO(add_2082_carry[7]), 
	.CI(add_2082_carry[6]), 
	.B(n5802), 
	.A(add_2082_A_6_));
   FA_X1 add_2082_U1_7 (.S(add_2073_A_7_), 
	.CO(add_2082_carry[8]), 
	.CI(add_2082_carry[7]), 
	.B(n5817), 
	.A(add_2082_A_7_));
   FA_X1 add_2082_U1_8 (.S(add_2073_A_8_), 
	.CO(add_2082_carry[9]), 
	.CI(add_2082_carry[8]), 
	.B(n5821), 
	.A(add_2082_A_8_));
   FA_X1 add_2082_U1_9 (.S(add_2073_A_9_), 
	.CO(add_2082_carry[10]), 
	.CI(add_2082_carry[9]), 
	.B(n5819), 
	.A(add_2082_A_9_));
   FA_X1 add_2082_U1_10 (.S(add_2073_A_10_), 
	.CO(add_2082_carry[11]), 
	.CI(add_2082_carry[10]), 
	.B(n5805), 
	.A(add_2082_A_10_));
   FA_X1 add_2082_U1_11 (.S(add_2073_A_11_), 
	.CO(add_2082_carry[12]), 
	.CI(add_2082_carry[11]), 
	.B(n5804), 
	.A(add_2082_A_11_));
   FA_X1 add_2082_U1_12 (.S(add_2073_A_12_), 
	.CO(add_2082_carry[13]), 
	.CI(add_2082_carry[12]), 
	.B(n5820), 
	.A(add_2082_A_12_));
   FA_X1 add_2082_U1_13 (.S(add_2073_A_13_), 
	.CO(add_2082_carry[14]), 
	.CI(add_2082_carry[13]), 
	.B(n5807), 
	.A(add_2082_A_13_));
   FA_X1 add_2082_U1_14 (.S(add_2073_A_14_), 
	.CO(add_2082_carry[15]), 
	.CI(add_2082_carry[14]), 
	.B(n5808), 
	.A(add_2082_A_14_));
   FA_X1 add_2082_U1_15 (.S(add_2073_A_15_), 
	.CO(add_2082_carry[16]), 
	.CI(add_2082_carry[15]), 
	.B(n5809), 
	.A(add_2082_A_15_));
   FA_X1 add_2082_U1_16 (.S(add_2073_A_16_), 
	.CO(add_2082_carry[17]), 
	.CI(add_2082_carry[16]), 
	.B(n5818), 
	.A(add_2082_A_16_));
   FA_X1 add_2082_U1_17 (.S(add_2073_A_17_), 
	.CO(add_2082_carry[18]), 
	.CI(add_2082_carry[17]), 
	.B(n5810), 
	.A(add_2082_A_17_));
   FA_X1 add_2082_U1_18 (.S(add_2073_A_18_), 
	.CO(add_2082_carry[19]), 
	.CI(add_2082_carry[18]), 
	.B(n5811), 
	.A(add_2082_A_18_));
   FA_X1 add_2082_U1_19 (.S(add_2073_A_19_), 
	.CO(add_2082_carry[20]), 
	.CI(add_2082_carry[19]), 
	.B(n5812), 
	.A(add_2082_A_19_));
   FA_X1 add_2082_U1_20 (.S(add_2073_A_20_), 
	.CO(add_2082_carry[21]), 
	.CI(add_2082_carry[20]), 
	.B(n5813), 
	.A(add_2082_A_20_));
   FA_X1 add_2082_U1_21 (.S(add_2073_A_21_), 
	.CO(add_2082_carry[22]), 
	.CI(add_2082_carry[21]), 
	.B(n5814), 
	.A(add_2082_A_21_));
   FA_X1 add_2082_U1_22 (.S(add_2073_A_22_), 
	.CO(add_2082_carry[23]), 
	.CI(add_2082_carry[22]), 
	.B(n5815), 
	.A(add_2082_A_22_));
   FA_X1 add_2082_U1_23 (.S(add_2073_A_23_), 
	.CO(add_2082_carry[24]), 
	.CI(add_2082_carry[23]), 
	.B(n5816), 
	.A(add_2082_A_23_));
   FA_X1 add_2082_U1_24 (.S(add_2073_A_24_), 
	.CO(add_2082_carry[25]), 
	.CI(add_2082_carry[24]), 
	.B(n5803), 
	.A(add_2082_A_24_));
   FA_X1 add_2082_U1_25 (.S(add_2073_A_25_), 
	.CO(add_2082_carry[26]), 
	.CI(add_2082_carry[25]), 
	.B(U163_Z_0), 
	.A(add_2082_A_25_));
   FA_X1 add_2082_U1_26 (.S(add_2073_A_26_), 
	.CO(add_2082_carry[27]), 
	.CI(add_2082_carry[26]), 
	.B(n4951), 
	.A(add_2082_A_26_));
   FA_X1 add_2082_U1_27 (.S(add_2073_A_27_), 
	.CO(add_2082_carry[28]), 
	.CI(add_2082_carry[27]), 
	.B(n4952), 
	.A(add_2082_A_27_));
   FA_X1 add_2082_U1_28 (.S(add_2073_A_28_), 
	.CO(add_2082_carry[29]), 
	.CI(add_2082_carry[28]), 
	.B(U175_Z_0), 
	.A(add_2082_A_28_));
   FA_X1 add_2082_U1_29 (.S(add_2073_A_29_), 
	.CO(add_2082_carry[30]), 
	.CI(add_2082_carry[29]), 
	.B(U189_Z_0), 
	.A(add_2082_A_29_));
   FA_X1 add_2082_U1_30 (.S(add_2073_A_30_), 
	.CO(add_2082_carry[31]), 
	.CI(add_2082_carry[30]), 
	.B(U158_Z_0), 
	.A(add_2082_A_30_));
   FA_X1 add_2082_U1_31 (.S(add_2073_A_31_), 
	.CO(add_2082_carry[32]), 
	.CI(add_2082_carry[31]), 
	.B(U180_Z_0), 
	.A(add_2082_A_31_));
   FA_X1 add_2082_U1_32 (.S(add_2073_A_32_), 
	.CO(add_2082_carry[33]), 
	.CI(add_2082_carry[32]), 
	.B(U186_Z_0), 
	.A(n4949));
   NOR2_X1 U3 (.ZN(sub_2069_A_8_), 
	.A2(n2), 
	.A1(n5034));
   NOR2_X1 U4 (.ZN(sub_2069_A_7_), 
	.A2(n3), 
	.A1(n5034));
   NOR2_X1 U5 (.ZN(sub_2069_A_6_), 
	.A2(n4), 
	.A1(n5034));
   NOR2_X1 U6 (.ZN(sub_2069_A_5_), 
	.A2(n5), 
	.A1(n5034));
   NOR2_X1 U8 (.ZN(sub_2069_A_4_), 
	.A2(n6), 
	.A1(n5034));
   NOR2_X1 U9 (.ZN(sub_2069_A_3_), 
	.A2(n7), 
	.A1(n5034));
   NOR2_X1 U10 (.ZN(sub_2069_A_2_), 
	.A2(n8), 
	.A1(n5034));
   NOR2_X1 U11 (.ZN(sub_2069_A_1_), 
	.A2(n9), 
	.A1(n5034));
   OAI21_X1 U13 (.ZN(n5654), 
	.B2(n12), 
	.B1(n11), 
	.A(FE_PHN3615_n4746));
   NAND4_X1 U14 (.ZN(n12), 
	.A4(n15), 
	.A3(hwdata_o[2]), 
	.A2(n14), 
	.A1(n13));
   NOR4_X1 U15 (.ZN(n15), 
	.A4(n19), 
	.A3(n18), 
	.A2(n17), 
	.A1(n16));
   INV_X1 U16 (.ZN(n16), 
	.A(n20));
   NAND4_X1 U17 (.ZN(n11), 
	.A4(n23), 
	.A3(n22), 
	.A2(hwdata_o[17]), 
	.A1(n21));
   NOR4_X1 U18 (.ZN(n23), 
	.A4(n25), 
	.A3(n24), 
	.A2(hwdata_o[30]), 
	.A1(hwdata_o[29]));
   OAI221_X1 U19 (.ZN(n5655), 
	.C2(n29), 
	.C1(FE_PHN711_n28), 
	.B2(n27), 
	.B1(n16644), 
	.A(n30));
   AOI221_X1 U20 (.ZN(n30), 
	.C2(n5006), 
	.C1(n33), 
	.B2(vis_pc_o[30]), 
	.B1(n31), 
	.A(n17120));
   AND2_X1 U21 (.ZN(n33), 
	.A2(add_2071_carry[30]), 
	.A1(n17117));
   OAI21_X1 U22 (.ZN(n31), 
	.B2(n36), 
	.B1(add_2071_carry[30]), 
	.A(n37));
   OAI211_X1 U24 (.ZN(n5656), 
	.C2(n29), 
	.C1(n39), 
	.B(n41), 
	.A(n40));
   AOI22_X1 U25 (.ZN(n41), 
	.B2(vis_pc_o[6]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_6_));
   AOI21_X1 U27 (.ZN(n40), 
	.B2(n17116), 
	.B1(n16726), 
	.A(n17120));
   OAI211_X1 U28 (.ZN(n5657), 
	.C2(n29), 
	.C1(FE_PHN703_n44), 
	.B(n46), 
	.A(n45));
   AOI22_X1 U29 (.ZN(n46), 
	.B2(vis_pc_o[22]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_22_));
   AOI21_X1 U31 (.ZN(n45), 
	.B2(n17116), 
	.B1(n16705), 
	.A(n17120));
   OAI211_X1 U32 (.ZN(n5658), 
	.C2(n29), 
	.C1(n48), 
	.B(n50), 
	.A(n49));
   AOI22_X1 U33 (.ZN(n50), 
	.B2(FE_PHN1341_SYNOPSYS_UNCONNECTED_531), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_14_));
   AOI21_X1 U34 (.ZN(n49), 
	.B2(n17116), 
	.B1(n16715), 
	.A(n17120));
   OAI211_X1 U35 (.ZN(n5659), 
	.C2(n37), 
	.C1(FE_PHN3099_n5601), 
	.B(n53), 
	.A(n52));
   AOI222_X1 U36 (.ZN(n53), 
	.C2(n55), 
	.C1(n54), 
	.B2(n17116), 
	.B1(n16706), 
	.A2(n17117), 
	.A1(add_2071_SUM_19_));
   OAI211_X1 U37 (.ZN(n5660), 
	.C2(n37), 
	.C1(FE_PHN3100_n5573), 
	.B(n56), 
	.A(n52));
   AOI222_X1 U38 (.ZN(n56), 
	.C2(n57), 
	.C1(n54), 
	.B2(n17116), 
	.B1(n16668), 
	.A2(n17117), 
	.A1(add_2071_SUM_20_));
   INV_X1 U39 (.ZN(n57), 
	.A(n58));
   OAI211_X1 U40 (.ZN(n5661), 
	.C2(n37), 
	.C1(FE_PHN3098_n5238), 
	.B(n59), 
	.A(n52));
   AOI222_X1 U41 (.ZN(n59), 
	.C2(n60), 
	.C1(n54), 
	.B2(n17116), 
	.B1(n16702), 
	.A2(n17117), 
	.A1(add_2071_SUM_21_));
   INV_X1 U42 (.ZN(n60), 
	.A(n61));
   OAI211_X1 U43 (.ZN(n5662), 
	.C2(n37), 
	.C1(FE_PHN3102_n5237), 
	.B(n62), 
	.A(n52));
   AOI222_X1 U44 (.ZN(n62), 
	.C2(n63), 
	.C1(n54), 
	.B2(n17116), 
	.B1(n16672), 
	.A2(n17117), 
	.A1(add_2071_SUM_17_));
   INV_X1 U45 (.ZN(n63), 
	.A(n64));
   OAI211_X1 U46 (.ZN(n5663), 
	.C2(n37), 
	.C1(FE_PHN3097_n5236), 
	.B(n65), 
	.A(n52));
   AOI222_X1 U47 (.ZN(n65), 
	.C2(n66), 
	.C1(n54), 
	.B2(n17116), 
	.B1(n16710), 
	.A2(n17117), 
	.A1(add_2071_SUM_16_));
   OAI211_X1 U48 (.ZN(n5664), 
	.C2(n37), 
	.C1(FE_PHN3101_n5235), 
	.B(n67), 
	.A(n52));
   AOI222_X1 U49 (.ZN(n67), 
	.C2(n68), 
	.C1(n54), 
	.B2(n17116), 
	.B1(n16711), 
	.A2(n17117), 
	.A1(add_2071_SUM_15_));
   OAI211_X1 U50 (.ZN(n5665), 
	.C2(n37), 
	.C1(FE_PHN1717_n5114), 
	.B(n69), 
	.A(n52));
   AOI222_X1 U51 (.ZN(n69), 
	.C2(n70), 
	.C1(n54), 
	.B2(n17116), 
	.B1(n16709), 
	.A2(n17117), 
	.A1(add_2071_SUM_18_));
   AOI21_X1 U52 (.ZN(n52), 
	.B2(FE_OFN383_n71), 
	.B1(n54), 
	.A(n17120));
   OAI211_X1 U53 (.ZN(n5666), 
	.C2(n29), 
	.C1(FE_PHN768_n72), 
	.B(n74), 
	.A(n73));
   AOI22_X1 U54 (.ZN(n74), 
	.B2(vis_pc_o[28]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_28_));
   AOI21_X1 U55 (.ZN(n73), 
	.B2(n17116), 
	.B1(n16693), 
	.A(n17120));
   OAI211_X1 U56 (.ZN(n5667), 
	.C2(n29), 
	.C1(n76), 
	.B(n78), 
	.A(n77));
   AOI22_X1 U57 (.ZN(n78), 
	.B2(FE_PHN1320_SYNOPSYS_UNCONNECTED_518), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_27_));
   AOI21_X1 U58 (.ZN(n77), 
	.B2(n17116), 
	.B1(n16695), 
	.A(n17120));
   OAI22_X1 U59 (.ZN(n5668), 
	.B2(n83), 
	.B1(n82), 
	.A2(FE_PHN675_n17126), 
	.A1(n80));
   AOI21_X1 U61 (.ZN(n82), 
	.B2(n85), 
	.B1(n84), 
	.A(FE_PHN674_n17127));
   AOI221_X1 U62 (.ZN(n80), 
	.C2(n89), 
	.C1(n88), 
	.B2(n87), 
	.B1(n86), 
	.A(n90));
   AND3_X1 U63 (.ZN(n90), 
	.A3(n84), 
	.A2(n92), 
	.A1(n91));
   OAI33_X1 U64 (.ZN(n91), 
	.B3(n94), 
	.B2(n16688), 
	.B1(n93), 
	.A3(n4949), 
	.A2(U186_Z_0), 
	.A1(n27));
   INV_X1 U65 (.ZN(n87), 
	.A(n76));
   OAI211_X1 U66 (.ZN(n5669), 
	.C2(n29), 
	.C1(n95), 
	.B(n97), 
	.A(n96));
   AOI22_X1 U67 (.ZN(n97), 
	.B2(vis_pc_o[26]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_26_));
   AOI21_X1 U69 (.ZN(n96), 
	.B2(n17116), 
	.B1(n16698), 
	.A(n17120));
   INV_X1 U70 (.ZN(n95), 
	.A(n99));
   OAI211_X1 U71 (.ZN(n5670), 
	.C2(n29), 
	.C1(FE_PHN735_n100), 
	.B(n102), 
	.A(n101));
   AOI22_X1 U72 (.ZN(n102), 
	.B2(vis_pc_o[25]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_25_));
   AOI21_X1 U74 (.ZN(n101), 
	.B2(n17116), 
	.B1(n16663), 
	.A(n17120));
   OAI211_X1 U75 (.ZN(n5671), 
	.C2(n29), 
	.C1(n104), 
	.B(n106), 
	.A(n105));
   AOI22_X1 U76 (.ZN(n106), 
	.B2(vis_pc_o[24]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_24_));
   AOI21_X1 U78 (.ZN(n105), 
	.B2(n17116), 
	.B1(n16655), 
	.A(n17120));
   INV_X1 U79 (.ZN(n104), 
	.A(n108));
   OAI211_X1 U80 (.ZN(n5672), 
	.C2(n29), 
	.C1(n109), 
	.B(n111), 
	.A(n110));
   AOI22_X1 U81 (.ZN(n111), 
	.B2(FE_PHN1331_SYNOPSYS_UNCONNECTED_522), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_23_));
   AOI21_X1 U82 (.ZN(n110), 
	.B2(n17116), 
	.B1(n16701), 
	.A(n17120));
   OAI211_X1 U83 (.ZN(n5673), 
	.C2(n29), 
	.C1(n113), 
	.B(n115), 
	.A(n114));
   AOI22_X1 U84 (.ZN(n115), 
	.B2(vis_pc_o[29]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_29_));
   AOI21_X1 U86 (.ZN(n114), 
	.B2(n17116), 
	.B1(add_2073_SUM_31_), 
	.A(n17120));
   INV_X1 U87 (.ZN(n113), 
	.A(n117));
   OAI211_X1 U88 (.ZN(n5674), 
	.C2(n29), 
	.C1(FE_OFN384_n118), 
	.B(n120), 
	.A(n119));
   AOI22_X1 U89 (.ZN(n120), 
	.B2(vis_pc_o[12]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_12_));
   AOI21_X1 U91 (.ZN(n119), 
	.B2(n17116), 
	.B1(n16679), 
	.A(n17120));
   OAI211_X1 U92 (.ZN(n5675), 
	.C2(n29), 
	.C1(n122), 
	.B(n124), 
	.A(n123));
   AOI22_X1 U93 (.ZN(n124), 
	.B2(vis_pc_o[10]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_10_));
   AOI21_X1 U95 (.ZN(n123), 
	.B2(n17116), 
	.B1(n16719), 
	.A(n17120));
   INV_X1 U96 (.ZN(n122), 
	.A(n126));
   OAI211_X1 U97 (.ZN(n5676), 
	.C2(n29), 
	.C1(n127), 
	.B(n129), 
	.A(n128));
   AOI22_X1 U98 (.ZN(n129), 
	.B2(vis_pc_o[8]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_8_));
   AOI21_X1 U100 (.ZN(n128), 
	.B2(n17116), 
	.B1(n16727), 
	.A(n17120));
   OAI211_X1 U101 (.ZN(n5677), 
	.C2(n29), 
	.C1(n131), 
	.B(n133), 
	.A(n132));
   AOI22_X1 U102 (.ZN(n133), 
	.B2(vis_pc_o[13]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_13_));
   AOI21_X1 U104 (.ZN(n132), 
	.B2(n17116), 
	.B1(n16658), 
	.A(n17120));
   INV_X1 U105 (.ZN(n131), 
	.A(n135));
   OAI211_X1 U106 (.ZN(n5678), 
	.C2(n29), 
	.C1(n136), 
	.B(n138), 
	.A(n137));
   AOI22_X1 U107 (.ZN(n138), 
	.B2(vis_pc_o[11]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_11_));
   AOI21_X1 U109 (.ZN(n137), 
	.B2(n17116), 
	.B1(n16653), 
	.A(n17120));
   OAI211_X1 U110 (.ZN(n5679), 
	.C2(n29), 
	.C1(FE_PHN770_n140), 
	.B(n142), 
	.A(n141));
   AOI22_X1 U111 (.ZN(n142), 
	.B2(vis_pc_o[9]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_9_));
   AOI21_X1 U113 (.ZN(n141), 
	.B2(n17116), 
	.B1(n16723), 
	.A(n17120));
   OAI211_X1 U114 (.ZN(n5680), 
	.C2(n29), 
	.C1(n144), 
	.B(n146), 
	.A(n145));
   AOI22_X1 U115 (.ZN(n146), 
	.B2(vis_pc_o[7]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_7_));
   AOI21_X1 U116 (.ZN(n145), 
	.B2(n17116), 
	.B1(n16722), 
	.A(n17120));
   OAI211_X1 U117 (.ZN(n5681), 
	.C2(n29), 
	.C1(n148), 
	.B(n150), 
	.A(n149));
   AOI22_X1 U118 (.ZN(n150), 
	.B2(FE_PHN1339_SYNOPSYS_UNCONNECTED_540), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_5_));
   AOI21_X1 U119 (.ZN(n149), 
	.B2(n17116), 
	.B1(add_2073_SUM_7_), 
	.A(n17120));
   OAI211_X1 U120 (.ZN(n5682), 
	.C2(n29), 
	.C1(FE_PHN783_n152), 
	.B(n154), 
	.A(n153));
   AOI22_X1 U121 (.ZN(n154), 
	.B2(vis_pc_o[4]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_4_));
   AOI21_X1 U122 (.ZN(n153), 
	.B2(n17116), 
	.B1(n16731), 
	.A(n17120));
   OAI222_X1 U123 (.ZN(n5683), 
	.C2(n159), 
	.C1(n158), 
	.B2(n157), 
	.B1(n5240), 
	.A2(n156), 
	.A1(FE_PHN783_n152));
   OAI211_X1 U125 (.ZN(n5684), 
	.C2(n29), 
	.C1(FE_PHN778_n160), 
	.B(n162), 
	.A(n161));
   AOI22_X1 U126 (.ZN(n162), 
	.B2(vis_pc_o[3]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_3_));
   AOI21_X1 U127 (.ZN(n161), 
	.B2(n17116), 
	.B1(n16730), 
	.A(n17120));
   OAI222_X1 U128 (.ZN(n5685), 
	.C2(n165), 
	.C1(n158), 
	.B2(n164), 
	.B1(n157), 
	.A2(n156), 
	.A1(FE_PHN778_n160));
   OAI211_X1 U129 (.ZN(n5686), 
	.C2(n29), 
	.C1(FE_PHN693_n166), 
	.B(n168), 
	.A(n167));
   AOI22_X1 U130 (.ZN(n168), 
	.B2(vis_pc_o[2]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_2_));
   AOI21_X1 U131 (.ZN(n167), 
	.B2(n17116), 
	.B1(n16682), 
	.A(n17120));
   OAI222_X1 U132 (.ZN(n5687), 
	.C2(n170), 
	.C1(n158), 
	.B2(n157), 
	.B1(FE_PHN3500_n5099), 
	.A2(n156), 
	.A1(FE_PHN693_n166));
   OAI211_X1 U133 (.ZN(n5688), 
	.C2(n29), 
	.C1(FE_PHN2916_n171), 
	.B(n173), 
	.A(n172));
   AOI22_X1 U134 (.ZN(n173), 
	.B2(vis_pc_o[1]), 
	.B1(n42), 
	.A2(n17117), 
	.A1(add_2071_SUM_1_));
   AOI21_X1 U136 (.ZN(n172), 
	.B2(n17116), 
	.B1(n16729), 
	.A(n17120));
   OAI222_X1 U138 (.ZN(n5689), 
	.C2(n176), 
	.C1(n158), 
	.B2(n175), 
	.B1(n157), 
	.A2(n156), 
	.A1(FE_PHN2916_n171));
   OAI221_X1 U139 (.ZN(n5690), 
	.C2(n37), 
	.C1(n4973), 
	.B2(vis_pc_o[0]), 
	.B1(n36), 
	.A(n178));
   AOI221_X1 U140 (.ZN(n178), 
	.C2(n17116), 
	.C1(n16732), 
	.B2(n179), 
	.B1(n54), 
	.A(n17120));
   OAI221_X1 U142 (.ZN(n180), 
	.C2(n184), 
	.C1(n183), 
	.B2(n182), 
	.B1(n181), 
	.A(n185));
   OR2_X1 U143 (.ZN(n182), 
	.A2(n5234), 
	.A1(n186));
   NAND2_X1 U146 (.ZN(n36), 
	.A2(n37), 
	.A1(n189));
   OAI222_X1 U147 (.ZN(n5691), 
	.C2(n191), 
	.C1(n158), 
	.B2(n157), 
	.B1(n5025), 
	.A2(n156), 
	.A1(FE_PHN719_n190));
   OAI222_X1 U148 (.ZN(n5692), 
	.C2(n186), 
	.C1(n158), 
	.B2(n157), 
	.B1(n4966), 
	.A2(n156), 
	.A1(n192));
   NAND2_X1 U149 (.ZN(n157), 
	.A2(n194), 
	.A1(n193));
   NAND2_X1 U150 (.ZN(n156), 
	.A2(n195), 
	.A1(n158));
   INV_X1 U151 (.ZN(n158), 
	.A(n196));
   NAND2_X1 U152 (.ZN(n5693), 
	.A2(n198), 
	.A1(n197));
   OAI221_X1 U153 (.ZN(n198), 
	.C2(n202), 
	.C1(n201), 
	.B2(n200), 
	.B1(n199), 
	.A(n203));
   INV_X1 U154 (.ZN(n197), 
	.A(n204));
   OAI21_X1 U155 (.ZN(n5694), 
	.B2(n202), 
	.B1(n205), 
	.A(n206));
   OAI221_X1 U156 (.ZN(n206), 
	.C2(n202), 
	.C1(n208), 
	.B2(n200), 
	.B1(n207), 
	.A(n209));
   OAI21_X1 U157 (.ZN(n5695), 
	.B2(n211), 
	.B1(n210), 
	.A(n212));
   OAI21_X1 U158 (.ZN(n212), 
	.B2(n210), 
	.B1(n213), 
	.A(FE_PHN2035_n214));
   OAI21_X1 U160 (.ZN(n5696), 
	.B2(n211), 
	.B1(n215), 
	.A(FE_PHN2047_n216));
   OAI21_X1 U161 (.ZN(n216), 
	.B2(n213), 
	.B1(n215), 
	.A(n217));
   OAI21_X1 U162 (.ZN(n5697), 
	.B2(n218), 
	.B1(n211), 
	.A(n219));
   OAI21_X1 U163 (.ZN(n219), 
	.B2(n218), 
	.B1(n213), 
	.A(FE_PHN2041_n220));
   OAI21_X1 U164 (.ZN(n5698), 
	.B2(n221), 
	.B1(n211), 
	.A(FE_PHN3411_n222));
   OAI21_X1 U165 (.ZN(n222), 
	.B2(n221), 
	.B1(n213), 
	.A(n223));
   OAI21_X1 U166 (.ZN(n5699), 
	.B2(n224), 
	.B1(n211), 
	.A(n225));
   OAI21_X1 U167 (.ZN(n225), 
	.B2(n224), 
	.B1(n213), 
	.A(n4799));
   OAI21_X1 U168 (.ZN(n5700), 
	.B2(n226), 
	.B1(n211), 
	.A(FE_PHN2048_n227));
   OAI21_X1 U169 (.ZN(n227), 
	.B2(n226), 
	.B1(n213), 
	.A(n228));
   OAI21_X1 U170 (.ZN(n5701), 
	.B2(n229), 
	.B1(n211), 
	.A(FE_PHN2043_n230));
   OAI21_X1 U171 (.ZN(n230), 
	.B2(n229), 
	.B1(n213), 
	.A(n231));
   OAI22_X1 U172 (.ZN(n5702), 
	.B2(n233), 
	.B1(n4796), 
	.A2(n211), 
	.A1(n232));
   NOR2_X1 U173 (.ZN(n233), 
	.A2(n213), 
	.A1(n232));
   OAI22_X1 U174 (.ZN(n5703), 
	.B2(n235), 
	.B1(n5578), 
	.A2(n211), 
	.A1(n234));
   NOR2_X1 U175 (.ZN(n235), 
	.A2(n213), 
	.A1(n234));
   OAI22_X1 U176 (.ZN(n5704), 
	.B2(n237), 
	.B1(n5537), 
	.A2(n211), 
	.A1(n236));
   NOR2_X1 U177 (.ZN(n237), 
	.A2(n213), 
	.A1(n236));
   OAI22_X1 U178 (.ZN(n5705), 
	.B2(n239), 
	.B1(n5570), 
	.A2(n211), 
	.A1(n238));
   NOR2_X1 U179 (.ZN(n239), 
	.A2(n213), 
	.A1(n238));
   OAI22_X1 U180 (.ZN(n5706), 
	.B2(n241), 
	.B1(n4795), 
	.A2(n211), 
	.A1(n240));
   NOR2_X1 U181 (.ZN(n241), 
	.A2(n213), 
	.A1(n240));
   OAI22_X1 U182 (.ZN(n5707), 
	.B2(n244), 
	.B1(n243), 
	.A2(n211), 
	.A1(n242));
   NOR2_X1 U183 (.ZN(n243), 
	.A2(n213), 
	.A1(n242));
   OAI22_X1 U184 (.ZN(n5708), 
	.B2(n246), 
	.B1(FE_PHN2672_n5538), 
	.A2(n245), 
	.A1(n211));
   NOR2_X1 U185 (.ZN(n246), 
	.A2(n245), 
	.A1(n213));
   OAI22_X1 U186 (.ZN(n5709), 
	.B2(n248), 
	.B1(FE_PHN2675_n5539), 
	.A2(n247), 
	.A1(n211));
   NOR2_X1 U187 (.ZN(n248), 
	.A2(n247), 
	.A1(n213));
   OAI22_X1 U188 (.ZN(n5710), 
	.B2(n250), 
	.B1(n5540), 
	.A2(n249), 
	.A1(n211));
   NOR2_X1 U189 (.ZN(n250), 
	.A2(n249), 
	.A1(n213));
   OAI211_X1 U192 (.ZN(n5711), 
	.C2(n17122), 
	.C1(n4905), 
	.B(n255), 
	.A(n254));
   OAI21_X1 U193 (.ZN(n254), 
	.B2(haddr_o[2]), 
	.B1(haddr_o[7]), 
	.A(n256));
   OAI33_X1 U194 (.ZN(n5712), 
	.B3(n260), 
	.B2(FE_PHN3501_n5516), 
	.B1(n259), 
	.A3(n258), 
	.A2(n5068), 
	.A1(n257));
   NOR3_X1 U195 (.ZN(n257), 
	.A3(n261), 
	.A2(n251), 
	.A1(n253));
   OAI221_X1 U196 (.ZN(n5713), 
	.C2(n17107), 
	.C1(n264), 
	.B2(n17109), 
	.B1(FE_PHN3496_n262), 
	.A(n266));
   NAND2_X1 U199 (.ZN(n269), 
	.A2(n17106), 
	.A1(sub_2068_SUM_22_));
   OAI221_X1 U201 (.ZN(n5715), 
	.C2(n17107), 
	.C1(FE_PHN3808_n270), 
	.B2(n17109), 
	.B1(FE_PHN2385_n5625), 
	.A(n271));
   NAND2_X1 U202 (.ZN(n271), 
	.A2(n17106), 
	.A1(sub_2068_SUM_21_));
   OAI221_X1 U203 (.ZN(n5716), 
	.C2(n265), 
	.C1(n272), 
	.B2(n17109), 
	.B1(FE_PHN2378_n5618), 
	.A(n273));
   NAND2_X1 U204 (.ZN(n273), 
	.A2(n17106), 
	.A1(sub_2068_SUM_20_));
   OAI221_X1 U205 (.ZN(n5717), 
	.C2(n265), 
	.C1(n274), 
	.B2(n17109), 
	.B1(FE_PHN2245_n5033), 
	.A(n275));
   NAND2_X1 U206 (.ZN(n275), 
	.A2(n17106), 
	.A1(sub_2068_SUM_19_));
   OAI221_X1 U207 (.ZN(n5718), 
	.C2(n265), 
	.C1(FE_PHN4748_n276), 
	.B2(n17109), 
	.B1(FE_PHN2270_n5067), 
	.A(n277));
   NAND2_X1 U208 (.ZN(n277), 
	.A2(n17106), 
	.A1(sub_2068_SUM_18_));
   OAI221_X1 U209 (.ZN(n5719), 
	.C2(n17107), 
	.C1(FE_PHN3717_n278), 
	.B2(n17109), 
	.B1(FE_PHN2364_n5639), 
	.A(n279));
   NAND2_X1 U210 (.ZN(n279), 
	.A2(n17106), 
	.A1(sub_2068_SUM_17_));
   NAND2_X1 U212 (.ZN(n281), 
	.A2(n17106), 
	.A1(sub_2068_SUM_16_));
   OAI221_X1 U214 (.ZN(n5721), 
	.C2(n265), 
	.C1(FE_PHN3641_n282), 
	.B2(n17109), 
	.B1(FE_PHN2429_n5505), 
	.A(n283));
   NAND2_X1 U215 (.ZN(n283), 
	.A2(n17106), 
	.A1(sub_2068_SUM_15_));
   OAI221_X1 U216 (.ZN(n5722), 
	.C2(n265), 
	.C1(FE_PHN3735_n284), 
	.B2(n17109), 
	.B1(FE_PHN2106_n5506), 
	.A(n285));
   NAND2_X1 U217 (.ZN(n285), 
	.A2(n17106), 
	.A1(sub_2068_SUM_14_));
   OAI221_X1 U218 (.ZN(n5723), 
	.C2(n265), 
	.C1(FE_PHN3779_n286), 
	.B2(n17109), 
	.B1(FE_PHN2333_n5600), 
	.A(n287));
   NAND2_X1 U219 (.ZN(n287), 
	.A2(n17106), 
	.A1(sub_2068_SUM_13_));
   OAI221_X1 U220 (.ZN(n5724), 
	.C2(n17107), 
	.C1(FE_PHN3611_n288), 
	.B2(n17109), 
	.B1(FE_PHN2428_n5507), 
	.A(n289));
   NAND2_X1 U221 (.ZN(n289), 
	.A2(n17106), 
	.A1(sub_2068_SUM_12_));
   NAND2_X1 U223 (.ZN(n291), 
	.A2(n17106), 
	.A1(sub_2068_SUM_11_));
   NAND2_X1 U226 (.ZN(n293), 
	.A2(n17106), 
	.A1(sub_2068_SUM_10_));
   OAI221_X1 U228 (.ZN(n5727), 
	.C2(n17107), 
	.C1(FE_PHN3631_n294), 
	.B2(n17109), 
	.B1(FE_PHN2330_n5579), 
	.A(n295));
   NAND2_X1 U229 (.ZN(n295), 
	.A2(n17106), 
	.A1(sub_2068_SUM_9_));
   OAI221_X1 U230 (.ZN(n5728), 
	.C2(n17107), 
	.C1(n296), 
	.B2(n17109), 
	.B1(FE_PHN2426_n5581), 
	.A(n297));
   NAND2_X1 U231 (.ZN(n297), 
	.A2(n17106), 
	.A1(sub_2068_SUM_8_));
   OAI221_X1 U232 (.ZN(n5729), 
	.C2(n17107), 
	.C1(n298), 
	.B2(n17109), 
	.B1(FE_PHN2430_n5520), 
	.A(n299));
   NAND2_X1 U233 (.ZN(n299), 
	.A2(n17106), 
	.A1(sub_2068_SUM_7_));
   NAND2_X1 U235 (.ZN(n301), 
	.A2(n17106), 
	.A1(sub_2068_SUM_6_));
   NAND2_X1 U238 (.ZN(n303), 
	.A2(n17106), 
	.A1(sub_2068_SUM_5_));
   NAND2_X1 U241 (.ZN(n305), 
	.A2(n17106), 
	.A1(sub_2068_SUM_4_));
   OAI221_X1 U243 (.ZN(n5733), 
	.C2(n17107), 
	.C1(n306), 
	.B2(n17109), 
	.B1(FE_PHN2347_n5513), 
	.A(n307));
   NAND2_X1 U244 (.ZN(n307), 
	.A2(n17106), 
	.A1(sub_2068_SUM_3_));
   OAI221_X1 U245 (.ZN(n5734), 
	.C2(n265), 
	.C1(n308), 
	.B2(n17109), 
	.B1(FE_PHN2412_n5512), 
	.A(n309));
   NAND2_X1 U246 (.ZN(n309), 
	.A2(n17106), 
	.A1(sub_2068_SUM_2_));
   OAI221_X1 U247 (.ZN(n5735), 
	.C2(n265), 
	.C1(n310), 
	.B2(n17109), 
	.B1(FE_PHN2232_n5511), 
	.A(n311));
   NAND2_X1 U248 (.ZN(n311), 
	.A2(n17106), 
	.A1(sub_2068_SUM_1_));
   OAI222_X1 U249 (.ZN(n5736), 
	.C2(n17107), 
	.C1(n260), 
	.B2(n16647), 
	.B1(sub_2068_A_0_), 
	.A2(n17109), 
	.A1(FE_PHN3512_n5510));
   INV_X1 U252 (.ZN(n258), 
	.A(n315));
   NOR2_X1 U255 (.ZN(n314), 
	.A2(sub_2068_A_0_), 
	.A1(n259));
   NAND2_X1 U256 (.ZN(n265), 
	.A2(n315), 
	.A1(FE_PHN3501_n5516));
   NAND2_X1 U257 (.ZN(n315), 
	.A2(n253), 
	.A1(n316));
   OAI221_X1 U258 (.ZN(n5737), 
	.C2(n17102), 
	.C1(n4971), 
	.B2(n17103), 
	.B1(n317), 
	.A(n320));
   AOI22_X1 U259 (.ZN(n320), 
	.B2(vis_tbit_o), 
	.B1(n322), 
	.A2(FE_PHN1331_SYNOPSYS_UNCONNECTED_522), 
	.A1(n16738));
   OAI221_X1 U261 (.ZN(n5738), 
	.C2(n17102), 
	.C1(n5101), 
	.B2(n324), 
	.B1(n186), 
	.A(n325));
   OAI21_X1 U262 (.ZN(n325), 
	.B2(n327), 
	.B1(n326), 
	.A(n17104));
   AOI21_X1 U263 (.ZN(n326), 
	.B2(n330), 
	.B1(n329), 
	.A(n4922));
   NAND3_X1 U264 (.ZN(n330), 
	.A3(n333), 
	.A2(n16686), 
	.A1(n16657));
   OAI221_X1 U265 (.ZN(n5739), 
	.C2(n336), 
	.C1(n16803), 
	.B2(n335), 
	.B1(n334), 
	.A(n337));
   AOI222_X1 U266 (.ZN(n337), 
	.C2(hrdata_i[14]), 
	.C1(n341), 
	.B2(hrdata_i[30]), 
	.B1(n16646), 
	.A2(n339), 
	.A1(n338));
   OAI221_X1 U268 (.ZN(n5740), 
	.C2(n336), 
	.C1(n16795), 
	.B2(n334), 
	.B1(n3), 
	.A(n342));
   AOI222_X1 U269 (.ZN(n342), 
	.C2(hrdata_i[12]), 
	.C1(n341), 
	.B2(hrdata_i[28]), 
	.B1(n16646), 
	.A2(n343), 
	.A1(n338));
   OAI221_X1 U271 (.ZN(n5741), 
	.C2(n336), 
	.C1(n16814), 
	.B2(n334), 
	.B1(n4), 
	.A(n344));
   AOI222_X1 U272 (.ZN(n344), 
	.C2(hrdata_i[11]), 
	.C1(n341), 
	.B2(hrdata_i[27]), 
	.B1(n16646), 
	.A2(n345), 
	.A1(n338));
   OAI221_X1 U274 (.ZN(n5742), 
	.C2(n336), 
	.C1(n16816), 
	.B2(n334), 
	.B1(n5), 
	.A(n346));
   AOI222_X1 U275 (.ZN(n346), 
	.C2(hrdata_i[10]), 
	.C1(n341), 
	.B2(hrdata_i[26]), 
	.B1(n16646), 
	.A2(n347), 
	.A1(n338));
   OAI221_X1 U277 (.ZN(n5743), 
	.C2(n336), 
	.C1(n16796), 
	.B2(n334), 
	.B1(n6), 
	.A(n348));
   AOI222_X1 U278 (.ZN(n348), 
	.C2(hrdata_i[9]), 
	.C1(n341), 
	.B2(hrdata_i[25]), 
	.B1(n16646), 
	.A2(n349), 
	.A1(n338));
   OAI221_X1 U280 (.ZN(n5744), 
	.C2(n336), 
	.C1(n16797), 
	.B2(n334), 
	.B1(n7), 
	.A(n350));
   AOI222_X1 U281 (.ZN(n350), 
	.C2(hrdata_i[8]), 
	.C1(n341), 
	.B2(hrdata_i[24]), 
	.B1(n16646), 
	.A2(n351), 
	.A1(n338));
   OAI221_X1 U283 (.ZN(n5745), 
	.C2(n336), 
	.C1(n16799), 
	.B2(n334), 
	.B1(n8), 
	.A(n352));
   AOI222_X1 U284 (.ZN(n352), 
	.C2(hrdata_i[7]), 
	.C1(n341), 
	.B2(hrdata_i[23]), 
	.B1(n16646), 
	.A2(n353), 
	.A1(n338));
   OAI221_X1 U286 (.ZN(n5746), 
	.C2(n336), 
	.C1(n16801), 
	.B2(n334), 
	.B1(n9), 
	.A(n354));
   AOI222_X1 U287 (.ZN(n354), 
	.C2(hrdata_i[6]), 
	.C1(n341), 
	.B2(hrdata_i[22]), 
	.B1(n16646), 
	.A2(n355), 
	.A1(n338));
   OAI221_X1 U289 (.ZN(n5747), 
	.C2(n336), 
	.C1(n5244), 
	.B2(n334), 
	.B1(n5240), 
	.A(n356));
   AOI222_X1 U290 (.ZN(n356), 
	.C2(hrdata_i[5]), 
	.C1(n341), 
	.B2(hrdata_i[21]), 
	.B1(n16646), 
	.A2(n357), 
	.A1(n338));
   OAI221_X1 U292 (.ZN(n5748), 
	.C2(n336), 
	.C1(n5243), 
	.B2(n334), 
	.B1(n164), 
	.A(n358));
   AOI222_X1 U293 (.ZN(n358), 
	.C2(hrdata_i[4]), 
	.C1(n341), 
	.B2(hrdata_i[20]), 
	.B1(n16646), 
	.A2(n359), 
	.A1(n338));
   OAI221_X1 U295 (.ZN(n5749), 
	.C2(n336), 
	.C1(n16794), 
	.B2(n334), 
	.B1(FE_PHN3500_n5099), 
	.A(n360));
   AOI222_X1 U296 (.ZN(n360), 
	.C2(hrdata_i[3]), 
	.C1(n341), 
	.B2(hrdata_i[19]), 
	.B1(n16646), 
	.A2(n361), 
	.A1(n338));
   OAI221_X1 U298 (.ZN(n5750), 
	.C2(n336), 
	.C1(n5241), 
	.B2(n334), 
	.B1(n175), 
	.A(n362));
   AOI222_X1 U299 (.ZN(n362), 
	.C2(hrdata_i[2]), 
	.C1(n341), 
	.B2(hrdata_i[18]), 
	.B1(n16646), 
	.A2(n363), 
	.A1(n338));
   OAI221_X1 U301 (.ZN(n5751), 
	.C2(n336), 
	.C1(n5026), 
	.B2(n334), 
	.B1(n5025), 
	.A(n364));
   AOI222_X1 U302 (.ZN(n364), 
	.C2(hrdata_i[1]), 
	.C1(n341), 
	.B2(hrdata_i[17]), 
	.B1(n16646), 
	.A2(n365), 
	.A1(n338));
   OAI221_X1 U304 (.ZN(n5752), 
	.C2(n336), 
	.C1(n4967), 
	.B2(n334), 
	.B1(n4966), 
	.A(n366));
   AOI222_X1 U305 (.ZN(n366), 
	.C2(hrdata_i[0]), 
	.C1(n341), 
	.B2(hrdata_i[16]), 
	.B1(n16646), 
	.A2(n367), 
	.A1(n338));
   OAI221_X1 U307 (.ZN(n5753), 
	.C2(n336), 
	.C1(n16807), 
	.B2(n334), 
	.B1(n2), 
	.A(n368));
   AOI222_X1 U308 (.ZN(n368), 
	.C2(hrdata_i[13]), 
	.C1(n341), 
	.B2(hrdata_i[29]), 
	.B1(n16646), 
	.A2(n369), 
	.A1(n338));
   OAI221_X1 U310 (.ZN(n5754), 
	.C2(n336), 
	.C1(n16811), 
	.B2(n370), 
	.B1(n334), 
	.A(n371));
   AOI222_X1 U311 (.ZN(n371), 
	.C2(hrdata_i[15]), 
	.C1(n341), 
	.B2(hrdata_i[31]), 
	.B1(n16646), 
	.A2(n372), 
	.A1(n338));
   NAND2_X1 U314 (.ZN(n374), 
	.A2(vis_pc_o[0]), 
	.A1(n16868));
   OAI22_X1 U317 (.ZN(n5755), 
	.B2(n381), 
	.B1(FE_PHN4701_n380), 
	.A2(n379), 
	.A1(n335));
   INV_X1 U318 (.ZN(n380), 
	.A(hrdata_i[14]));
   OAI221_X1 U320 (.ZN(n5756), 
	.C2(n379), 
	.C1(n2), 
	.B2(n381), 
	.B1(n382), 
	.A(n383));
   NAND2_X1 U321 (.ZN(n383), 
	.A2(n384), 
	.A1(sub_2069_SUM_8_));
   OAI221_X1 U322 (.ZN(n5757), 
	.C2(n379), 
	.C1(n3), 
	.B2(n381), 
	.B1(FE_PHN4725_n385), 
	.A(n386));
   NAND2_X1 U323 (.ZN(n386), 
	.A2(n384), 
	.A1(sub_2069_SUM_7_));
   INV_X1 U324 (.ZN(n385), 
	.A(hrdata_i[12]));
   OAI221_X1 U325 (.ZN(n5758), 
	.C2(n379), 
	.C1(n4), 
	.B2(n381), 
	.B1(FE_PHN4700_n387), 
	.A(n388));
   NAND2_X1 U326 (.ZN(n388), 
	.A2(n384), 
	.A1(sub_2069_SUM_6_));
   INV_X1 U327 (.ZN(n387), 
	.A(hrdata_i[11]));
   OAI221_X1 U328 (.ZN(n5759), 
	.C2(n379), 
	.C1(n5), 
	.B2(n381), 
	.B1(FE_PHN4693_n389), 
	.A(n390));
   NAND2_X1 U329 (.ZN(n390), 
	.A2(n384), 
	.A1(sub_2069_SUM_5_));
   INV_X1 U330 (.ZN(n389), 
	.A(hrdata_i[10]));
   OAI221_X1 U331 (.ZN(n5760), 
	.C2(n379), 
	.C1(n6), 
	.B2(n381), 
	.B1(n391), 
	.A(n392));
   NAND2_X1 U332 (.ZN(n392), 
	.A2(n384), 
	.A1(sub_2069_SUM_4_));
   OAI221_X1 U333 (.ZN(n5761), 
	.C2(n379), 
	.C1(n7), 
	.B2(n381), 
	.B1(FE_PHN904_n393), 
	.A(n394));
   NAND2_X1 U334 (.ZN(n394), 
	.A2(n384), 
	.A1(sub_2069_SUM_3_));
   OAI221_X1 U335 (.ZN(n5762), 
	.C2(n379), 
	.C1(n8), 
	.B2(n381), 
	.B1(FE_PHN4695_n395), 
	.A(n396));
   NAND2_X1 U336 (.ZN(n396), 
	.A2(n384), 
	.A1(sub_2069_SUM_2_));
   INV_X1 U337 (.ZN(n395), 
	.A(hrdata_i[7]));
   OAI221_X1 U338 (.ZN(n5763), 
	.C2(n379), 
	.C1(n9), 
	.B2(n381), 
	.B1(n397), 
	.A(n398));
   NAND2_X1 U339 (.ZN(n398), 
	.A2(n384), 
	.A1(sub_2069_SUM_1_));
   AOI21_X1 U340 (.ZN(n384), 
	.B2(n5648), 
	.B1(n399), 
	.A(n400));
   OR4_X1 U341 (.ZN(n399), 
	.A4(n404), 
	.A3(n403), 
	.A2(n402), 
	.A1(n401));
   XOR2_X1 U342 (.Z(n404), 
	.B(n406), 
	.A(n405));
   NOR2_X1 U343 (.ZN(n406), 
	.A2(n164), 
	.A1(n5034));
   XOR2_X1 U344 (.Z(n402), 
	.B(n407), 
	.A(n4804));
   OAI221_X1 U345 (.ZN(n401), 
	.C2(n410), 
	.C1(n5025), 
	.B2(n409), 
	.B1(n408), 
	.A(n411));
   AOI21_X1 U346 (.ZN(n411), 
	.B2(n413), 
	.B1(n412), 
	.A(n414));
   XOR2_X1 U347 (.Z(n414), 
	.B(n416), 
	.A(n415));
   AOI21_X1 U348 (.ZN(n409), 
	.B2(n417), 
	.B1(n4966), 
	.A(n410));
   AOI211_X1 U349 (.ZN(n408), 
	.C2(n417), 
	.C1(n4966), 
	.B(n5034), 
	.A(n5025));
   OAI22_X1 U350 (.ZN(n5764), 
	.B2(n381), 
	.B1(FE_PHN3000_n419), 
	.A2(n418), 
	.A1(n5240));
   INV_X1 U351 (.ZN(n419), 
	.A(hrdata_i[5]));
   OAI222_X1 U352 (.ZN(n5765), 
	.C2(n422), 
	.C1(n421), 
	.B2(n381), 
	.B1(FE_PHN870_n420), 
	.A2(n418), 
	.A1(n164));
   OAI222_X1 U354 (.ZN(n5766), 
	.C2(n422), 
	.C1(n424), 
	.B2(n381), 
	.B1(FE_PHN875_n423), 
	.A2(n418), 
	.A1(FE_PHN3500_n5099));
   OAI222_X1 U355 (.ZN(n5767), 
	.C2(n422), 
	.C1(n426), 
	.B2(n381), 
	.B1(FE_PHN844_n425), 
	.A2(n418), 
	.A1(n175));
   OAI222_X1 U356 (.ZN(n5768), 
	.C2(n422), 
	.C1(n428), 
	.B2(n381), 
	.B1(FE_PHN869_n427), 
	.A2(n418), 
	.A1(n5025));
   INV_X1 U357 (.ZN(n428), 
	.A(n410));
   OAI222_X1 U358 (.ZN(n5769), 
	.C2(n422), 
	.C1(n412), 
	.B2(n381), 
	.B1(FE_PHN804_n429), 
	.A2(n418), 
	.A1(n4966));
   OAI21_X1 U360 (.ZN(n418), 
	.B2(n431), 
	.B1(n430), 
	.A(n422));
   OAI221_X1 U361 (.ZN(n5770), 
	.C2(n434), 
	.C1(n5254), 
	.B2(n433), 
	.B1(n432), 
	.A(n435));
   AOI21_X1 U362 (.ZN(n434), 
	.B2(n437), 
	.B1(n436), 
	.A(n433));
   AOI221_X1 U363 (.ZN(n432), 
	.C2(n16817), 
	.C1(n440), 
	.B2(n16734), 
	.B1(n438), 
	.A(n442));
   OAI33_X1 U364 (.ZN(n442), 
	.B3(n445), 
	.B2(n16814), 
	.B1(n16681), 
	.A3(n444), 
	.A2(n16795), 
	.A1(n443));
   OAI221_X1 U365 (.ZN(n5771), 
	.C2(n447), 
	.C1(n5162), 
	.B2(n433), 
	.B1(n446), 
	.A(n435));
   AOI222_X1 U366 (.ZN(n446), 
	.C2(n451), 
	.C1(n450), 
	.B2(n17098), 
	.B1(n449), 
	.A2(n16798), 
	.A1(n440));
   OAI221_X1 U367 (.ZN(n5772), 
	.C2(n433), 
	.C1(n453), 
	.B2(n452), 
	.B1(n5253), 
	.A(n435));
   AOI222_X1 U368 (.ZN(n453), 
	.C2(n454), 
	.C1(n450), 
	.B2(n16817), 
	.B1(n449), 
	.A2(n16657), 
	.A1(n440));
   AOI21_X1 U369 (.ZN(n452), 
	.B2(n455), 
	.B1(n436), 
	.A(n433));
   OAI221_X1 U370 (.ZN(n5773), 
	.C2(n433), 
	.C1(n457), 
	.B2(n456), 
	.B1(n5003), 
	.A(n435));
   NAND2_X1 U371 (.ZN(n435), 
	.A2(n458), 
	.A1(n447));
   OAI21_X1 U372 (.ZN(n458), 
	.B2(n459), 
	.B1(n16799), 
	.A(n460));
   INV_X1 U373 (.ZN(n447), 
	.A(n433));
   AOI222_X1 U374 (.ZN(n457), 
	.C2(n461), 
	.C1(n450), 
	.B2(n16657), 
	.B1(n449), 
	.A2(n17098), 
	.A1(n440));
   NAND3_X1 U375 (.ZN(n450), 
	.A3(n464), 
	.A2(n463), 
	.A1(n462));
   AOI21_X1 U376 (.ZN(n464), 
	.B2(n466), 
	.B1(n465), 
	.A(n438));
   NAND2_X1 U377 (.ZN(n438), 
	.A2(n468), 
	.A1(n467));
   NAND3_X1 U378 (.ZN(n467), 
	.A3(n471), 
	.A2(n16725), 
	.A1(n469));
   AOI21_X1 U379 (.ZN(n471), 
	.B2(n16657), 
	.B1(n16733), 
	.A(n443));
   OAI211_X1 U380 (.ZN(n463), 
	.C2(n474), 
	.C1(n473), 
	.B(n475), 
	.A(n16820));
   NAND3_X1 U381 (.ZN(n462), 
	.A3(n476), 
	.A2(n16725), 
	.A1(n16816));
   OAI221_X1 U382 (.ZN(n449), 
	.C2(n479), 
	.C1(n478), 
	.B2(n443), 
	.B1(n477), 
	.A(n480));
   AOI22_X1 U383 (.ZN(n480), 
	.B2(n466), 
	.B1(n482), 
	.A2(n481), 
	.A1(n16820));
   INV_X1 U384 (.ZN(n481), 
	.A(n445));
   NOR2_X1 U385 (.ZN(n445), 
	.A2(n484), 
	.A1(n483));
   NOR2_X1 U386 (.ZN(n477), 
	.A2(n16795), 
	.A1(n485));
   AOI21_X1 U387 (.ZN(n456), 
	.B2(n486), 
	.B1(n436), 
	.A(n433));
   NAND2_X1 U388 (.ZN(n433), 
	.A2(n487), 
	.A1(n17124));
   NAND4_X1 U389 (.ZN(n487), 
	.A4(n491), 
	.A3(n490), 
	.A2(n489), 
	.A1(n488));
   NOR4_X1 U390 (.ZN(n491), 
	.A4(n495), 
	.A3(n494), 
	.A2(n493), 
	.A1(n492));
   OAI221_X1 U391 (.ZN(n492), 
	.C2(n499), 
	.C1(n498), 
	.B2(n497), 
	.B1(n496), 
	.A(n500));
   NAND4_X1 U392 (.ZN(n500), 
	.A4(FE_OFN21_n503), 
	.A3(n502), 
	.A2(n501), 
	.A1(n483));
   AOI21_X1 U393 (.ZN(n496), 
	.B2(n16817), 
	.B1(n504), 
	.A(n505));
   AOI221_X1 U394 (.ZN(n490), 
	.C2(n16802), 
	.C1(n508), 
	.B2(n507), 
	.B1(n506), 
	.A(n510));
   OAI211_X1 U395 (.ZN(n508), 
	.C2(n329), 
	.C1(n16733), 
	.B(n512), 
	.A(n511));
   NAND3_X1 U396 (.ZN(n511), 
	.A3(n16811), 
	.A2(n16871), 
	.A1(n16733));
   AOI21_X1 U397 (.ZN(n436), 
	.B2(n17097), 
	.B1(n514), 
	.A(n515));
   OAI22_X1 U398 (.ZN(n5774), 
	.B2(FE_PHN675_n17126), 
	.B1(n516), 
	.A2(FE_OFN667_n17122), 
	.A1(n16854));
   NOR4_X1 U399 (.ZN(n516), 
	.A4(n520), 
	.A3(n519), 
	.A2(n518), 
	.A1(n517));
   OAI221_X1 U400 (.ZN(n520), 
	.C2(n524), 
	.C1(n16864), 
	.B2(n522), 
	.B1(n16859), 
	.A(n525));
   AOI22_X1 U401 (.ZN(n525), 
	.B2(n529), 
	.B1(n528), 
	.A2(n527), 
	.A1(n526));
   OAI221_X1 U402 (.ZN(n519), 
	.C2(n532), 
	.C1(n531), 
	.B2(n530), 
	.B1(n16795), 
	.A(n533));
   AOI222_X1 U403 (.ZN(n533), 
	.C2(n538), 
	.C1(n16820), 
	.B2(n537), 
	.B1(n536), 
	.A2(n535), 
	.A1(n534));
   INV_X1 U404 (.ZN(n538), 
	.A(n539));
   AOI221_X1 U405 (.ZN(n539), 
	.C2(n543), 
	.C1(n542), 
	.B2(n541), 
	.B1(n540), 
	.A(n544));
   OR2_X1 U406 (.ZN(n544), 
	.A2(n546), 
	.A1(n545));
   NAND3_X1 U407 (.ZN(n537), 
	.A3(n549), 
	.A2(n548), 
	.A1(n547));
   NAND3_X1 U408 (.ZN(n549), 
	.A3(n551), 
	.A2(n16797), 
	.A1(n550));
   INV_X1 U409 (.ZN(n536), 
	.A(n552));
   AOI211_X1 U410 (.ZN(n531), 
	.C2(n553), 
	.C1(n466), 
	.B(n555), 
	.A(n554));
   AOI21_X1 U411 (.ZN(n555), 
	.B2(n557), 
	.B1(n556), 
	.A(n558));
   OAI21_X1 U412 (.ZN(n557), 
	.B2(n16824), 
	.B1(n559), 
	.A(n16862));
   NAND2_X1 U413 (.ZN(n554), 
	.A2(n561), 
	.A1(n560));
   NAND3_X1 U414 (.ZN(n561), 
	.A3(n563), 
	.A2(FE_OFN85_n16839), 
	.A1(n16820));
   OAI21_X1 U415 (.ZN(n560), 
	.B2(n565), 
	.B1(n564), 
	.A(n566));
   INV_X1 U416 (.ZN(n564), 
	.A(n567));
   OAI21_X1 U417 (.ZN(n553), 
	.B2(n569), 
	.B1(n568), 
	.A(n570));
   NAND3_X1 U418 (.ZN(n570), 
	.A3(n5228), 
	.A2(n16826), 
	.A1(FE_OFN628_n16833));
   AOI221_X1 U419 (.ZN(n530), 
	.C2(n473), 
	.C1(n574), 
	.B2(n573), 
	.B1(n572), 
	.A(n575));
   OAI33_X1 U420 (.ZN(n575), 
	.B3(n580), 
	.B2(n579), 
	.B1(n578), 
	.A3(n577), 
	.A2(n5243), 
	.A1(n576));
   NAND2_X1 U421 (.ZN(n578), 
	.A2(n581), 
	.A1(n16680));
   OAI22_X1 U422 (.ZN(n581), 
	.B2(n583), 
	.B1(n16796), 
	.A2(n582), 
	.A1(n16797));
   OAI21_X1 U423 (.ZN(n573), 
	.B2(n16812), 
	.B1(n16801), 
	.A(n16798));
   OAI221_X1 U424 (.ZN(n518), 
	.C2(n586), 
	.C1(FE_OFN70_n16867), 
	.B2(FE_OFN107_n585), 
	.B1(n584), 
	.A(n587));
   AOI222_X1 U425 (.ZN(n587), 
	.C2(n593), 
	.C1(n592), 
	.B2(n591), 
	.B1(n590), 
	.A2(n589), 
	.A1(n588));
   OAI22_X1 U426 (.ZN(n593), 
	.B2(n596), 
	.B1(n595), 
	.A2(n16734), 
	.A1(n594));
   AOI221_X1 U427 (.ZN(n595), 
	.C2(n598), 
	.C1(n16833), 
	.B2(n16862), 
	.B1(n597), 
	.A(n599));
   OAI21_X1 U428 (.ZN(n598), 
	.B2(n16839), 
	.B1(n16680), 
	.A(n600));
   OAI21_X1 U429 (.ZN(n600), 
	.B2(n602), 
	.B1(n601), 
	.A(n483));
   INV_X1 U430 (.ZN(n601), 
	.A(n603));
   OAI21_X1 U431 (.ZN(n591), 
	.B2(n605), 
	.B1(n604), 
	.A(n606));
   INV_X1 U432 (.ZN(n588), 
	.A(n607));
   AOI222_X1 U433 (.ZN(n586), 
	.C2(n589), 
	.C1(n611), 
	.B2(n610), 
	.B1(n609), 
	.A2(n563), 
	.A1(n608));
   AOI221_X1 U434 (.ZN(n584), 
	.C2(n614), 
	.C1(n613), 
	.B2(n5228), 
	.B1(n612), 
	.A(n615));
   NOR2_X1 U435 (.ZN(n613), 
	.A2(n617), 
	.A1(n616));
   NAND4_X1 U436 (.ZN(n517), 
	.A4(n621), 
	.A3(n620), 
	.A2(n619), 
	.A1(n618));
   AOI21_X1 U437 (.ZN(n621), 
	.B2(n622), 
	.B1(n574), 
	.A(n623));
   NOR4_X1 U438 (.ZN(n623), 
	.A4(n625), 
	.A3(FE_OFN21_n503), 
	.A2(n579), 
	.A1(n624));
   OAI21_X1 U439 (.ZN(n622), 
	.B2(n626), 
	.B1(n16812), 
	.A(n627));
   AOI21_X1 U440 (.ZN(n626), 
	.B2(n16657), 
	.B1(FE_OFN419_n628), 
	.A(n629));
   NAND4_X1 U441 (.ZN(n620), 
	.A4(n632), 
	.A3(n483), 
	.A2(n631), 
	.A1(n630));
   OAI22_X1 U442 (.ZN(n5775), 
	.B2(FE_PHN675_n17126), 
	.B1(n633), 
	.A2(FE_OFN667_n17122), 
	.A1(n16868));
   NOR4_X1 U443 (.ZN(n633), 
	.A4(n637), 
	.A3(n636), 
	.A2(n635), 
	.A1(n634));
   OAI221_X1 U444 (.ZN(n637), 
	.C2(FE_OFN422_n641), 
	.C1(n640), 
	.B2(n639), 
	.B1(n638), 
	.A(n642));
   OAI222_X1 U445 (.ZN(n636), 
	.C2(n648), 
	.C1(n647), 
	.B2(n646), 
	.B1(FE_OFN627_n16828), 
	.A2(n644), 
	.A1(n643));
   INV_X1 U446 (.ZN(n647), 
	.A(n535));
   OAI21_X1 U447 (.ZN(n535), 
	.B2(n514), 
	.B1(n649), 
	.A(n650));
   AOI221_X1 U448 (.ZN(n643), 
	.C2(FE_OFN627_n16828), 
	.C1(n16824), 
	.B2(n651), 
	.B1(n16861), 
	.A(n652));
   OAI33_X1 U449 (.ZN(n652), 
	.B3(n655), 
	.B2(n16810), 
	.B1(n654), 
	.A3(n16836), 
	.A2(n16854), 
	.A1(n653));
   OAI222_X1 U450 (.ZN(n635), 
	.C2(n576), 
	.C1(n658), 
	.B2(n610), 
	.B1(n657), 
	.A2(n552), 
	.A1(n656));
   INV_X1 U451 (.ZN(n658), 
	.A(n577));
   NAND3_X1 U452 (.ZN(n577), 
	.A3(n16801), 
	.A2(FE_OFN426_n659), 
	.A1(n16800));
   AOI222_X1 U453 (.ZN(n657), 
	.C2(n661), 
	.C1(n590), 
	.B2(n16836), 
	.B1(n609), 
	.A2(n195), 
	.A1(n660));
   OAI221_X1 U454 (.ZN(n661), 
	.C2(n665), 
	.C1(n664), 
	.B2(n663), 
	.B1(n662), 
	.A(n666));
   NAND2_X1 U455 (.ZN(n665), 
	.A2(FE_OFN629_n16850), 
	.A1(n667));
   NAND2_X1 U456 (.ZN(n663), 
	.A2(FE_OFN79_n16834), 
	.A1(n16680));
   AOI222_X1 U457 (.ZN(n656), 
	.C2(n669), 
	.C1(n16816), 
	.B2(n668), 
	.B1(n17099), 
	.A2(n17098), 
	.A1(n16796));
   OR3_X1 U458 (.ZN(n634), 
	.A3(n672), 
	.A2(n671), 
	.A1(n670));
   OAI33_X1 U459 (.ZN(n672), 
	.B3(FE_OFN429_n673), 
	.B2(n16845), 
	.B1(n514), 
	.A3(FE_OFN95_n16864), 
	.A2(n4956), 
	.A1(n650));
   NOR4_X1 U460 (.ZN(n671), 
	.A4(n459), 
	.A3(n16808), 
	.A2(n674), 
	.A1(n485));
   NOR4_X1 U461 (.ZN(n670), 
	.A4(n677), 
	.A3(n443), 
	.A2(n17098), 
	.A1(n676));
   AOI21_X1 U462 (.ZN(n676), 
	.B2(n504), 
	.B1(n678), 
	.A(n679));
   INV_X1 U463 (.ZN(n678), 
	.A(n680));
   OAI221_X1 U464 (.ZN(n5776), 
	.C2(n17102), 
	.C1(n5255), 
	.B2(n324), 
	.B1(n191), 
	.A(n681));
   AOI21_X1 U465 (.ZN(n681), 
	.B2(vis_pc_o[0]), 
	.B1(n16738), 
	.A(n682));
   NOR4_X1 U466 (.ZN(n682), 
	.A4(n17103), 
	.A3(n684), 
	.A2(n628), 
	.A1(n683));
   INV_X1 U467 (.ZN(n628), 
	.A(n638));
   OAI221_X1 U469 (.ZN(n5777), 
	.C2(FE_OFN667_n17122), 
	.C1(n16833), 
	.B2(FE_PHN675_n17126), 
	.B1(n685), 
	.A(n686));
   NAND3_X1 U470 (.ZN(n686), 
	.A3(n687), 
	.A2(n16851), 
	.A1(n529));
   NOR4_X1 U471 (.ZN(n685), 
	.A4(n691), 
	.A3(n690), 
	.A2(n689), 
	.A1(n688));
   OAI22_X1 U472 (.ZN(n691), 
	.B2(n694), 
	.B1(n5230), 
	.A2(n693), 
	.A1(n692));
   INV_X1 U473 (.ZN(n693), 
	.A(n695));
   OAI33_X1 U474 (.ZN(n690), 
	.B3(n478), 
	.B2(n697), 
	.B1(n677), 
	.A3(n605), 
	.A2(n5165), 
	.A1(n696));
   OAI221_X1 U475 (.ZN(n689), 
	.C2(n699), 
	.C1(FE_OFN95_n16864), 
	.B2(n16808), 
	.B1(n698), 
	.A(n700));
   INV_X1 U476 (.ZN(n700), 
	.A(n701));
   NOR4_X1 U477 (.ZN(n698), 
	.A4(n705), 
	.A3(n704), 
	.A2(n703), 
	.A1(n702));
   AOI21_X1 U478 (.ZN(n705), 
	.B2(n707), 
	.B1(n706), 
	.A(n16807));
   NAND4_X1 U479 (.ZN(n707), 
	.A4(n710), 
	.A3(n709), 
	.A2(n708), 
	.A1(n485));
   NOR3_X1 U480 (.ZN(n710), 
	.A3(n712), 
	.A2(n711), 
	.A1(FE_OFN426_n659));
   INV_X1 U481 (.ZN(n485), 
	.A(n444));
   NAND3_X1 U482 (.ZN(n706), 
	.A3(n629), 
	.A2(n16813), 
	.A1(n475));
   NOR3_X1 U483 (.ZN(n704), 
	.A3(n582), 
	.A2(n580), 
	.A1(n711));
   OAI33_X1 U484 (.ZN(n703), 
	.B3(FE_OFN21_n503), 
	.B2(n716), 
	.B1(n478), 
	.A3(FE_OFN104_n715), 
	.A2(n714), 
	.A1(n713));
   AOI22_X1 U485 (.ZN(n716), 
	.B2(n679), 
	.B1(n718), 
	.A2(n717), 
	.A1(n16814));
   INV_X1 U486 (.ZN(n717), 
	.A(n719));
   AOI211_X1 U487 (.ZN(n719), 
	.C2(n721), 
	.C1(n720), 
	.B(n722), 
	.A(n16804));
   OAI221_X1 U488 (.ZN(n702), 
	.C2(n725), 
	.C1(n724), 
	.B2(n723), 
	.B1(FE_OFN414_n556), 
	.A(n726));
   AOI22_X1 U489 (.ZN(n726), 
	.B2(n730), 
	.B1(n729), 
	.A2(n728), 
	.A1(n727));
   AOI221_X1 U490 (.ZN(n724), 
	.C2(n733), 
	.C1(n732), 
	.B2(n333), 
	.B1(n731), 
	.A(n734));
   INV_X1 U491 (.ZN(n733), 
	.A(n735));
   AOI21_X1 U492 (.ZN(n735), 
	.B2(n505), 
	.B1(n16733), 
	.A(n736));
   NAND4_X1 U493 (.ZN(n688), 
	.A4(n740), 
	.A3(n739), 
	.A2(n738), 
	.A1(n737));
   NOR4_X1 U494 (.ZN(n740), 
	.A4(n545), 
	.A3(n493), 
	.A2(n742), 
	.A1(n741));
   NOR3_X1 U495 (.ZN(n545), 
	.A3(n594), 
	.A2(n16836), 
	.A1(n16828));
   NAND3_X1 U496 (.ZN(n739), 
	.A3(n744), 
	.A2(FE_OFN82_n16856), 
	.A1(n16826));
   OAI21_X1 U497 (.ZN(n744), 
	.B2(n745), 
	.B1(n16820), 
	.A(n640));
   NAND3_X1 U498 (.ZN(n737), 
	.A3(n746), 
	.A2(n16821), 
	.A1(n16824));
   OAI22_X1 U499 (.ZN(n5778), 
	.B2(n748), 
	.B1(n17097), 
	.A2(FE_PHN675_n17126), 
	.A1(n747));
   AOI211_X1 U500 (.ZN(n748), 
	.C2(n16854), 
	.C1(n16680), 
	.B(n534), 
	.A(FE_PHN675_n17126));
   AOI211_X1 U501 (.ZN(n747), 
	.C2(n16821), 
	.C1(n526), 
	.B(n750), 
	.A(n749));
   OAI22_X1 U502 (.ZN(n750), 
	.B2(n696), 
	.B1(n751), 
	.A2(n692), 
	.A1(n499));
   OAI211_X1 U503 (.ZN(n749), 
	.C2(n753), 
	.C1(n752), 
	.B(n755), 
	.A(n754));
   OAI211_X1 U504 (.ZN(n754), 
	.C2(n757), 
	.C1(n756), 
	.B(n16802), 
	.A(FE_OFN21_n503));
   NOR2_X1 U505 (.ZN(n756), 
	.A2(n759), 
	.A1(n758));
   AOI21_X1 U506 (.ZN(n752), 
	.B2(n760), 
	.B1(n543), 
	.A(n761));
   NOR3_X1 U507 (.ZN(n761), 
	.A3(FE_OFN91_n16864), 
	.A2(n16843), 
	.A1(n762));
   OAI22_X1 U508 (.ZN(n5779), 
	.B2(n766), 
	.B1(FE_PHN1586_n5256), 
	.A2(n765), 
	.A1(n764));
   AOI21_X1 U509 (.ZN(n766), 
	.B2(n768), 
	.B1(n767), 
	.A(n765));
   AOI221_X1 U510 (.ZN(n764), 
	.C2(n659), 
	.C1(n770), 
	.B2(n403), 
	.B1(n769), 
	.A(n771));
   OAI22_X1 U511 (.ZN(n771), 
	.B2(n773), 
	.B1(n5243), 
	.A2(n772), 
	.A1(n16816));
   OAI22_X1 U513 (.ZN(n5780), 
	.B2(n775), 
	.B1(n16810), 
	.A2(n765), 
	.A1(n774));
   AOI21_X1 U514 (.ZN(n775), 
	.B2(n776), 
	.B1(n767), 
	.A(n765));
   NOR3_X1 U515 (.ZN(n774), 
	.A3(FE_PHN1501_n779), 
	.A2(n778), 
	.A1(n777));
   INV_X1 U516 (.ZN(n779), 
	.A(n780));
   AOI22_X1 U517 (.ZN(n780), 
	.B2(n769), 
	.B1(n4806), 
	.A2(n770), 
	.A1(n781));
   AOI21_X1 U518 (.ZN(n769), 
	.B2(n783), 
	.B1(n782), 
	.A(n5034));
   NOR2_X1 U519 (.ZN(n783), 
	.A2(n785), 
	.A1(n784));
   OAI33_X1 U520 (.ZN(n778), 
	.B3(n790), 
	.B2(n16816), 
	.B1(n16659), 
	.A3(n788), 
	.A2(n16957), 
	.A1(n786));
   AOI21_X1 U521 (.ZN(n790), 
	.B2(n466), 
	.B1(n791), 
	.A(n792));
   XNOR2_X1 U522 (.ZN(n786), 
	.B(n654), 
	.A(n793));
   NAND2_X1 U523 (.ZN(n654), 
	.A2(n795), 
	.A1(n794));
   NAND2_X1 U524 (.ZN(n793), 
	.A2(FE_OFN15_n16671), 
	.A1(n17097));
   OAI221_X1 U525 (.ZN(n777), 
	.C2(n772), 
	.C1(n16796), 
	.B2(n773), 
	.B1(n16794), 
	.A(n460));
   AOI21_X1 U526 (.ZN(n460), 
	.B2(n798), 
	.B1(n797), 
	.A(n799));
   INV_X1 U527 (.ZN(n773), 
	.A(n800));
   OAI22_X1 U528 (.ZN(n5781), 
	.B2(FE_PHN675_n17126), 
	.B1(n801), 
	.A2(FE_OFN667_n17122), 
	.A1(n16851));
   NOR2_X1 U529 (.ZN(n801), 
	.A2(n803), 
	.A1(n802));
   OAI211_X1 U530 (.ZN(n803), 
	.C2(n16821), 
	.C1(n804), 
	.B(n806), 
	.A(n805));
   AOI22_X1 U531 (.ZN(n806), 
	.B2(n16826), 
	.B1(n809), 
	.A2(FE_OFN450_n808), 
	.A1(n807));
   OAI21_X1 U532 (.ZN(n805), 
	.B2(n811), 
	.B1(n810), 
	.A(n16855));
   OAI33_X1 U533 (.ZN(n811), 
	.B3(n16859), 
	.B2(n812), 
	.B1(n640), 
	.A3(n16843), 
	.A2(FE_OFN627_n16828), 
	.A1(n514));
   AOI21_X1 U534 (.ZN(n810), 
	.B2(n16851), 
	.B1(n5165), 
	.A(n813));
   NOR4_X1 U535 (.ZN(n804), 
	.A4(n817), 
	.A3(n816), 
	.A2(n815), 
	.A1(n814));
   OAI221_X1 U536 (.ZN(n817), 
	.C2(n16813), 
	.C1(n819), 
	.B2(n818), 
	.B1(n499), 
	.A(n820));
   AOI22_X1 U537 (.ZN(n820), 
	.B2(n16659), 
	.B1(n629), 
	.A2(n822), 
	.A1(n821));
   OAI211_X1 U538 (.ZN(n816), 
	.C2(n16659), 
	.C1(n823), 
	.B(n825), 
	.A(n824));
   AOI22_X1 U539 (.ZN(n825), 
	.B2(n827), 
	.B1(n543), 
	.A2(n16871), 
	.A1(n826));
   OAI211_X1 U540 (.ZN(n826), 
	.C2(n625), 
	.C1(n16802), 
	.B(n828), 
	.A(n16680));
   AOI221_X1 U541 (.ZN(n828), 
	.C2(n830), 
	.C1(n16811), 
	.B2(n829), 
	.B1(n821), 
	.A(n831));
   NOR3_X1 U542 (.ZN(n831), 
	.A3(n832), 
	.A2(n16801), 
	.A1(n711));
   OAI22_X1 U543 (.ZN(n830), 
	.B2(n625), 
	.B1(n833), 
	.A2(n582), 
	.A1(n16803));
   NAND3_X1 U544 (.ZN(n829), 
	.A3(n834), 
	.A2(n16657), 
	.A1(n833));
   OAI21_X1 U545 (.ZN(n824), 
	.B2(n731), 
	.B1(n835), 
	.A(n474));
   NOR3_X1 U546 (.ZN(n835), 
	.A3(n16798), 
	.A2(n16796), 
	.A1(n16674));
   AOI221_X1 U547 (.ZN(n823), 
	.C2(n791), 
	.C1(n505), 
	.B2(n16683), 
	.B1(n474), 
	.A(n684));
   INV_X1 U548 (.ZN(n474), 
	.A(n329));
   OAI211_X1 U549 (.ZN(n815), 
	.C2(n610), 
	.C1(n838), 
	.B(n840), 
	.A(n839));
   AOI22_X1 U550 (.ZN(n840), 
	.B2(n597), 
	.B1(n842), 
	.A2(n473), 
	.A1(n841));
   AOI21_X1 U551 (.ZN(n842), 
	.B2(n606), 
	.B1(n16843), 
	.A(n16838));
   AOI21_X1 U552 (.ZN(n841), 
	.B2(n832), 
	.B1(n843), 
	.A(n16814));
   NAND3_X1 U553 (.ZN(n839), 
	.A3(n730), 
	.A2(FE_OFN608_n16686), 
	.A1(n16816));
   AOI21_X1 U554 (.ZN(n838), 
	.B2(n632), 
	.B1(n844), 
	.A(n845));
   NOR3_X1 U555 (.ZN(n845), 
	.A3(n617), 
	.A2(FE_OFN107_n585), 
	.A1(n846));
   OR4_X1 U556 (.ZN(n814), 
	.A4(n848), 
	.A3(n482), 
	.A2(n484), 
	.A1(n847));
   NOR3_X1 U557 (.ZN(n847), 
	.A3(n567), 
	.A2(n16871), 
	.A1(n849));
   OAI211_X1 U558 (.ZN(n802), 
	.C2(n851), 
	.C1(n850), 
	.B(n853), 
	.A(n852));
   NOR3_X1 U559 (.ZN(n853), 
	.A3(n856), 
	.A2(n855), 
	.A1(n854));
   NOR3_X1 U560 (.ZN(n856), 
	.A3(n857), 
	.A2(FE_OFN104_n715), 
	.A1(n664));
   NOR3_X1 U561 (.ZN(n854), 
	.A3(n849), 
	.A2(n604), 
	.A1(FE_OFN425_n650));
   OAI21_X1 U562 (.ZN(n852), 
	.B2(n807), 
	.B1(n858), 
	.A(n16862));
   NOR3_X1 U563 (.ZN(n858), 
	.A3(n860), 
	.A2(n16820), 
	.A1(n859));
   AOI21_X1 U564 (.ZN(n850), 
	.B2(n861), 
	.B1(n597), 
	.A(n599));
   NOR3_X1 U565 (.ZN(n599), 
	.A3(n16847), 
	.A2(FE_OFN70_n16867), 
	.A1(n16680));
   OAI21_X1 U566 (.ZN(n861), 
	.B2(n16843), 
	.B1(FE_OFN627_n16828), 
	.A(n863));
   OAI221_X1 U567 (.ZN(n5782), 
	.C2(n324), 
	.C1(n4948), 
	.B2(n16792), 
	.B1(n5006), 
	.A(n865));
   AOI22_X1 U568 (.ZN(n865), 
	.B2(n867), 
	.B1(n866), 
	.A2(FE_OFN118_HADDR_31_), 
	.A1(n17104));
   INV_X1 U569 (.ZN(n5783), 
	.A(n868));
   AOI221_X1 U570 (.ZN(n868), 
	.C2(n866), 
	.C1(n869), 
	.B2(n17104), 
	.B1(haddr_o[9]), 
	.A(n870));
   OAI22_X1 U571 (.ZN(n870), 
	.B2(n5546), 
	.B1(n324), 
	.A2(n4814), 
	.A1(n16792));
   AOI22_X1 U573 (.ZN(n872), 
	.B2(vis_ipsr_o[3]), 
	.B1(n322), 
	.A2(vis_pc_o[2]), 
	.A1(n16738));
   INV_X1 U574 (.ZN(n871), 
	.A(haddr_o[3]));
   INV_X1 U575 (.ZN(n5785), 
	.A(n873));
   AOI221_X1 U576 (.ZN(n873), 
	.C2(n866), 
	.C1(n874), 
	.B2(n17104), 
	.B1(FE_OFN112_HADDR_30_), 
	.A(n875));
   OAI22_X1 U577 (.ZN(n875), 
	.B2(n4954), 
	.B1(n324), 
	.A2(n4817), 
	.A1(n16792));
   AOI22_X1 U579 (.ZN(n877), 
	.B2(vis_ipsr_o[2]), 
	.B1(n322), 
	.A2(vis_pc_o[1]), 
	.A1(n16738));
   OAI221_X1 U580 (.ZN(n5787), 
	.C2(n17102), 
	.C1(n5626), 
	.B2(n17103), 
	.B1(n878), 
	.A(n879));
   AOI22_X1 U581 (.ZN(n879), 
	.B2(vis_apsr_o[0]), 
	.B1(n322), 
	.A2(FE_PHN1320_SYNOPSYS_UNCONNECTED_518), 
	.A1(n16738));
   OAI221_X1 U583 (.ZN(n5788), 
	.C2(n324), 
	.C1(n4953), 
	.B2(n16792), 
	.B1(n5239), 
	.A(n880));
   AOI22_X1 U584 (.ZN(n880), 
	.B2(n881), 
	.B1(n866), 
	.A2(FE_OFN115_HADDR_29_), 
	.A1(n17104));
   OAI221_X1 U585 (.ZN(n5789), 
	.C2(n17122), 
	.C1(n16862), 
	.B2(FE_PHN675_n17126), 
	.B1(n882), 
	.A(n883));
   NAND3_X1 U586 (.ZN(n883), 
	.A3(n884), 
	.A2(n592), 
	.A1(n4974));
   NOR4_X1 U587 (.ZN(n882), 
	.A4(n888), 
	.A3(n887), 
	.A2(n886), 
	.A1(n885));
   OAI33_X1 U588 (.ZN(n888), 
	.B3(FE_OFN21_n503), 
	.B2(n16847), 
	.B1(n889), 
	.A3(n532), 
	.A2(n851), 
	.A1(n653));
   NAND2_X1 U589 (.ZN(n889), 
	.A2(n483), 
	.A1(n631));
   NOR3_X1 U590 (.ZN(n887), 
	.A3(FE_OFN104_n715), 
	.A2(n714), 
	.A1(n650));
   NAND4_X1 U591 (.ZN(n886), 
	.A4(n892), 
	.A3(n891), 
	.A2(n618), 
	.A1(FE_OFN461_n890));
   NAND3_X1 U592 (.ZN(n885), 
	.A3(n895), 
	.A2(n894), 
	.A1(n893));
   AOI221_X1 U593 (.ZN(n895), 
	.C2(n799), 
	.C1(n649), 
	.B2(n728), 
	.B1(n809), 
	.A(n896));
   AOI22_X1 U594 (.ZN(n894), 
	.B2(FE_OFN95_n16864), 
	.B1(n899), 
	.A2(n898), 
	.A1(n897));
   OAI21_X1 U595 (.ZN(n899), 
	.B2(n900), 
	.B1(n813), 
	.A(n522));
   NAND2_X1 U596 (.ZN(n900), 
	.A2(n610), 
	.A1(n16838));
   OAI22_X1 U597 (.ZN(n898), 
	.B2(n901), 
	.B1(n846), 
	.A2(n673), 
	.A1(n762));
   NAND2_X1 U598 (.ZN(n901), 
	.A2(FE_OFN82_n16856), 
	.A1(n632));
   AOI22_X1 U599 (.ZN(n893), 
	.B2(n903), 
	.B1(n16820), 
	.A2(n902), 
	.A1(n466));
   NAND4_X1 U600 (.ZN(n903), 
	.A4(n907), 
	.A3(n906), 
	.A2(n905), 
	.A1(n904));
   NOR3_X1 U601 (.ZN(n907), 
	.A3(n910), 
	.A2(n909), 
	.A1(n908));
   NOR3_X1 U602 (.ZN(n910), 
	.A3(n859), 
	.A2(FE_OFN104_n715), 
	.A1(n911));
   OAI33_X1 U603 (.ZN(n908), 
	.B3(FE_OFN634_n16871), 
	.B2(n16833), 
	.B1(n912), 
	.A3(n651), 
	.A2(n16854), 
	.A1(n694));
   AOI222_X1 U604 (.ZN(n906), 
	.C2(n916), 
	.C1(n597), 
	.B2(n915), 
	.B1(n914), 
	.A2(n913), 
	.A1(n708));
   OAI21_X1 U605 (.ZN(n916), 
	.B2(n918), 
	.B1(n917), 
	.A(n919));
   OAI21_X1 U606 (.ZN(n915), 
	.B2(n653), 
	.B1(n714), 
	.A(FE_OFN72_n16867));
   OAI22_X1 U607 (.ZN(n913), 
	.B2(n921), 
	.B1(n16807), 
	.A2(n920), 
	.A1(n16795));
   AOI22_X1 U608 (.ZN(n921), 
	.B2(n17098), 
	.B1(n923), 
	.A2(n922), 
	.A1(n5243));
   AOI221_X1 U609 (.ZN(n920), 
	.C2(n16816), 
	.C1(n721), 
	.B2(n16733), 
	.B1(n720), 
	.A(n924));
   XOR2_X1 U610 (.Z(n924), 
	.B(n731), 
	.A(n17098));
   AOI221_X1 U611 (.ZN(n905), 
	.C2(n926), 
	.C1(n483), 
	.B2(n925), 
	.B1(n4974), 
	.A(n927));
   AOI21_X1 U612 (.ZN(n927), 
	.B2(n16816), 
	.B1(n928), 
	.A(n580));
   XOR2_X1 U613 (.Z(n928), 
	.B(n16796), 
	.A(n16798));
   OAI211_X1 U614 (.ZN(n926), 
	.C2(n711), 
	.C1(n16847), 
	.B(n16854), 
	.A(n929));
   NAND3_X1 U615 (.ZN(n929), 
	.A3(n16862), 
	.A2(n596), 
	.A1(n930));
   OAI221_X1 U616 (.ZN(n925), 
	.C2(n582), 
	.C1(n932), 
	.B2(n931), 
	.B1(n819), 
	.A(n933));
   AOI21_X1 U617 (.ZN(n933), 
	.B2(n935), 
	.B1(n934), 
	.A(n494));
   INV_X1 U618 (.ZN(n494), 
	.A(n627));
   NAND2_X1 U619 (.ZN(n627), 
	.A2(FE_OFN625_n16814), 
	.A1(n936));
   OAI211_X1 U620 (.ZN(n935), 
	.C2(n16657), 
	.C1(n16800), 
	.B(n938), 
	.A(n937));
   AOI221_X1 U621 (.ZN(n938), 
	.C2(n16817), 
	.C1(n668), 
	.B2(n16816), 
	.B1(n721), 
	.A(n939));
   XOR2_X1 U622 (.Z(n937), 
	.B(n469), 
	.A(n17098));
   AOI222_X1 U623 (.ZN(n904), 
	.C2(n482), 
	.C1(n16797), 
	.B2(n475), 
	.B1(n684), 
	.A2(n16659), 
	.A1(n934));
   INV_X1 U624 (.ZN(n684), 
	.A(n940));
   NAND4_X1 U625 (.ZN(n902), 
	.A4(n942), 
	.A3(n512), 
	.A2(n819), 
	.A1(n941));
   AOI221_X1 U626 (.ZN(n942), 
	.C2(n16734), 
	.C1(n943), 
	.B2(n16683), 
	.B1(FE_OFN456_n822), 
	.A(n944));
   NOR3_X1 U627 (.ZN(n944), 
	.A3(n16659), 
	.A2(n16862), 
	.A1(n945));
   OAI221_X1 U628 (.ZN(n5790), 
	.C2(n17122), 
	.C1(n5502), 
	.B2(n946), 
	.B1(haddr_o[4]), 
	.A(n255));
   OAI221_X1 U629 (.ZN(n5791), 
	.C2(n17122), 
	.C1(FE_PHN1894_n5149), 
	.B2(n946), 
	.B1(n947), 
	.A(n255));
   XOR2_X1 U630 (.Z(n947), 
	.B(n948), 
	.A(haddr_o[3]));
   OAI211_X1 U631 (.ZN(n5792), 
	.C2(n17122), 
	.C1(n5096), 
	.B(n255), 
	.A(n949));
   OAI21_X1 U632 (.ZN(n949), 
	.B2(haddr_o[3]), 
	.B1(haddr_o[5]), 
	.A(n256));
   OAI221_X1 U633 (.ZN(n5793), 
	.C2(n17122), 
	.C1(n5017), 
	.B2(n946), 
	.B1(haddr_o[8]), 
	.A(n255));
   OAI21_X1 U634 (.ZN(n255), 
	.B2(n951), 
	.B1(n950), 
	.A(n256));
   NAND4_X1 U635 (.ZN(n951), 
	.A4(n954), 
	.A3(n953), 
	.A2(n952), 
	.A1(haddr_o[15]));
   NOR4_X1 U636 (.ZN(n954), 
	.A4(n958), 
	.A3(n957), 
	.A2(n956), 
	.A1(n955));
   AOI22_X1 U637 (.ZN(n958), 
	.B2(n962), 
	.B1(n961), 
	.A2(n960), 
	.A1(n959));
   NOR4_X1 U638 (.ZN(n962), 
	.A4(haddr_o[5]), 
	.A3(haddr_o[6]), 
	.A2(haddr_o[7]), 
	.A1(haddr_o[9]));
   AOI221_X1 U639 (.ZN(n961), 
	.C2(haddr_o[11]), 
	.C1(n964), 
	.B2(n963), 
	.B1(haddr_o[8]), 
	.A(n965));
   NOR3_X1 U640 (.ZN(n965), 
	.A3(haddr_o[3]), 
	.A2(haddr_o[4]), 
	.A1(haddr_o[10]));
   NAND3_X1 U641 (.ZN(n964), 
	.A3(haddr_o[10]), 
	.A2(haddr_o[2]), 
	.A1(haddr_o[8]));
   NOR3_X1 U642 (.ZN(n960), 
	.A3(haddr_o[3]), 
	.A2(haddr_o[6]), 
	.A1(n966));
   AOI21_X1 U643 (.ZN(n966), 
	.B2(n967), 
	.B1(n876), 
	.A(n968));
   AOI21_X1 U644 (.ZN(n959), 
	.B2(n970), 
	.B1(n969), 
	.A(n971));
   XNOR2_X1 U645 (.ZN(n971), 
	.B(haddr_o[8]), 
	.A(haddr_o[9]));
   NAND4_X1 U646 (.ZN(n970), 
	.A4(n972), 
	.A3(n876), 
	.A2(n968), 
	.A1(n967));
   NOR2_X1 U647 (.ZN(n972), 
	.A2(haddr_o[11]), 
	.A1(haddr_o[10]));
   NOR3_X1 U649 (.ZN(n953), 
	.A3(haddr_o[17]), 
	.A2(haddr_o[18]), 
	.A1(haddr_o[16]));
   NAND4_X1 U650 (.ZN(n950), 
	.A4(n975), 
	.A3(n974), 
	.A2(n317), 
	.A1(n973));
   NOR4_X1 U651 (.ZN(n975), 
	.A4(haddr_o[19]), 
	.A3(haddr_o[20]), 
	.A2(haddr_o[21]), 
	.A1(haddr_o[22]));
   NOR3_X1 U652 (.ZN(n974), 
	.A3(haddr_o[26]), 
	.A2(haddr_o[27]), 
	.A1(haddr_o[25]));
   NAND2_X1 U653 (.ZN(n5794), 
	.A2(n977), 
	.A1(n976));
   NAND3_X1 U654 (.ZN(n977), 
	.A3(n980), 
	.A2(n979), 
	.A1(n978));
   OAI21_X1 U655 (.ZN(n976), 
	.B2(n16808), 
	.B1(1'b0), 
	.A(FE_PHN674_n17127));
   OAI22_X1 U665 (.ZN(n5795), 
	.B2(n999), 
	.B1(FE_PHN674_n17127), 
	.A2(n17122), 
	.A1(n5231));
   OAI21_X1 U666 (.ZN(n5796), 
	.B2(n431), 
	.B1(n430), 
	.A(FE_PHN2045_n1000));
   NAND4_X1 U667 (.ZN(n1000), 
	.A4(n1002), 
	.A3(n334), 
	.A2(n1001), 
	.A1(n430));
   OAI21_X1 U668 (.ZN(n5797), 
	.B2(n1003), 
	.B1(n5233), 
	.A(n1004));
   NAND2_X1 U669 (.ZN(n5798), 
	.A2(n1006), 
	.A1(n1005));
   OAI211_X1 U670 (.ZN(n1006), 
	.C2(n1007), 
	.C1(n189), 
	.B(n17124), 
	.A(n1008));
   OAI21_X1 U671 (.ZN(n1005), 
	.B2(n42), 
	.B1(n189), 
	.A(n1009));
   INV_X4 U672 (.ZN(n42), 
	.A(n37));
   INV_X1 U673 (.ZN(n189), 
	.A(n1010));
   OAI21_X1 U674 (.ZN(n5799), 
	.B2(n1011), 
	.B1(n5229), 
	.A(n1012));
   NOR3_X1 U675 (.ZN(n1011), 
	.A3(n181), 
	.A2(n186), 
	.A1(n200));
   OAI22_X1 U676 (.ZN(n5800), 
	.B2(FE_PHN675_n17126), 
	.B1(n1013), 
	.A2(n17122), 
	.A1(n4947));
   NOR4_X1 U677 (.ZN(n1013), 
	.A4(n1017), 
	.A3(n1016), 
	.A2(n1015), 
	.A1(n1014));
   OAI33_X1 U678 (.ZN(n1017), 
	.B3(n1020), 
	.B2(n16795), 
	.B1(n1019), 
	.A3(n552), 
	.A2(n1018), 
	.A1(n843));
   NOR2_X1 U679 (.ZN(n1020), 
	.A2(n1021), 
	.A1(n16812));
   AOI21_X1 U680 (.ZN(n1018), 
	.B2(n16798), 
	.B1(n1022), 
	.A(n922));
   INV_X1 U681 (.ZN(n922), 
	.A(n712));
   NOR3_X1 U682 (.ZN(n1016), 
	.A3(n1023), 
	.A2(FE_OFN85_n16839), 
	.A1(n699));
   NAND3_X1 U683 (.ZN(n1015), 
	.A3(n1026), 
	.A2(n1025), 
	.A1(n1024));
   OAI211_X1 U684 (.ZN(n1026), 
	.C2(n465), 
	.C1(n333), 
	.B(n574), 
	.A(n16804));
   OAI211_X1 U685 (.ZN(n1014), 
	.C2(n514), 
	.C1(n1027), 
	.B(n1029), 
	.A(n1028));
   AOI222_X1 U686 (.ZN(n1029), 
	.C2(n1032), 
	.C1(n728), 
	.B2(n1031), 
	.B1(n991), 
	.A2(n1030), 
	.A1(n563));
   OAI22_X1 U687 (.ZN(n1032), 
	.B2(n1033), 
	.B1(n808), 
	.A2(n650), 
	.A1(FE_OFN627_n16828));
   NAND2_X1 U688 (.ZN(n1033), 
	.A2(FE_OFN469_n1034), 
	.A1(n528));
   OAI21_X1 U689 (.ZN(n1031), 
	.B2(n1035), 
	.B1(n994), 
	.A(n646));
   OAI221_X1 U690 (.ZN(n1030), 
	.C2(n692), 
	.C1(FE_OFN411_n499), 
	.B2(n699), 
	.B1(n610), 
	.A(n1036));
   INV_X1 U691 (.ZN(n1036), 
	.A(n1037));
   OAI22_X1 U692 (.ZN(n5823), 
	.B2(n1038), 
	.B1(n422), 
	.A2(n193), 
	.A1(n16820));
   OAI21_X1 U693 (.ZN(n1038), 
	.B2(n1040), 
	.B1(n1039), 
	.A(n17122));
   NOR2_X1 U694 (.ZN(n1039), 
	.A2(n1042), 
	.A1(n1041));
   AOI21_X1 U695 (.ZN(n193), 
	.B2(n641), 
	.B1(n1043), 
	.A(n196));
   OAI22_X1 U696 (.ZN(n5824), 
	.B2(n1047), 
	.B1(n1046), 
	.A2(n1045), 
	.A1(n1044));
   INV_X1 U697 (.ZN(n1046), 
	.A(n1048));
   INV_X1 U698 (.ZN(n1044), 
	.A(n1047));
   NAND2_X1 U699 (.ZN(n1047), 
	.A2(n1049), 
	.A1(n17124));
   OAI21_X1 U700 (.ZN(n5825), 
	.B2(n930), 
	.B1(n1050), 
	.A(FE_PHN2042_n1051));
   OAI21_X1 U701 (.ZN(n1051), 
	.B2(n200), 
	.B1(n1052), 
	.A(n1053));
   OAI21_X1 U702 (.ZN(n5826), 
	.B2(n1054), 
	.B1(n5234), 
	.A(n1055));
   OAI211_X1 U703 (.ZN(n1055), 
	.C2(n1057), 
	.C1(n1056), 
	.B(n5167), 
	.A(n16808));
   NOR3_X1 U704 (.ZN(n1057), 
	.A3(n196), 
	.A2(FE_OFN75_n16806), 
	.A1(vis_pc_o[1]));
   NAND2_X1 U705 (.ZN(n196), 
	.A2(n1058), 
	.A1(n17124));
   NOR4_X1 U706 (.ZN(n1056), 
	.A4(n1058), 
	.A3(n1059), 
	.A2(n181), 
	.A1(n186));
   OAI22_X1 U707 (.ZN(n5827), 
	.B2(n1060), 
	.B1(n1059), 
	.A2(n184), 
	.A1(n1054));
   OAI21_X1 U708 (.ZN(n1060), 
	.B2(n1062), 
	.B1(n1061), 
	.A(n16808));
   NOR2_X1 U709 (.ZN(n1062), 
	.A2(n5228), 
	.A1(n5167));
   NOR3_X1 U710 (.ZN(n1061), 
	.A3(n1058), 
	.A2(n183), 
	.A1(FE_OFN19_n1063));
   OAI22_X1 U712 (.ZN(n5828), 
	.B2(FE_PHN675_n17126), 
	.B1(n1064), 
	.A2(n17122), 
	.A1(n5230));
   AOI22_X1 U713 (.ZN(n1064), 
	.B2(n1066), 
	.B1(n183), 
	.A2(n181), 
	.A1(n1065));
   OAI21_X1 U714 (.ZN(n1065), 
	.B2(n1068), 
	.B1(n1067), 
	.A(n5229));
   INV_X1 U715 (.ZN(n1068), 
	.A(n1069));
   OAI22_X1 U716 (.ZN(n4854), 
	.B2(n1071), 
	.B1(n4826), 
	.A2(n1070), 
	.A1(n19));
   OAI22_X1 U717 (.ZN(n4855), 
	.B2(n17095), 
	.B1(FE_PHN2140_n5515), 
	.A2(n16781), 
	.A1(n19));
   OAI22_X1 U718 (.ZN(n4856), 
	.B2(n17095), 
	.B1(FE_PHN2429_n5505), 
	.A2(n17094), 
	.A1(n247));
   OAI22_X1 U719 (.ZN(n4857), 
	.B2(n17095), 
	.B1(FE_PHN2430_n5520), 
	.A2(n17094), 
	.A1(n229));
   OAI22_X1 U720 (.ZN(n4858), 
	.B2(n17095), 
	.B1(FE_PHN2106_n5506), 
	.A2(n16781), 
	.A1(n245));
   OAI22_X1 U721 (.ZN(n4859), 
	.B2(n17095), 
	.B1(FE_PHN2180_n5517), 
	.A2(n16781), 
	.A1(n226));
   OAI22_X1 U722 (.ZN(n4860), 
	.B2(n1075), 
	.B1(n249), 
	.A2(n1074), 
	.A1(FE_PHN3501_n5516));
   OAI22_X1 U723 (.ZN(n4861), 
	.B2(n17095), 
	.B1(FE_PHN3512_n5510), 
	.A2(n17094), 
	.A1(n249));
   OAI22_X1 U724 (.ZN(n4862), 
	.B2(n1078), 
	.B1(n1077), 
	.A2(n1076), 
	.A1(n5503));
   OAI22_X1 U725 (.ZN(n4863), 
	.B2(n1080), 
	.B1(n221), 
	.A2(n1079), 
	.A1(FE_PHN4850_n5168));
   OAI22_X1 U726 (.ZN(n4864), 
	.B2(n1080), 
	.B1(n215), 
	.A2(n1079), 
	.A1(FE_PHN3602_n4829));
   OAI22_X1 U727 (.ZN(n4865), 
	.B2(n17095), 
	.B1(FE_PHN2428_n5507), 
	.A2(n16781), 
	.A1(n240));
   OAI22_X1 U728 (.ZN(n4866), 
	.B2(n17095), 
	.B1(FE_PHN2223_n5508), 
	.A2(n16781), 
	.A1(n236));
   OAI22_X1 U729 (.ZN(n4867), 
	.B2(n17095), 
	.B1(FE_PHN2302_n5509), 
	.A2(n16781), 
	.A1(n221));
   OAI22_X1 U730 (.ZN(n4868), 
	.B2(n17095), 
	.B1(FE_PHN2232_n5511), 
	.A2(n16781), 
	.A1(n210));
   OAI22_X1 U731 (.ZN(n4869), 
	.B2(n17095), 
	.B1(FE_PHN2412_n5512), 
	.A2(n16781), 
	.A1(n215));
   OAI22_X1 U732 (.ZN(n4870), 
	.B2(n17095), 
	.B1(FE_PHN2347_n5513), 
	.A2(n16781), 
	.A1(n218));
   OAI22_X1 U733 (.ZN(n4871), 
	.B2(n17095), 
	.B1(FE_PHN2240_n5514), 
	.A2(n16781), 
	.A1(n224));
   OAI22_X1 U734 (.ZN(n4872), 
	.B2(n17095), 
	.B1(FE_PHN2376_n5571), 
	.A2(n17094), 
	.A1(n238));
   OAI22_X1 U735 (.ZN(n4873), 
	.B2(n17095), 
	.B1(FE_PHN2333_n5600), 
	.A2(n17094), 
	.A1(n242));
   OAI22_X1 U736 (.ZN(n4874), 
	.B2(n1075), 
	.B1(n210), 
	.A2(n1074), 
	.A1(n4833));
   INV_X1 U737 (.ZN(n1075), 
	.A(n1074));
   NOR3_X1 U738 (.ZN(n1074), 
	.A3(n261), 
	.A2(FE_PHN1037_n5007), 
	.A1(n251));
   OAI21_X1 U739 (.ZN(n4875), 
	.B2(n17122), 
	.B1(n4834), 
	.A(n1081));
   NAND4_X1 U740 (.ZN(n1081), 
	.A4(n1084), 
	.A3(n1083), 
	.A2(n422), 
	.A1(n1082));
   AOI221_X1 U741 (.ZN(n1084), 
	.C2(n1087), 
	.C1(FE_OFN100_n1086), 
	.B2(n651), 
	.B1(n1085), 
	.A(FE_PHN675_n17126));
   OAI22_X1 U743 (.ZN(n1085), 
	.B2(n16826), 
	.B1(n1088), 
	.A2(n696), 
	.A1(n16854));
   INV_X1 U744 (.ZN(n1083), 
	.A(n1089));
   AOI21_X1 U745 (.ZN(n1089), 
	.B2(n1090), 
	.B1(n590), 
	.A(n1091));
   AOI221_X1 U746 (.ZN(n1091), 
	.C2(n1087), 
	.C1(n1093), 
	.B2(n1092), 
	.B1(FE_OFN95_n16864), 
	.A(n1094));
   NAND3_X1 U747 (.ZN(n1082), 
	.A3(n1097), 
	.A2(n1096), 
	.A1(n1095));
   OAI22_X1 U748 (.ZN(n4876), 
	.B2(n687), 
	.B1(n5165), 
	.A2(n1059), 
	.A1(n5829));
   OAI21_X1 U749 (.ZN(n5829), 
	.B2(n1099), 
	.B1(n1098), 
	.A(n194));
   NAND4_X1 U750 (.ZN(n1099), 
	.A4(n2), 
	.A3(n9), 
	.A2(n8), 
	.A1(n7));
   NAND4_X1 U755 (.ZN(n1098), 
	.A4(n6), 
	.A3(n5), 
	.A2(n4), 
	.A1(n3));
   OAI21_X1 U760 (.ZN(n4878), 
	.B2(n17122), 
	.B1(n4843), 
	.A(n1100));
   OAI21_X1 U761 (.ZN(n1100), 
	.B2(n1102), 
	.B1(n1101), 
	.A(n17122));
   NOR3_X1 U762 (.ZN(n1102), 
	.A3(FE_OFN98_n1104), 
	.A2(n16821), 
	.A1(n1103));
   NOR4_X1 U763 (.ZN(n1101), 
	.A4(n568), 
	.A3(n616), 
	.A2(n556), 
	.A1(n532));
   OAI21_X1 U764 (.ZN(n4879), 
	.B2(n17122), 
	.B1(n4845), 
	.A(n1105));
   OAI211_X1 U765 (.ZN(n1105), 
	.C2(n1009), 
	.C1(n1106), 
	.B(n17124), 
	.A(n1107));
   OAI22_X1 U766 (.ZN(n4880), 
	.B2(n687), 
	.B1(n5228), 
	.A2(n1059), 
	.A1(n181));
   OAI22_X1 U767 (.ZN(n4881), 
	.B2(n1109), 
	.B1(FE_PHN3103_n4847), 
	.A2(FE_PHN776_n1108), 
	.A1(n373));
   OAI22_X1 U768 (.ZN(n4882), 
	.B2(n1080), 
	.B1(n210), 
	.A2(n1079), 
	.A1(FE_PHN5123_n4848));
   INV_X1 U769 (.ZN(n1079), 
	.A(n1080));
   NAND3_X1 U770 (.ZN(n1080), 
	.A3(n1111), 
	.A2(n253), 
	.A1(n1110));
   OAI22_X1 U771 (.ZN(n4883), 
	.B2(n1071), 
	.B1(FE_PHN2826_n5097), 
	.A2(n1070), 
	.A1(n1077));
   OAI22_X1 U772 (.ZN(n4884), 
	.B2(n17095), 
	.B1(FE_PHN2426_n5581), 
	.A2(n17094), 
	.A1(n232));
   OAI22_X1 U773 (.ZN(n4885), 
	.B2(n17095), 
	.B1(FE_PHN2364_n5639), 
	.A2(n17094), 
	.A1(n1112));
   OAI22_X1 U774 (.ZN(n4886), 
	.B2(FE_PHN675_n17126), 
	.B1(n1113), 
	.A2(n17122), 
	.A1(n5167));
   OAI22_X1 U775 (.ZN(n4887), 
	.B2(n17095), 
	.B1(FE_PHN2245_n5033), 
	.A2(n17094), 
	.A1(n1114));
   OAI22_X1 U776 (.ZN(n4888), 
	.B2(n17095), 
	.B1(FE_PHN2270_n5067), 
	.A2(n17094), 
	.A1(n1115));
   OAI22_X1 U777 (.ZN(n4889), 
	.B2(n17095), 
	.B1(FE_PHN2330_n5579), 
	.A2(n17094), 
	.A1(n234));
   OAI22_X1 U778 (.ZN(n4890), 
	.B2(n17095), 
	.B1(FE_PHN2385_n5625), 
	.A2(n17094), 
	.A1(n1116));
   OAI22_X1 U779 (.ZN(n4891), 
	.B2(n17095), 
	.B1(FE_PHN2378_n5618), 
	.A2(n17094), 
	.A1(n1117));
   OAI22_X1 U780 (.ZN(n4892), 
	.B2(n17095), 
	.B1(FE_PHN2254_n5074), 
	.A2(n17094), 
	.A1(n1118));
   AOI21_X1 U781 (.ZN(n4902), 
	.B2(n1120), 
	.B1(n17092), 
	.A(n1121));
   AOI21_X1 U782 (.ZN(n4903), 
	.B2(n1122), 
	.B1(n17092), 
	.A(n1123));
   AOI221_X1 U783 (.ZN(n4904), 
	.C2(n1126), 
	.C1(n1125), 
	.B2(hwdata_o[9]), 
	.B1(n1124), 
	.A(FE_PHN1665_n1127));
   OAI21_X1 U784 (.ZN(n1127), 
	.B2(n1129), 
	.B1(n1128), 
	.A(FE_PHN4637_IRQ_9_));
   OAI22_X1 U786 (.ZN(n4906), 
	.B2(n1131), 
	.B1(FE_PHN4697_n1130), 
	.A2(n1109), 
	.A1(n4777));
   INV_X1 U787 (.ZN(n1130), 
	.A(hrdata_i[16]));
   OAI22_X1 U788 (.ZN(n4907), 
	.B2(n1131), 
	.B1(FE_PHN4699_n1132), 
	.A2(n1109), 
	.A1(n4778));
   INV_X1 U789 (.ZN(n1132), 
	.A(hrdata_i[17]));
   OAI22_X1 U790 (.ZN(n4908), 
	.B2(n1131), 
	.B1(FE_PHN4698_n1133), 
	.A2(n1109), 
	.A1(n4779));
   INV_X1 U791 (.ZN(n1133), 
	.A(hrdata_i[18]));
   OAI22_X1 U792 (.ZN(n4909), 
	.B2(n1131), 
	.B1(FE_PHN5207_n1134), 
	.A2(n1109), 
	.A1(n4780));
   INV_X1 U793 (.ZN(n1134), 
	.A(hrdata_i[19]));
   OAI22_X1 U794 (.ZN(n4910), 
	.B2(n1131), 
	.B1(FE_PHN4722_n1135), 
	.A2(n1109), 
	.A1(n4781));
   INV_X1 U795 (.ZN(n1135), 
	.A(hrdata_i[20]));
   OAI22_X1 U796 (.ZN(n4911), 
	.B2(n1131), 
	.B1(FE_PHN4724_n1136), 
	.A2(n1109), 
	.A1(n4782));
   INV_X1 U797 (.ZN(n1136), 
	.A(hrdata_i[21]));
   OAI22_X1 U798 (.ZN(n4912), 
	.B2(n1131), 
	.B1(FE_PHN5206_n1137), 
	.A2(n1109), 
	.A1(n4783));
   INV_X1 U799 (.ZN(n1137), 
	.A(hrdata_i[22]));
   OAI22_X1 U800 (.ZN(n4913), 
	.B2(n1131), 
	.B1(FE_PHN4720_n1138), 
	.A2(n1109), 
	.A1(n4784));
   INV_X1 U801 (.ZN(n1138), 
	.A(hrdata_i[23]));
   OAI22_X1 U802 (.ZN(n4914), 
	.B2(n1131), 
	.B1(FE_PHN4696_n1139), 
	.A2(n1109), 
	.A1(n4785));
   INV_X1 U803 (.ZN(n1139), 
	.A(hrdata_i[24]));
   OAI22_X1 U804 (.ZN(n4915), 
	.B2(n1131), 
	.B1(FE_PHN763_n1140), 
	.A2(n1109), 
	.A1(n4786));
   OAI22_X1 U805 (.ZN(n4916), 
	.B2(n1131), 
	.B1(FE_PHN4721_n1141), 
	.A2(n1109), 
	.A1(n4787));
   INV_X1 U806 (.ZN(n1141), 
	.A(hrdata_i[26]));
   OAI22_X1 U807 (.ZN(n4917), 
	.B2(n1131), 
	.B1(FE_PHN755_n1142), 
	.A2(n1109), 
	.A1(n4788));
   OAI22_X1 U808 (.ZN(n4918), 
	.B2(n1131), 
	.B1(FE_PHN806_n1143), 
	.A2(n1109), 
	.A1(n4789));
   OAI22_X1 U809 (.ZN(n4919), 
	.B2(n1131), 
	.B1(FE_PHN765_n1144), 
	.A2(n1109), 
	.A1(n4790));
   OAI22_X1 U810 (.ZN(n4920), 
	.B2(n1131), 
	.B1(FE_PHN2928_n1145), 
	.A2(n1109), 
	.A1(n4791));
   OAI22_X1 U811 (.ZN(n4921), 
	.B2(n1131), 
	.B1(FE_PHN4702_n1146), 
	.A2(n1109), 
	.A1(n4792));
   INV_X1 U813 (.ZN(n1146), 
	.A(hrdata_i[31]));
   OAI222_X1 U816 (.ZN(n4925), 
	.C2(n17102), 
	.C1(n4762), 
	.B2(n16792), 
	.B1(n4820), 
	.A2(n17103), 
	.A1(n1149));
   INV_X1 U818 (.ZN(n4927), 
	.A(n1151));
   AOI222_X1 U819 (.ZN(n1151), 
	.C2(n866), 
	.C1(n1152), 
	.B2(n16738), 
	.B1(FE_PHN1339_SYNOPSYS_UNCONNECTED_540), 
	.A2(n17104), 
	.A1(haddr_o[6]));
   OAI222_X1 U821 (.ZN(n4928), 
	.C2(n17102), 
	.C1(n4764), 
	.B2(n16792), 
	.B1(FE_PHN3098_n5238), 
	.A2(n318), 
	.A1(n1153));
   OAI222_X1 U822 (.ZN(n4929), 
	.C2(n17102), 
	.C1(n4765), 
	.B2(n16792), 
	.B1(FE_PHN3100_n5573), 
	.A2(n318), 
	.A1(n1154));
   OAI222_X1 U823 (.ZN(n4930), 
	.C2(n17102), 
	.C1(n4766), 
	.B2(n16792), 
	.B1(FE_PHN3099_n5601), 
	.A2(n318), 
	.A1(n1155));
   OAI222_X1 U824 (.ZN(n4931), 
	.C2(n17102), 
	.C1(n4767), 
	.B2(n16792), 
	.B1(FE_PHN1717_n5114), 
	.A2(n318), 
	.A1(n1156));
   INV_X1 U825 (.ZN(n1156), 
	.A(haddr_o[19]));
   OAI222_X1 U826 (.ZN(n4932), 
	.C2(n17102), 
	.C1(n4768), 
	.B2(n16792), 
	.B1(FE_PHN3102_n5237), 
	.A2(n318), 
	.A1(n1157));
   OAI222_X1 U827 (.ZN(n4933), 
	.C2(n17102), 
	.C1(n4769), 
	.B2(n16792), 
	.B1(FE_PHN3097_n5236), 
	.A2(n318), 
	.A1(n1158));
   OAI222_X1 U828 (.ZN(n4934), 
	.C2(n17102), 
	.C1(n4770), 
	.B2(n16792), 
	.B1(FE_PHN3101_n5235), 
	.A2(n318), 
	.A1(n1159));
   OAI222_X1 U831 (.ZN(n4937), 
	.C2(n17102), 
	.C1(n4830), 
	.B2(n16792), 
	.B1(n4812), 
	.A2(n318), 
	.A1(n952));
   INV_X1 U833 (.ZN(n963), 
	.A(haddr_o[11]));
   OAI222_X1 U834 (.ZN(n4939), 
	.C2(n17102), 
	.C1(n4771), 
	.B2(n16792), 
	.B1(n4811), 
	.A2(n17103), 
	.A1(n948));
   INV_X1 U835 (.ZN(n4940), 
	.A(n1160));
   AOI222_X1 U836 (.ZN(n1160), 
	.C2(n866), 
	.C1(n1161), 
	.B2(n16738), 
	.B1(vis_pc_o[7]), 
	.A2(n17104), 
	.A1(haddr_o[8]));
   INV_X1 U838 (.ZN(n4941), 
	.A(n1162));
   AOI222_X1 U839 (.ZN(n1162), 
	.C2(n866), 
	.C1(n1163), 
	.B2(n16738), 
	.B1(FE_PHN1341_SYNOPSYS_UNCONNECTED_531), 
	.A2(n17104), 
	.A1(haddr_o[15]));
   AOI22_X1 U844 (.ZN(n1164), 
	.B2(vis_ipsr_o[5]), 
	.B1(n322), 
	.A2(vis_pc_o[4]), 
	.A1(n16738));
   AOI22_X1 U847 (.ZN(n1165), 
	.B2(vis_ipsr_o[4]), 
	.B1(n322), 
	.A2(vis_pc_o[3]), 
	.A1(n16738));
   INV_X1 U848 (.ZN(n322), 
	.A(n324));
   NAND2_X1 U849 (.ZN(n324), 
	.A2(n17102), 
	.A1(n784));
   NAND2_X2 U853 (.ZN(n318), 
	.A2(n1166), 
	.A1(n17102));
   OAI211_X1 U854 (.ZN(n1166), 
	.C2(n692), 
	.C1(n16843), 
	.B(n762), 
	.A(n1167));
   OAI21_X1 U855 (.ZN(n1167), 
	.B2(n931), 
	.B1(n16659), 
	.A(n17097));
   AOI222_X1 U859 (.ZN(n1171), 
	.C2(n1175), 
	.C1(n16820), 
	.B2(FE_OFN631_n16851), 
	.B1(n1174), 
	.A2(n1173), 
	.A1(n1172));
   OAI221_X1 U860 (.ZN(n1175), 
	.C2(n1027), 
	.C1(n846), 
	.B2(n1176), 
	.B1(n16811), 
	.A(n1177));
   OAI211_X1 U861 (.ZN(n1168), 
	.C2(n1178), 
	.C1(FE_OFN84_n16839), 
	.B(n1180), 
	.A(n1179));
   NOR3_X1 U862 (.ZN(n1180), 
	.A3(n1183), 
	.A2(n1182), 
	.A1(n1181));
   AOI211_X1 U863 (.ZN(n1183), 
	.C2(n548), 
	.C1(n679), 
	.B(n478), 
	.A(n479));
   NOR3_X1 U864 (.ZN(n1181), 
	.A3(n1184), 
	.A2(n16795), 
	.A1(n580));
   NAND3_X1 U865 (.ZN(n1179), 
	.A3(n506), 
	.A2(FE_OFN87_n16848), 
	.A1(n16854));
   OAI22_X1 U866 (.ZN(n4945), 
	.B2(n1186), 
	.B1(hprot_o[3]), 
	.A2(n1185), 
	.A1(n4846));
   INV_X1 U867 (.ZN(n1186), 
	.A(n1185));
   NOR2_X1 U868 (.ZN(n1185), 
	.A2(FE_PHN674_n17127), 
	.A1(n999));
   OAI21_X1 U869 (.ZN(n5649), 
	.B2(n200), 
	.B1(FE_PHN674_n17127), 
	.A(n194));
   INV_X1 U870 (.ZN(n5648), 
	.A(n422));
   OAI22_X1 U871 (.ZN(n5650), 
	.B2(n1187), 
	.B1(n1078), 
	.A2(n1076), 
	.A1(n5504));
   INV_X1 U872 (.ZN(n1076), 
	.A(n1078));
   NAND3_X1 U873 (.ZN(n1078), 
	.A3(n1189), 
	.A2(n253), 
	.A1(n1188));
   OAI22_X1 U874 (.ZN(n5651), 
	.B2(n1071), 
	.B1(n5098), 
	.A2(n1187), 
	.A1(n1070));
   OAI22_X1 U875 (.ZN(n5652), 
	.B2(n1071), 
	.B1(n4961), 
	.A2(n1070), 
	.A1(n1190));
   INV_X1 U876 (.ZN(n1071), 
	.A(n1070));
   NAND2_X1 U877 (.ZN(n1070), 
	.A2(n253), 
	.A1(n1191));
   OAI22_X1 U878 (.ZN(n5653), 
	.B2(FE_PHN3496_n262), 
	.B1(n17095), 
	.A2(n17094), 
	.A1(n1190));
   AOI21_X1 U881 (.ZN(n9972), 
	.B2(FE_PHN674_n17127), 
	.B1(n16837), 
	.A(n1192));
   NOR4_X1 U882 (.ZN(n1192), 
	.A4(n1196), 
	.A3(n1195), 
	.A2(n1194), 
	.A1(n1193));
   OAI221_X1 U883 (.ZN(n1196), 
	.C2(n988), 
	.C1(FE_OFN82_n16856), 
	.B2(n1198), 
	.B1(n1197), 
	.A(n1199));
   AOI21_X1 U884 (.ZN(n1199), 
	.B2(n16820), 
	.B1(n1200), 
	.A(n1201));
   AOI22_X1 U885 (.ZN(n1197), 
	.B2(n469), 
	.B1(n630), 
	.A2(n1203), 
	.A1(n1202));
   OAI211_X1 U886 (.ZN(n1203), 
	.C2(n16674), 
	.C1(n16814), 
	.B(n17099), 
	.A(n669));
   OAI221_X1 U887 (.ZN(n1195), 
	.C2(n1087), 
	.C1(n1205), 
	.B2(n1204), 
	.B1(n16803), 
	.A(n1206));
   AOI221_X1 U888 (.ZN(n1206), 
	.C2(n1208), 
	.C1(n714), 
	.B2(n1207), 
	.B1(n844), 
	.A(n1209));
   NOR3_X1 U889 (.ZN(n1209), 
	.A3(FE_OFN95_n16864), 
	.A2(FE_OFN634_n16871), 
	.A1(n1210));
   OAI22_X1 U890 (.ZN(n1208), 
	.B2(n1212), 
	.B1(n846), 
	.A2(n1211), 
	.A1(n818));
   NAND2_X1 U891 (.ZN(n1212), 
	.A2(n16862), 
	.A1(n1213));
   INV_X1 U892 (.ZN(n844), 
	.A(n1214));
   OR2_X1 U893 (.ZN(n1087), 
	.A2(n16854), 
	.A1(n1092));
   AOI222_X1 U894 (.ZN(n1204), 
	.C2(n708), 
	.C1(n1216), 
	.B2(n630), 
	.B1(n1215), 
	.A2(n732), 
	.A1(n550));
   NOR2_X1 U895 (.ZN(n1215), 
	.A2(FE_OFN608_n16686), 
	.A1(n16868));
   OAI221_X1 U896 (.ZN(n1194), 
	.C2(n945), 
	.C1(n1218), 
	.B2(n1217), 
	.B1(n797), 
	.A(n1219));
   AOI22_X1 U897 (.ZN(n1219), 
	.B2(n482), 
	.B1(n16814), 
	.A2(n16813), 
	.A1(n1220));
   OAI221_X1 U898 (.ZN(n1193), 
	.C2(n16659), 
	.C1(n1222), 
	.B2(n713), 
	.B1(n1221), 
	.A(n1223));
   AOI222_X1 U899 (.ZN(n1223), 
	.C2(n1226), 
	.C1(n821), 
	.B2(n1225), 
	.B1(n914), 
	.A2(n1224), 
	.A1(n597));
   OAI21_X1 U900 (.ZN(n1226), 
	.B2(n1228), 
	.B1(n1227), 
	.A(n941));
   NOR3_X1 U901 (.ZN(n1227), 
	.A3(n16799), 
	.A2(n5244), 
	.A1(n1229));
   OAI21_X1 U902 (.ZN(n1229), 
	.B2(n781), 
	.B1(n16674), 
	.A(n16816));
   OAI21_X1 U903 (.ZN(n1225), 
	.B2(n1230), 
	.B1(n649), 
	.A(n1231));
   NAND4_X1 U904 (.ZN(n1231), 
	.A4(FE_OFN72_n16867), 
	.A3(FE_OFN85_n16839), 
	.A2(n610), 
	.A1(n1232));
   NAND2_X1 U905 (.ZN(n1232), 
	.A2(n1043), 
	.A1(n994));
   OAI222_X1 U906 (.ZN(n1224), 
	.C2(n617), 
	.C1(FE_OFN627_n16828), 
	.B2(n1234), 
	.B1(n16837), 
	.A2(n1233), 
	.A1(FE_OFN106_n585));
   AOI221_X1 U907 (.ZN(n1222), 
	.C2(n16817), 
	.C1(n333), 
	.B2(n16803), 
	.B1(n473), 
	.A(n1235));
   OAI221_X1 U908 (.ZN(n1235), 
	.C2(n638), 
	.C1(n16813), 
	.B2(n941), 
	.B1(n1236), 
	.A(n1237));
   NAND3_X1 U909 (.ZN(n1237), 
	.A3(n1202), 
	.A2(n16871), 
	.A1(n469));
   INV_X1 U910 (.ZN(n1202), 
	.A(n711));
   NAND2_X1 U911 (.ZN(n638), 
	.A2(n16871), 
	.A1(n16803));
   AOI221_X1 U912 (.ZN(n1236), 
	.C2(n16657), 
	.C1(n16801), 
	.B2(n1238), 
	.B1(n16796), 
	.A(n1239));
   OR2_X1 U913 (.ZN(n1239), 
	.A2(n718), 
	.A1(n833));
   AOI221_X1 U914 (.ZN(n1221), 
	.C2(n16839), 
	.C1(n16845), 
	.B2(n664), 
	.B1(n526), 
	.A(n1240));
   OAI21_X1 U915 (.ZN(n1240), 
	.B2(n16839), 
	.B1(FE_OFN98_n1104), 
	.A(n567));
   NAND2_X1 U916 (.ZN(n567), 
	.A2(n753), 
	.A1(n16845));
   AOI22_X1 U917 (.ZN(n9796), 
	.B2(FE_PHN675_n17126), 
	.B1(n16824), 
	.A2(n1242), 
	.A1(n1241));
   NOR4_X1 U918 (.ZN(n1242), 
	.A4(n1246), 
	.A3(n1245), 
	.A2(n1244), 
	.A1(n1243));
   OAI33_X1 U919 (.ZN(n1246), 
	.B3(n16821), 
	.B2(n1248), 
	.B1(n677), 
	.A3(n1247), 
	.A2(n16804), 
	.A1(n552));
   AOI21_X1 U920 (.ZN(n1248), 
	.B2(n473), 
	.B1(n1249), 
	.A(n734));
   INV_X1 U921 (.ZN(n734), 
	.A(n1176));
   NAND2_X1 U922 (.ZN(n1176), 
	.A2(n16683), 
	.A1(n934));
   NOR2_X1 U923 (.ZN(n1249), 
	.A2(FE_OFN608_n16686), 
	.A1(n931));
   NOR3_X1 U924 (.ZN(n1247), 
	.A3(n720), 
	.A2(n1251), 
	.A1(n1250));
   INV_X1 U925 (.ZN(n1251), 
	.A(n547));
   NAND3_X1 U926 (.ZN(n547), 
	.A3(n731), 
	.A2(n17098), 
	.A1(n16799));
   OAI33_X1 U927 (.ZN(n1250), 
	.B3(n718), 
	.B2(n16800), 
	.B1(n16687), 
	.A3(n16657), 
	.A2(n17098), 
	.A1(n668));
   NAND3_X1 U928 (.ZN(n552), 
	.A3(n574), 
	.A2(n16807), 
	.A1(n934));
   OAI33_X1 U929 (.ZN(n1245), 
	.B3(n723), 
	.B2(n579), 
	.B1(n569), 
	.A3(n616), 
	.A2(n1252), 
	.A1(n580));
   AOI21_X1 U930 (.ZN(n1252), 
	.B2(n16802), 
	.B1(n16725), 
	.A(n1253));
   NOR3_X1 U931 (.ZN(n1253), 
	.A3(n16796), 
	.A2(n16807), 
	.A1(n583));
   OAI33_X1 U932 (.ZN(n1244), 
	.B3(FE_OFN426_n659), 
	.B2(n576), 
	.B1(n1255), 
	.A3(n759), 
	.A2(n851), 
	.A1(n1254));
   NAND3_X1 U933 (.ZN(n576), 
	.A3(n1256), 
	.A2(n540), 
	.A1(n709));
   NOR3_X1 U934 (.ZN(n1256), 
	.A3(n444), 
	.A2(n16797), 
	.A1(n443));
   OAI21_X1 U935 (.ZN(n1255), 
	.B2(n5243), 
	.B1(n16801), 
	.A(n16799));
   OAI211_X1 U936 (.ZN(n1243), 
	.C2(n16808), 
	.C1(n1257), 
	.B(n1259), 
	.A(n1258));
   NAND4_X1 U937 (.ZN(n1259), 
	.A4(n16813), 
	.A3(n1260), 
	.A2(n16804), 
	.A1(n574));
   OAI21_X1 U938 (.ZN(n1260), 
	.B2(n843), 
	.B1(n1261), 
	.A(n478));
   INV_X1 U939 (.ZN(n574), 
	.A(n639));
   NAND2_X1 U940 (.ZN(n639), 
	.A2(n1262), 
	.A1(n475));
   INV_X1 U941 (.ZN(n1258), 
	.A(n1263));
   AOI211_X1 U942 (.ZN(n1257), 
	.C2(n1265), 
	.C1(n1264), 
	.B(n1182), 
	.A(n1266));
   NOR2_X1 U943 (.ZN(n1182), 
	.A2(n731), 
	.A1(n459));
   OAI22_X1 U944 (.ZN(n1266), 
	.B2(n640), 
	.B1(n16825), 
	.A2(n459), 
	.A1(n16797));
   NAND2_X1 U945 (.ZN(n459), 
	.A2(n482), 
	.A1(n631));
   NOR2_X1 U946 (.ZN(n1264), 
	.A2(n1267), 
	.A1(n16813));
   NOR4_X1 U947 (.ZN(n1241), 
	.A4(n1271), 
	.A3(n1270), 
	.A2(n1269), 
	.A1(n1268));
   INV_X1 U948 (.ZN(n1270), 
	.A(n1028));
   AOI221_X1 U949 (.ZN(n1028), 
	.C2(n534), 
	.C1(n528), 
	.B2(n1174), 
	.B1(n16862), 
	.A(n1272));
   INV_X1 U950 (.ZN(n1174), 
	.A(n857));
   OAI21_X1 U951 (.ZN(n1269), 
	.B2(n610), 
	.B1(n1273), 
	.A(n642));
   AOI221_X1 U952 (.ZN(n642), 
	.C2(n572), 
	.C1(n1021), 
	.B2(n612), 
	.B1(n695), 
	.A(n1274));
   NOR3_X1 U953 (.ZN(n1274), 
	.A3(n677), 
	.A2(n16725), 
	.A1(n443));
   INV_X1 U954 (.ZN(n572), 
	.A(n1019));
   NAND4_X1 U955 (.ZN(n1019), 
	.A4(n16797), 
	.A3(n505), 
	.A2(n476), 
	.A1(n540));
   AOI211_X1 U956 (.ZN(n1273), 
	.C2(n1275), 
	.C1(n660), 
	.B(n1277), 
	.A(n1276));
   NOR3_X1 U957 (.ZN(n1277), 
	.A3(n846), 
	.A2(n16821), 
	.A1(n1027));
   NOR4_X1 U958 (.ZN(n1276), 
	.A4(n664), 
	.A3(n912), 
	.A2(n650), 
	.A1(FE_OFN627_n16828));
   OAI21_X1 U959 (.ZN(n1275), 
	.B2(FE_OFN458_n860), 
	.B1(FE_OFN85_n16839), 
	.A(n607));
   OAI221_X1 U960 (.ZN(n1268), 
	.C2(n1279), 
	.C1(n605), 
	.B2(n644), 
	.B1(n1278), 
	.A(n1280));
   AOI22_X1 U961 (.ZN(n1280), 
	.B2(n1282), 
	.B1(n827), 
	.A2(n1281), 
	.A1(n751));
   OAI22_X1 U962 (.ZN(n1282), 
	.B2(n1035), 
	.B1(n16854), 
	.A2(n692), 
	.A1(n16825));
   NAND2_X1 U963 (.ZN(n1281), 
	.A2(n644), 
	.A1(n699));
   OAI22_X1 U964 (.ZN(n8706), 
	.B2(n765), 
	.B1(n1284), 
	.A2(n1283), 
	.A1(n5257));
   AOI22_X1 U965 (.ZN(n1284), 
	.B2(n659), 
	.B1(n800), 
	.A2(n16674), 
	.A1(n770));
   NAND2_X1 U966 (.ZN(n770), 
	.A2(n443), 
	.A1(n1285));
   AOI21_X1 U967 (.ZN(n1283), 
	.B2(n1286), 
	.B1(n767), 
	.A(n765));
   OAI22_X1 U968 (.ZN(n8698), 
	.B2(n765), 
	.B1(n1288), 
	.A2(n1287), 
	.A1(n5258));
   AOI22_X1 U969 (.ZN(n1288), 
	.B2(n16674), 
	.B1(n800), 
	.A2(n16798), 
	.A1(n1289));
   OAI21_X1 U970 (.ZN(n800), 
	.B2(n1184), 
	.B1(n819), 
	.A(n892));
   OAI21_X1 U971 (.ZN(n1289), 
	.B2(n443), 
	.B1(n16816), 
	.A(n1285));
   INV_X1 U972 (.ZN(n1285), 
	.A(n1290));
   OAI211_X1 U973 (.ZN(n1290), 
	.C2(n945), 
	.C1(n16821), 
	.B(n1292), 
	.A(n1291));
   AOI21_X1 U974 (.ZN(n1292), 
	.B2(n631), 
	.B1(n541), 
	.A(n1293));
   INV_X1 U975 (.ZN(n1293), 
	.A(n468));
   NAND2_X1 U976 (.ZN(n468), 
	.A2(n631), 
	.A1(n1220));
   AOI21_X1 U977 (.ZN(n1287), 
	.B2(n1294), 
	.B1(n767), 
	.A(n765));
   OAI21_X1 U978 (.ZN(n765), 
	.B2(n1296), 
	.B1(n1295), 
	.A(n17122));
   OAI211_X1 U979 (.ZN(n1296), 
	.C2(n1297), 
	.C1(n16683), 
	.B(n1298), 
	.A(n489));
   INV_X1 U980 (.ZN(n1298), 
	.A(n1299));
   AOI221_X1 U981 (.ZN(n489), 
	.C2(n1301), 
	.C1(n914), 
	.B2(n543), 
	.B1(n1300), 
	.A(n1302));
   INV_X1 U982 (.ZN(n1301), 
	.A(n1303));
   OAI221_X1 U983 (.ZN(n1295), 
	.C2(FE_OFN429_n673), 
	.C1(n498), 
	.B2(n1304), 
	.B1(n696), 
	.A(n1305));
   AOI22_X1 U984 (.ZN(n1305), 
	.B2(n990), 
	.B1(n809), 
	.A2(n195), 
	.A1(n1306));
   NAND2_X1 U985 (.ZN(n1304), 
	.A2(n808), 
	.A1(n1042));
   OAI211_X1 U986 (.ZN(n767), 
	.C2(n1307), 
	.C1(n851), 
	.B(n1309), 
	.A(n1308));
   AOI221_X1 U988 (.ZN(n1313), 
	.C2(n1316), 
	.C1(n1315), 
	.B2(n249), 
	.B1(n1314), 
	.A(n1317));
   INV_X1 U989 (.ZN(n1312), 
	.A(FE_PHN2985_IRQ_0_));
   NAND2_X1 U990 (.ZN(n1311), 
	.A2(n1318), 
	.A1(n17092));
   OAI221_X1 U991 (.ZN(n14934), 
	.C2(FE_PHN1551_n1319), 
	.C1(n379), 
	.B2(n430), 
	.B1(n373), 
	.A(n400));
   INV_X1 U992 (.ZN(n430), 
	.A(n379));
   OAI211_X1 U993 (.ZN(n14928), 
	.C2(n378), 
	.C1(FE_PHN3103_n4847), 
	.B(n1321), 
	.A(n1320));
   INV_X1 U994 (.ZN(n1321), 
	.A(n1322));
   OAI22_X1 U995 (.ZN(n1322), 
	.B2(n4974), 
	.B1(n336), 
	.A2(n334), 
	.A1(FE_PHN1551_n1319));
   NAND3_X1 U998 (.ZN(n1320), 
	.A3(n336), 
	.A2(n375), 
	.A1(n377));
   NAND3_X1 U999 (.ZN(n378), 
	.A3(n336), 
	.A2(n1323), 
	.A1(n5231));
   OAI211_X1 U1001 (.ZN(n376), 
	.C2(n1324), 
	.C1(n1054), 
	.B(n1325), 
	.A(n1107));
   INV_X1 U1002 (.ZN(n1107), 
	.A(n1326));
   NOR3_X1 U1003 (.ZN(n1324), 
	.A3(n1106), 
	.A2(n1327), 
	.A1(FE_PHN776_n1108));
   NOR2_X1 U1004 (.ZN(n1054), 
	.A2(n16868), 
	.A1(FE_PHN675_n17126));
   OAI21_X1 U1005 (.ZN(n1323), 
	.B2(n1002), 
	.B1(n4973), 
	.A(n1001));
   OAI221_X1 U1007 (.ZN(n14825), 
	.C2(n1331), 
	.C1(n1330), 
	.B2(n1329), 
	.B1(n1328), 
	.A(n1332));
   NAND3_X1 U1008 (.ZN(n1332), 
	.A3(n1329), 
	.A2(vis_tbit_o), 
	.A1(n1331));
   NAND4_X1 U1009 (.ZN(n1331), 
	.A4(n185), 
	.A3(n1010), 
	.A2(n1333), 
	.A1(n37));
   NAND2_X1 U1010 (.ZN(n1010), 
	.A2(n188), 
	.A1(n187));
   OAI211_X1 U1011 (.ZN(n1333), 
	.C2(n797), 
	.C1(n16847), 
	.B(n1335), 
	.A(n1334));
   AOI22_X1 U1012 (.ZN(n1335), 
	.B2(FE_OFN81_n16856), 
	.B1(n16836), 
	.A2(n16842), 
	.A1(n16828));
   INV_X1 U1014 (.ZN(n1330), 
	.A(n1336));
   NAND2_X1 U1015 (.ZN(n1329), 
	.A2(n17124), 
	.A1(n86));
   NOR2_X1 U1016 (.ZN(n1328), 
	.A2(FE_PHN752_n1337), 
	.A1(n1336));
   OAI22_X1 U1017 (.ZN(n1336), 
	.B2(n188), 
	.B1(n192), 
	.A2(n16785), 
	.A1(n187));
   OAI211_X1 U1018 (.ZN(n14432), 
	.C2(n379), 
	.C1(n370), 
	.B(n400), 
	.A(n1339));
   NAND3_X1 U1019 (.ZN(n1339), 
	.A3(n373), 
	.A2(n379), 
	.A1(hrdata_i[15]));
   INV_X1 U1020 (.ZN(n373), 
	.A(n377));
   NAND3_X1 U1021 (.ZN(n377), 
	.A3(n4846), 
	.A2(vis_tbit_o), 
	.A1(1'b1));
   NAND4_X1 U1025 (.ZN(n1340), 
	.A4(n16868), 
	.A3(n1001), 
	.A2(n1327), 
	.A1(n1109));
   INV_X1 U1026 (.ZN(n1327), 
	.A(n1003));
   NAND2_X1 U1028 (.ZN(n1108), 
	.A2(n375), 
	.A1(n17124));
   INV_X1 U1029 (.ZN(n400), 
	.A(n431));
   NAND2_X1 U1030 (.ZN(n431), 
	.A2(n422), 
	.A1(n5034));
   AOI21_X1 U1032 (.ZN(n1341), 
	.B2(n1342), 
	.B1(n5229), 
	.A(n1343));
   NAND3_X1 U1033 (.ZN(n1342), 
	.A3(n1345), 
	.A2(n1344), 
	.A1(n1069));
   AOI22_X1 U1034 (.ZN(n1345), 
	.B2(n1346), 
	.B1(vis_primask_o), 
	.A2(n1049), 
	.A1(n1048));
   INV_X1 U1035 (.ZN(n1346), 
	.A(n1049));
   OAI33_X1 U1036 (.ZN(n1049), 
	.B3(n1350), 
	.B2(n16824), 
	.B1(n1349), 
	.A3(n1348), 
	.A2(n16810), 
	.A1(n16656));
   NAND2_X1 U1037 (.ZN(n1349), 
	.A2(n751), 
	.A1(n897));
   OAI21_X1 U1038 (.ZN(n1048), 
	.B2(n1348), 
	.B1(n1351), 
	.A(n1352));
   NAND3_X1 U1039 (.ZN(n1352), 
	.A3(n897), 
	.A2(n1353), 
	.A1(n751));
   INV_X1 U1040 (.ZN(n1351), 
	.A(n1354));
   INV_X1 U1041 (.ZN(n1344), 
	.A(n1067));
   OAI211_X1 U1042 (.ZN(n1069), 
	.C2(n1356), 
	.C1(n1355), 
	.B(n1358), 
	.A(n1357));
   OAI21_X1 U1043 (.ZN(n1357), 
	.B2(n1360), 
	.B1(n1359), 
	.A(n1361));
   NAND4_X1 U1044 (.ZN(n1361), 
	.A4(n1365), 
	.A3(n1364), 
	.A2(n1363), 
	.A1(n1362));
   INV_X1 U1045 (.ZN(n1364), 
	.A(n1366));
   OAI21_X1 U1046 (.ZN(n1366), 
	.B2(n5503), 
	.B1(n1052), 
	.A(n1367));
   AOI211_X1 U1047 (.ZN(n1360), 
	.C2(n1368), 
	.C1(n1355), 
	.B(n1370), 
	.A(n1369));
   AOI211_X1 U1048 (.ZN(n1359), 
	.C2(n1371), 
	.C1(n1355), 
	.B(n1373), 
	.A(n1372));
   INV_X1 U1049 (.ZN(n1356), 
	.A(n1374));
   OAI22_X1 U1050 (.ZN(n1374), 
	.B2(n1370), 
	.B1(n1368), 
	.A2(n1371), 
	.A1(n1372));
   NOR3_X1 U1052 (.ZN(n14001), 
	.A3(n1377), 
	.A2(n1376), 
	.A1(n1375));
   AOI21_X1 U1053 (.ZN(n1377), 
	.B2(n1378), 
	.B1(n17092), 
	.A(n1379));
   AOI211_X1 U1055 (.ZN(n1376), 
	.C2(n247), 
	.C1(n1314), 
	.B(n1380), 
	.A(n1317));
   AOI21_X1 U1056 (.ZN(n1380), 
	.B2(n1124), 
	.B1(hwdata_o[15]), 
	.A(n1378));
   INV_X1 U1057 (.ZN(n1375), 
	.A(FE_PHN5178_IRQ_15_));
   INV_X1 U1059 (.ZN(n1383), 
	.A(FE_PHN2993_IRQ_13_));
   OAI22_X1 U1060 (.ZN(n1382), 
	.B2(n1385), 
	.B1(n242), 
	.A2(n1314), 
	.A1(n1384));
   NAND2_X1 U1061 (.ZN(n1381), 
	.A2(n1386), 
	.A1(n17092));
   AOI221_X1 U1063 (.ZN(n1389), 
	.C2(n1391), 
	.C1(n1390), 
	.B2(n218), 
	.B1(n1314), 
	.A(n1317));
   INV_X1 U1064 (.ZN(n1388), 
	.A(FE_PHN2991_IRQ_3_));
   NAND2_X1 U1065 (.ZN(n1387), 
	.A2(n1392), 
	.A1(n17092));
   AOI221_X1 U1067 (.ZN(n1395), 
	.C2(n1397), 
	.C1(n1396), 
	.B2(n215), 
	.B1(n1314), 
	.A(n1317));
   INV_X1 U1068 (.ZN(n1394), 
	.A(FE_PHN2992_IRQ_2_));
   NAND2_X1 U1069 (.ZN(n1393), 
	.A2(n1398), 
	.A1(n17092));
   AOI221_X1 U1071 (.ZN(n1401), 
	.C2(n1403), 
	.C1(n1402), 
	.B2(n229), 
	.B1(n1314), 
	.A(n1317));
   INV_X1 U1072 (.ZN(n1400), 
	.A(FE_PHN2990_IRQ_7_));
   NAND2_X1 U1073 (.ZN(n1399), 
	.A2(n1404), 
	.A1(n17092));
   AOI221_X1 U1075 (.ZN(n1407), 
	.C2(n1409), 
	.C1(n1408), 
	.B2(n226), 
	.B1(n1314), 
	.A(n1317));
   INV_X1 U1076 (.ZN(n1406), 
	.A(FE_PHN2987_IRQ_6_));
   NAND2_X1 U1077 (.ZN(n1405), 
	.A2(n1410), 
	.A1(n17092));
   AOI221_X1 U1079 (.ZN(n1414), 
	.C2(n1416), 
	.C1(n1415), 
	.B2(n224), 
	.B1(n1314), 
	.A(n1317));
   INV_X1 U1080 (.ZN(n1413), 
	.A(FE_PHN2984_IRQ_5_));
   NAND2_X1 U1081 (.ZN(n1412), 
	.A2(n1419), 
	.A1(n17092));
   AOI221_X1 U1083 (.ZN(n1422), 
	.C2(n1424), 
	.C1(n1423), 
	.B2(n1314), 
	.B1(n221), 
	.A(n1317));
   INV_X1 U1084 (.ZN(n1421), 
	.A(FE_PHN2986_IRQ_4_));
   NAND2_X1 U1085 (.ZN(n1420), 
	.A2(n1425), 
	.A1(n17092));
   OAI21_X1 U1087 (.ZN(n1427), 
	.B2(n1314), 
	.B1(n183), 
	.A(FE_PHN4631_NMI));
   INV_X1 U1088 (.ZN(n1426), 
	.A(n1429));
   AOI221_X1 U1089 (.ZN(n13846), 
	.C2(n1430), 
	.C1(n1125), 
	.B2(hwdata_o[11]), 
	.B1(n1124), 
	.A(FE_PHN1599_n1431));
   OAI21_X1 U1090 (.ZN(n1431), 
	.B2(n4755), 
	.B1(n1432), 
	.A(FE_PHN5177_IRQ_11_));
   INV_X1 U1092 (.ZN(n1435), 
	.A(FE_PHN2989_IRQ_10_));
   OAI22_X1 U1093 (.ZN(n1434), 
	.B2(n1385), 
	.B1(n236), 
	.A2(n1314), 
	.A1(n1436));
   NAND2_X1 U1094 (.ZN(n1433), 
	.A2(n1122), 
	.A1(n17092));
   INV_X1 U1096 (.ZN(n1440), 
	.A(FE_PHN2995_IRQ_8_));
   OAI22_X1 U1097 (.ZN(n1439), 
	.B2(n1385), 
	.B1(n232), 
	.A2(n1314), 
	.A1(n1441));
   NAND2_X1 U1098 (.ZN(n1438), 
	.A2(n1120), 
	.A1(n17092));
   INV_X1 U1099 (.ZN(n1120), 
	.A(n1441));
   OAI22_X1 U1101 (.ZN(n1443), 
	.B2(n1385), 
	.B1(n240), 
	.A2(n1314), 
	.A1(n1445));
   NAND2_X1 U1102 (.ZN(n1442), 
	.A2(n1446), 
	.A1(n17092));
   AOI221_X1 U1104 (.ZN(n1450), 
	.C2(n1452), 
	.C1(n1451), 
	.B2(n210), 
	.B1(n1314), 
	.A(n1317));
   INV_X1 U1105 (.ZN(n1449), 
	.A(FE_PHN4634_IRQ_1_));
   NAND2_X1 U1106 (.ZN(n1448), 
	.A2(n1453), 
	.A1(n17092));
   AND3_X1 U1107 (.ZN(n13747), 
	.A3(n1455), 
	.A2(n1454), 
	.A1(FE_PHN4641_IRQ_14_));
   OAI21_X1 U1108 (.ZN(n1455), 
	.B2(n1456), 
	.B1(n200), 
	.A(n5619));
   INV_X1 U1109 (.ZN(n1454), 
	.A(n1457));
   AOI211_X1 U1110 (.ZN(n1457), 
	.C2(n245), 
	.C1(n1314), 
	.B(n1458), 
	.A(n1317));
   AOI21_X1 U1111 (.ZN(n1458), 
	.B2(n1124), 
	.B1(hwdata_o[14]), 
	.A(n1459));
   AOI22_X1 U1113 (.ZN(n11746), 
	.B2(FE_PHN675_n17126), 
	.B1(n4950), 
	.A2(n1461), 
	.A1(n1460));
   NOR3_X1 U1114 (.ZN(n1461), 
	.A3(n1464), 
	.A2(n1463), 
	.A1(n1462));
   OAI33_X1 U1115 (.ZN(n1464), 
	.B3(n617), 
	.B2(n1218), 
	.B1(n1254), 
	.A3(n16847), 
	.A2(n5165), 
	.A1(n1465));
   OAI33_X1 U1116 (.ZN(n1463), 
	.B3(n640), 
	.B2(n1467), 
	.B1(n1466), 
	.A3(n723), 
	.A2(n16802), 
	.A1(n569));
   NAND2_X1 U1117 (.ZN(n1466), 
	.A2(FE_OFN95_n16864), 
	.A1(FE_OFN82_n16856));
   NAND3_X1 U1118 (.ZN(n569), 
	.A3(n1469), 
	.A2(n632), 
	.A1(n1468));
   OR4_X1 U1119 (.ZN(n1462), 
	.A4(n1473), 
	.A3(n1472), 
	.A2(n1471), 
	.A1(n1470));
   NOR2_X1 U1120 (.ZN(n1460), 
	.A2(n1475), 
	.A1(n1474));
   OAI211_X1 U1121 (.ZN(n1475), 
	.C2(n694), 
	.C1(n605), 
	.B(n1477), 
	.A(n1476));
   INV_X1 U1122 (.ZN(n1477), 
	.A(n1271));
   NAND3_X1 U1123 (.ZN(n1271), 
	.A3(n17122), 
	.A2(n619), 
	.A1(n988));
   NAND2_X1 U1124 (.ZN(n988), 
	.A2(n16826), 
	.A1(n1478));
   OAI221_X1 U1125 (.ZN(n1474), 
	.C2(n16808), 
	.C1(n1480), 
	.B2(n624), 
	.B1(n1479), 
	.A(n1481));
   AOI22_X1 U1126 (.ZN(n1481), 
	.B2(n1483), 
	.B1(n540), 
	.A2(n1482), 
	.A1(n526));
   OAI211_X1 U1127 (.ZN(n1483), 
	.C2(n1485), 
	.C1(n1484), 
	.B(n941), 
	.A(n1486));
   NAND3_X1 U1128 (.ZN(n1485), 
	.A3(n834), 
	.A2(n473), 
	.A1(n833));
   XOR2_X1 U1129 (.Z(n834), 
	.B(n16801), 
	.A(FE_OFN426_n659));
   NAND3_X1 U1130 (.ZN(n1484), 
	.A3(n505), 
	.A2(n16802), 
	.A1(n16814));
   INV_X1 U1131 (.ZN(n540), 
	.A(n677));
   NAND2_X1 U1132 (.ZN(n677), 
	.A2(n16659), 
	.A1(n16680));
   OAI22_X1 U1133 (.ZN(n1482), 
	.B2(n640), 
	.B1(n1205), 
	.A2(n745), 
	.A1(n16820));
   INV_X1 U1134 (.ZN(n1205), 
	.A(n1487));
   NOR4_X1 U1135 (.ZN(n1480), 
	.A4(n1491), 
	.A3(n1490), 
	.A2(n1489), 
	.A1(n1488));
   AND3_X1 U1136 (.ZN(n1489), 
	.A3(n465), 
	.A2(n4974), 
	.A1(n697));
   INV_X1 U1137 (.ZN(n465), 
	.A(n478));
   NOR2_X1 U1138 (.ZN(n697), 
	.A2(n16812), 
	.A1(n16803));
   OAI22_X1 U1139 (.ZN(n1488), 
	.B2(n499), 
	.B1(n846), 
	.A2(n818), 
	.A1(FE_OFN458_n860));
   AOI222_X1 U1140 (.ZN(n1479), 
	.C2(n16659), 
	.C1(n1495), 
	.B2(n1494), 
	.B1(n475), 
	.A2(n1493), 
	.A1(n1492));
   OAI22_X1 U1141 (.ZN(n1495), 
	.B2(n1498), 
	.B1(n1497), 
	.A2(n16802), 
	.A1(n1496));
   NAND2_X1 U1142 (.ZN(n1498), 
	.A2(n444), 
	.A1(n16807));
   NAND2_X1 U1143 (.ZN(n444), 
	.A2(n16733), 
	.A1(n731));
   INV_X1 U1144 (.ZN(n1497), 
	.A(n674));
   XOR2_X1 U1145 (.Z(n674), 
	.B(n17099), 
	.A(n1499));
   OAI211_X1 U1146 (.ZN(n1499), 
	.C2(n1501), 
	.C1(n1500), 
	.B(n1503), 
	.A(n1502));
   XOR2_X1 U1147 (.Z(n1503), 
	.B(n1505), 
	.A(n1504));
   AND3_X1 U1148 (.ZN(n1505), 
	.A3(n680), 
	.A2(n843), 
	.A1(n1506));
   AOI22_X1 U1149 (.ZN(n1506), 
	.B2(n1510), 
	.B1(n1509), 
	.A2(n1508), 
	.A1(vis_apsr_o[3]));
   OAI211_X1 U1150 (.ZN(n1504), 
	.C2(n16733), 
	.C1(n731), 
	.B(n1511), 
	.A(n843));
   OAI22_X1 U1151 (.ZN(n1511), 
	.B2(n1512), 
	.B1(n85), 
	.A2(n92), 
	.A1(vis_apsr_o[0]));
   AOI222_X1 U1152 (.ZN(n1512), 
	.C2(n27), 
	.C1(n93), 
	.B2(n94), 
	.B1(n4949), 
	.A2(U186_Z_0), 
	.A1(n16688));
   INV_X1 U1153 (.ZN(n4949), 
	.A(n93));
   NAND2_X1 U1154 (.ZN(n93), 
	.A2(n1514), 
	.A1(n1513));
   INV_X1 U1155 (.ZN(n92), 
	.A(n85));
   NOR2_X1 U1156 (.ZN(n85), 
	.A2(n1516), 
	.A1(n1515));
   OAI33_X1 U1157 (.ZN(n1516), 
	.B3(FE_OFN485_n1519), 
	.B2(n16824), 
	.B1(n1518), 
	.A3(n653), 
	.A2(FE_OFN633_n16868), 
	.A1(n1517));
   OAI211_X1 U1158 (.ZN(n1502), 
	.C2(n16814), 
	.C1(n16796), 
	.B(n1520), 
	.A(n16816));
   AOI221_X1 U1159 (.ZN(n1520), 
	.C2(n1525), 
	.C1(n1524), 
	.B2(vis_apsr_o[1]), 
	.B1(n1521), 
	.A(n736));
   AOI21_X1 U1160 (.ZN(n1501), 
	.B2(n16733), 
	.B1(n16796), 
	.A(n720));
   AOI22_X1 U1161 (.ZN(n1500), 
	.B2(n1508), 
	.B1(n1527), 
	.A2(n1509), 
	.A1(n1526));
   XOR2_X1 U1162 (.Z(n1527), 
	.B(n4954), 
	.A(n931));
   INV_X1 U1163 (.ZN(n1509), 
	.A(n1508));
   XOR2_X1 U1164 (.Z(n1526), 
	.B(n1528), 
	.A(n679));
   INV_X1 U1165 (.ZN(n679), 
	.A(n931));
   NAND2_X2 U1166 (.ZN(n931), 
	.A2(n16812), 
	.A1(n16816));
   AOI221_X1 U1167 (.ZN(n1496), 
	.C2(n17099), 
	.C1(n736), 
	.B2(n1530), 
	.B1(n1529), 
	.A(n1531));
   NAND2_X1 U1168 (.ZN(n1531), 
	.A2(n16683), 
	.A1(n582));
   NOR2_X1 U1169 (.ZN(n736), 
	.A2(n16733), 
	.A1(n16657));
   NOR3_X1 U1170 (.ZN(n1530), 
	.A3(n16814), 
	.A2(n16816), 
	.A1(n923));
   NOR3_X1 U1171 (.ZN(n1529), 
	.A3(FE_OFN426_n659), 
	.A2(n712), 
	.A1(n781));
   NAND2_X1 U1172 (.ZN(n712), 
	.A2(n16799), 
	.A1(n1532));
   OAI21_X1 U1173 (.ZN(n1494), 
	.B2(n16795), 
	.B1(n16812), 
	.A(n16807));
   NAND3_X1 U1174 (.ZN(n1493), 
	.A3(n1533), 
	.A2(n16795), 
	.A1(n720));
   AOI221_X1 U1175 (.ZN(n1533), 
	.C2(n17098), 
	.C1(n721), 
	.B2(n16800), 
	.B1(n16797), 
	.A(n1238));
   INV_X1 U1176 (.ZN(n1238), 
	.A(n669));
   AOI21_X1 U1177 (.ZN(n10553), 
	.B2(FE_PHN674_n17127), 
	.B1(FE_OFN70_n16867), 
	.A(n1534));
   NOR4_X1 U1178 (.ZN(n1534), 
	.A4(n1538), 
	.A3(n1537), 
	.A2(n1536), 
	.A1(n1535));
   OAI221_X1 U1179 (.ZN(n1538), 
	.C2(n813), 
	.C1(FE_OFN104_n715), 
	.B2(n762), 
	.B1(n16859), 
	.A(n1539));
   AOI21_X1 U1180 (.ZN(n1539), 
	.B2(FE_OFN608_n16686), 
	.B1(n1540), 
	.A(n1201));
   OAI211_X1 U1181 (.ZN(n1201), 
	.C2(n1541), 
	.C1(FE_OFN107_n585), 
	.B(n1542), 
	.A(n17122));
   NOR3_X1 U1182 (.ZN(n1542), 
	.A3(n484), 
	.A2(n1471), 
	.A1(n1543));
   INV_X1 U1183 (.ZN(n484), 
	.A(n512));
   NOR3_X1 U1184 (.ZN(n1543), 
	.A3(n16680), 
	.A2(n16824), 
	.A1(FE_OFN82_n16856));
   OAI221_X1 U1185 (.ZN(n1537), 
	.C2(n1465), 
	.C1(n606), 
	.B2(n818), 
	.B1(n649), 
	.A(n1544));
   AOI222_X1 U1186 (.ZN(n1544), 
	.C2(n1546), 
	.C1(n708), 
	.B2(n1545), 
	.B1(n822), 
	.A2(FE_OFN70_n16867), 
	.A1(n1172));
   NAND4_X1 U1187 (.ZN(n1546), 
	.A4(n1548), 
	.A3(n1547), 
	.A2(n16799), 
	.A1(n731));
   AOI211_X1 U1188 (.ZN(n1548), 
	.C2(n16733), 
	.C1(n1549), 
	.B(n718), 
	.A(n5244));
   INV_X1 U1189 (.ZN(n718), 
	.A(n1550));
   NAND3_X1 U1190 (.ZN(n1549), 
	.A3(n5243), 
	.A2(n16801), 
	.A1(n709));
   INV_X1 U1191 (.ZN(n709), 
	.A(n923));
   NAND4_X1 U1192 (.ZN(n923), 
	.A4(n16794), 
	.A3(n5241), 
	.A2(n5026), 
	.A1(n4967));
   OAI211_X1 U1193 (.ZN(n1545), 
	.C2(n1551), 
	.C1(n16804), 
	.B(n16811), 
	.A(n1552));
   NOR3_X1 U1194 (.ZN(n1551), 
	.A3(n722), 
	.A2(n16733), 
	.A1(n1553));
   OAI21_X1 U1195 (.ZN(n722), 
	.B2(n832), 
	.B1(FE_OFN608_n16686), 
	.A(n1554));
   OAI21_X1 U1196 (.ZN(n1554), 
	.B2(FE_OFN608_n16686), 
	.B1(n551), 
	.A(n16817));
   INV_X1 U1197 (.ZN(n551), 
	.A(n668));
   NAND3_X1 U1198 (.ZN(n668), 
	.A3(n1555), 
	.A2(n454), 
	.A1(n16798));
   NAND2_X1 U1199 (.ZN(n832), 
	.A2(n16798), 
	.A1(n16657));
   OAI211_X1 U1200 (.ZN(n1553), 
	.C2(n1556), 
	.C1(n1550), 
	.B(n1557), 
	.A(n548));
   NAND3_X1 U1201 (.ZN(n1557), 
	.A3(n721), 
	.A2(n16686), 
	.A1(n16796));
   NAND2_X1 U1202 (.ZN(n548), 
	.A2(n16657), 
	.A1(n939));
   NAND2_X1 U1203 (.ZN(n1556), 
	.A2(n16800), 
	.A1(n720));
   NAND2_X1 U1204 (.ZN(n1550), 
	.A2(n17099), 
	.A1(n16801));
   OAI221_X1 U1205 (.ZN(n1536), 
	.C2(n1559), 
	.C1(n16803), 
	.B2(n1558), 
	.B1(FE_OFN70_n16867), 
	.A(n1560));
   AOI22_X1 U1206 (.ZN(n1560), 
	.B2(n1094), 
	.B1(n884), 
	.A2(n1561), 
	.A1(n543));
   AOI222_X1 U1207 (.ZN(n1559), 
	.C2(n732), 
	.C1(n720), 
	.B2(n16871), 
	.B1(n1216), 
	.A2(n791), 
	.A1(n731));
   INV_X1 U1208 (.ZN(n720), 
	.A(n843));
   NAND2_X1 U1209 (.ZN(n843), 
	.A2(n16816), 
	.A1(n16796));
   INV_X1 U1210 (.ZN(n1216), 
	.A(n1562));
   AOI221_X1 U1211 (.ZN(n1558), 
	.C2(n16868), 
	.C1(n1564), 
	.B2(n563), 
	.B1(n1563), 
	.A(n1565));
   OAI22_X1 U1212 (.ZN(n1565), 
	.B2(n995), 
	.B1(n5165), 
	.A2(n859), 
	.A1(n1467));
   NAND4_X1 U1213 (.ZN(n1535), 
	.A4(n1568), 
	.A3(n1567), 
	.A2(n1308), 
	.A1(n1566));
   AOI22_X1 U1214 (.ZN(n1568), 
	.B2(n1487), 
	.B1(n746), 
	.A2(n16813), 
	.A1(n936));
   NAND2_X1 U1215 (.ZN(n1487), 
	.A2(n16820), 
	.A1(n5230));
   OAI21_X1 U1216 (.ZN(n1567), 
	.B2(n527), 
	.B1(n1172), 
	.A(n16855));
   INV_X1 U1217 (.ZN(n1172), 
	.A(n699));
   OAI21_X1 U1218 (.ZN(n1566), 
	.B2(n483), 
	.B1(n1569), 
	.A(FE_OFN78_n16834));
   OAI211_X1 U1219 (.ZN(n10055), 
	.C2(FE_PHN675_n17126), 
	.C1(n1570), 
	.B(n1572), 
	.A(n1571));
   AOI22_X1 U1220 (.ZN(n1572), 
	.B2(n16843), 
	.B1(FE_PHN675_n17126), 
	.A2(n16862), 
	.A1(n1573));
   NAND3_X1 U1221 (.ZN(n1571), 
	.A3(n687), 
	.A2(FE_OFN81_n16856), 
	.A1(n1574));
   NOR4_X1 U1222 (.ZN(n1570), 
	.A4(n1578), 
	.A3(n1577), 
	.A2(n1576), 
	.A1(n1575));
   NOR4_X1 U1223 (.ZN(n1578), 
	.A4(n1035), 
	.A3(n1580), 
	.A2(FE_OFN486_n1579), 
	.A1(n714));
   INV_X1 U1224 (.ZN(n1035), 
	.A(n660));
   INV_X1 U1225 (.ZN(n714), 
	.A(n610));
   NOR4_X1 U1226 (.ZN(n1577), 
	.A4(n995), 
	.A3(n610), 
	.A2(n994), 
	.A1(FE_OFN70_n16867));
   OAI22_X1 U1227 (.ZN(n1576), 
	.B2(n1582), 
	.B1(n1254), 
	.A2(FE_OFN100_n1086), 
	.A1(n1581));
   NAND2_X1 U1228 (.ZN(n1582), 
	.A2(n632), 
	.A1(n592));
   NAND3_X1 U1229 (.ZN(n1254), 
	.A3(n630), 
	.A2(n16802), 
	.A1(n483));
   AOI22_X1 U1230 (.ZN(n1581), 
	.B2(FE_OFN70_n16867), 
	.B1(n1583), 
	.A2(n590), 
	.A1(n1090));
   NOR2_X1 U1231 (.ZN(n1090), 
	.A2(n16828), 
	.A1(n606));
   OAI221_X1 U1232 (.ZN(n1575), 
	.C2(n616), 
	.C1(n1585), 
	.B2(n16821), 
	.B1(n1584), 
	.A(n1586));
   AOI21_X1 U1233 (.ZN(n1586), 
	.B2(n1587), 
	.B1(n16680), 
	.A(n1588));
   AOI21_X1 U1234 (.ZN(n1588), 
	.B2(n1589), 
	.B1(n618), 
	.A(n16831));
   NAND3_X1 U1235 (.ZN(n1589), 
	.A3(n612), 
	.A2(n16854), 
	.A1(n827));
   INV_X1 U1236 (.ZN(n612), 
	.A(n644));
   NAND2_X1 U1237 (.ZN(n644), 
	.A2(n597), 
	.A1(n897));
   NAND2_X1 U1238 (.ZN(n618), 
	.A2(n897), 
	.A1(n483));
   OAI221_X1 U1239 (.ZN(n1587), 
	.C2(n892), 
	.C1(n16814), 
	.B2(n1562), 
	.B1(n443), 
	.A(n1590));
   OR3_X1 U1240 (.ZN(n1590), 
	.A3(n662), 
	.A2(n650), 
	.A1(n863));
   NOR4_X1 U1241 (.ZN(n1585), 
	.A4(n1593), 
	.A3(n730), 
	.A2(n1592), 
	.A1(n1591));
   NOR3_X1 U1242 (.ZN(n1593), 
	.A3(n603), 
	.A2(n1595), 
	.A1(n1594));
   AOI211_X1 U1243 (.ZN(n1595), 
	.C2(n17098), 
	.C1(n1596), 
	.B(n1597), 
	.A(n625));
   NOR3_X1 U1244 (.ZN(n1597), 
	.A3(n1532), 
	.A2(n16799), 
	.A1(n469));
   INV_X1 U1245 (.ZN(n1532), 
	.A(n1022));
   NAND2_X1 U1246 (.ZN(n1022), 
	.A2(FE_OFN608_n16686), 
	.A1(n16801));
   NAND3_X1 U1247 (.ZN(n1596), 
	.A3(n1598), 
	.A2(n669), 
	.A1(n582));
   AOI22_X1 U1248 (.ZN(n1598), 
	.B2(n16796), 
	.B1(n16801), 
	.A2(n16817), 
	.A1(n16800));
   OAI21_X1 U1249 (.ZN(n1592), 
	.B2(n1599), 
	.B1(n16812), 
	.A(n1600));
   NAND3_X1 U1250 (.ZN(n1600), 
	.A3(n16797), 
	.A2(n16807), 
	.A1(n708));
   AOI221_X1 U1251 (.ZN(n1599), 
	.C2(n16816), 
	.C1(n708), 
	.B2(n16683), 
	.B1(n629), 
	.A(n1601));
   OAI33_X1 U1252 (.ZN(n1601), 
	.B3(n16816), 
	.B2(n16868), 
	.B1(n711), 
	.A3(n16657), 
	.A2(FE_OFN21_n503), 
	.A1(n329));
   OAI222_X1 U1253 (.ZN(n1591), 
	.C2(n580), 
	.C1(n821), 
	.B2(n512), 
	.B1(n16802), 
	.A2(n329), 
	.A1(n725));
   NAND2_X1 U1254 (.ZN(n512), 
	.A2(FE_OFN21_n503), 
	.A1(n16871));
   NOR4_X1 U1255 (.ZN(n1584), 
	.A4(n1200), 
	.A3(n848), 
	.A2(n546), 
	.A1(n1602));
   NOR3_X1 U1256 (.ZN(n848), 
	.A3(n1603), 
	.A2(n649), 
	.A1(n713));
   OAI211_X1 U1257 (.ZN(n1602), 
	.C2(n1217), 
	.C1(n556), 
	.B(n1177), 
	.A(n1604));
   OAI21_X1 U1258 (.ZN(n1604), 
	.B2(n1606), 
	.B1(n1605), 
	.A(n543));
   INV_X1 U1261 (.ZN(n1609), 
	.A(hprot_o[3]));
   OAI21_X1 U1262 (.ZN(n1608), 
	.B2(n1610), 
	.B1(haddr_o[28]), 
	.A(n999));
   OR2_X1 U1263 (.ZN(n999), 
	.A2(hprot_o[0]), 
	.A1(n1611));
   AOI21_X1 U1268 (.ZN(n1616), 
	.B2(FE_OFN115_HADDR_29_), 
	.B1(n1618), 
	.A(n1619));
   INV_X1 U1269 (.ZN(n1619), 
	.A(n1620));
   AOI22_X1 U1272 (.ZN(n1623), 
	.B2(n17090), 
	.B1(add_2072_SUM_7_), 
	.A2(n16727), 
	.A1(n17088));
   AOI22_X1 U1274 (.ZN(n1626), 
	.B2(n16722), 
	.B1(n17088), 
	.A2(n17090), 
	.A1(add_2072_SUM_6_));
   AOI221_X1 U1276 (.ZN(n1147), 
	.C2(n17088), 
	.C1(n16726), 
	.B2(n1628), 
	.B1(n1627), 
	.A(n1629));
   AND2_X1 U1277 (.ZN(n1629), 
	.A2(n17090), 
	.A1(add_2072_SUM_5_));
   NAND2_X1 U1279 (.ZN(n1633), 
	.A2(n17090), 
	.A1(add_2072_SUM_4_));
   AND2_X1 U1282 (.ZN(n1635), 
	.A2(n17090), 
	.A1(add_2072_SUM_3_));
   AND2_X1 U1285 (.ZN(n1637), 
	.A2(n17090), 
	.A1(add_2072_SUM_2_));
   AOI22_X1 U1287 (.ZN(n1639), 
	.B2(n17090), 
	.B1(add_2072_SUM_1_), 
	.A2(n16682), 
	.A1(n17088));
   AND3_X1 U1290 (.ZN(n1641), 
	.A3(n17090), 
	.A2(n1004), 
	.A1(n1642));
   OR3_X1 U1291 (.ZN(n1004), 
	.A3(n1643), 
	.A2(n4973), 
	.A1(n1106));
   OAI21_X1 U1292 (.ZN(n1642), 
	.B2(n1106), 
	.B1(n4973), 
	.A(n1643));
   XOR2_X1 U1293 (.Z(n1643), 
	.B(vis_pc_o[1]), 
	.A(n1003));
   AOI222_X1 U1295 (.ZN(n1148), 
	.C2(n16698), 
	.C1(n17088), 
	.B2(n1644), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_25_));
   AND2_X1 U1298 (.ZN(n1646), 
	.A2(n17090), 
	.A1(add_2072_SUM_24_));
   AOI222_X1 U1300 (.ZN(n1150), 
	.C2(n16655), 
	.C1(n17088), 
	.B2(n1647), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_23_));
   AOI222_X1 U1302 (.ZN(n317), 
	.C2(n16701), 
	.C1(n17088), 
	.B2(n1648), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_22_));
   AOI222_X1 U1304 (.ZN(n973), 
	.C2(n16705), 
	.C1(n17088), 
	.B2(n1649), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_21_));
   AOI222_X1 U1306 (.ZN(n1153), 
	.C2(n16702), 
	.C1(n17088), 
	.B2(n1650), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_20_));
   AND2_X1 U1309 (.ZN(n1652), 
	.A2(n17090), 
	.A1(add_2072_SUM_19_));
   AOI222_X1 U1311 (.ZN(n1155), 
	.C2(n16706), 
	.C1(n17088), 
	.B2(n1653), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_18_));
   NAND2_X1 U1314 (.ZN(n1656), 
	.A2(n17090), 
	.A1(add_2072_SUM_17_));
   AOI222_X1 U1316 (.ZN(n1157), 
	.C2(n16672), 
	.C1(n17088), 
	.B2(n1657), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_16_));
   AND2_X1 U1319 (.ZN(n1659), 
	.A2(n17090), 
	.A1(add_2072_SUM_15_));
   AOI222_X1 U1321 (.ZN(n1159), 
	.C2(n16711), 
	.C1(n17088), 
	.B2(n1660), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_14_));
   AOI22_X1 U1323 (.ZN(n1662), 
	.B2(n16715), 
	.B1(n17088), 
	.A2(n17090), 
	.A1(add_2072_SUM_13_));
   AOI222_X1 U1325 (.ZN(n956), 
	.C2(n16658), 
	.C1(n17088), 
	.B2(n1663), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_12_));
   AOI222_X1 U1327 (.ZN(n957), 
	.C2(n16679), 
	.C1(n17088), 
	.B2(n1664), 
	.B1(n1628), 
	.A2(n17090), 
	.A1(add_2072_SUM_11_));
   AND2_X1 U1330 (.ZN(n1666), 
	.A2(n17090), 
	.A1(add_2072_SUM_10_));
   AND2_X1 U1333 (.ZN(n1668), 
	.A2(n17090), 
	.A1(add_2072_SUM_8_));
   NOR2_X1 U1335 (.ZN(add_2082_A_9_), 
	.A2(n1625), 
	.A1(n17083));
   NOR2_X1 U1336 (.ZN(add_2082_A_8_), 
	.A2(n1672), 
	.A1(n17083));
   NOR2_X1 U1337 (.ZN(add_2082_A_7_), 
	.A2(n1630), 
	.A1(n17083));
   NOR2_X1 U1338 (.ZN(add_2082_A_6_), 
	.A2(n1673), 
	.A1(n17083));
   NOR2_X1 U1339 (.ZN(add_2082_A_5_), 
	.A2(n1674), 
	.A1(n17083));
   NOR2_X1 U1340 (.ZN(add_2082_A_4_), 
	.A2(n1638), 
	.A1(n17083));
   NOR3_X1 U1341 (.ZN(add_2082_A_3_), 
	.A3(n1676), 
	.A2(n17083), 
	.A1(n1675));
   NOR3_X1 U1342 (.ZN(n1675), 
	.A3(n16847), 
	.A2(n4950), 
	.A1(n890));
   NOR2_X1 U1343 (.ZN(add_2082_A_31_), 
	.A2(n1677), 
	.A1(n17083));
   NOR2_X1 U1344 (.ZN(add_2082_A_30_), 
	.A2(n1678), 
	.A1(n17083));
   NOR2_X2 U1345 (.ZN(add_2082_A_2_), 
	.A2(n1679), 
	.A1(n17083));
   NOR2_X1 U1346 (.ZN(add_2082_A_29_), 
	.A2(n1680), 
	.A1(n17083));
   NOR2_X1 U1347 (.ZN(add_2082_A_28_), 
	.A2(n1681), 
	.A1(n17083));
   NOR2_X1 U1348 (.ZN(add_2082_A_27_), 
	.A2(n1682), 
	.A1(n17083));
   NOR2_X1 U1349 (.ZN(add_2082_A_26_), 
	.A2(n17083), 
	.A1(n1683));
   NOR2_X1 U1350 (.ZN(add_2082_A_25_), 
	.A2(n1684), 
	.A1(n17083));
   NOR2_X1 U1351 (.ZN(add_2082_A_24_), 
	.A2(n1685), 
	.A1(n17083));
   NOR2_X1 U1352 (.ZN(add_2082_A_23_), 
	.A2(n1686), 
	.A1(n17083));
   NOR2_X1 U1353 (.ZN(add_2082_A_22_), 
	.A2(n1687), 
	.A1(n17083));
   NOR2_X1 U1354 (.ZN(add_2082_A_21_), 
	.A2(n1688), 
	.A1(n17083));
   NOR2_X1 U1355 (.ZN(add_2082_A_20_), 
	.A2(n1654), 
	.A1(n17083));
   NOR2_X2 U1356 (.ZN(add_2082_A_1_), 
	.A2(n1689), 
	.A1(n17083));
   NOR2_X1 U1357 (.ZN(add_2082_A_19_), 
	.A2(n1690), 
	.A1(n17083));
   NOR2_X1 U1358 (.ZN(add_2082_A_18_), 
	.A2(n1691), 
	.A1(n17083));
   NOR2_X1 U1359 (.ZN(add_2082_A_17_), 
	.A2(n1692), 
	.A1(n17083));
   NOR2_X1 U1360 (.ZN(add_2082_A_16_), 
	.A2(n1661), 
	.A1(n17083));
   NOR2_X1 U1361 (.ZN(add_2082_A_15_), 
	.A2(n17083), 
	.A1(n1693));
   AND2_X1 U1362 (.ZN(add_2082_A_14_), 
	.A2(n1514), 
	.A1(n1664));
   NOR2_X1 U1363 (.ZN(add_2082_A_13_), 
	.A2(n1694), 
	.A1(n17083));
   NOR2_X1 U1364 (.ZN(add_2082_A_12_), 
	.A2(n1695), 
	.A1(n17083));
   NOR2_X1 U1365 (.ZN(add_2082_A_11_), 
	.A2(n1696), 
	.A1(n17083));
   NOR2_X1 U1366 (.ZN(add_2082_A_10_), 
	.A2(n1621), 
	.A1(n17083));
   NAND4_X2 U1368 (.ZN(n1514), 
	.A4(n1699), 
	.A3(n1698), 
	.A2(FE_OFN10_n1697), 
	.A1(n662));
   AOI221_X1 U1369 (.ZN(n1699), 
	.C2(n16859), 
	.C1(n1095), 
	.B2(n16828), 
	.B1(n827), 
	.A(n1700));
   OAI22_X1 U1370 (.ZN(n1700), 
	.B2(FE_OFN17_n16805), 
	.B1(FE_OFN107_n585), 
	.A2(n696), 
	.A1(n16859));
   AOI22_X1 U1371 (.ZN(n1698), 
	.B2(n1574), 
	.B1(n1097), 
	.A2(n1702), 
	.A1(n1701));
   OAI211_X1 U1372 (.ZN(n1702), 
	.C2(FE_OFN17_n16805), 
	.C1(n16854), 
	.B(n998), 
	.A(n1303));
   OAI21_X1 U1373 (.ZN(n1701), 
	.B2(n617), 
	.B1(n532), 
	.A(FE_OFN610_n16690));
   NAND2_X1 U1374 (.ZN(n662), 
	.A2(FE_OFN85_n16839), 
	.A1(n526));
   NOR2_X1 U1375 (.ZN(add_2073_B_1_), 
	.A2(n1703), 
	.A1(n4950));
   AOI211_X1 U1376 (.ZN(n1703), 
	.C2(n565), 
	.C1(n589), 
	.B(n1705), 
	.A(n1704));
   OAI221_X1 U1377 (.ZN(n1704), 
	.C2(n1708), 
	.C1(FE_OFN633_n16868), 
	.B2(n1707), 
	.B1(n1706), 
	.A(n1709));
   OR4_X1 U1378 (.ZN(n1709), 
	.A4(n16865), 
	.A3(n16844), 
	.A2(n653), 
	.A1(n1278));
   INV_X1 U1379 (.ZN(n1708), 
	.A(n1710));
   OAI22_X1 U1380 (.ZN(n1710), 
	.B2(n4953), 
	.B1(n1711), 
	.A2(n16837), 
	.A1(n863));
   AOI22_X1 U1381 (.ZN(n1711), 
	.B2(n1712), 
	.B1(FE_OFN70_n16867), 
	.A2(n16851), 
	.A1(n16828));
   NAND2_X1 U1382 (.ZN(n1707), 
	.A2(n16825), 
	.A1(n1564));
   OAI22_X1 U1383 (.ZN(U98_Z_0), 
	.B2(n1715), 
	.B1(n1714), 
	.A2(n1713), 
	.A1(n5259));
   AOI211_X1 U1384 (.ZN(n1714), 
	.C2(n659), 
	.C1(n1716), 
	.B(n1718), 
	.A(n1717));
   OAI22_X1 U1385 (.ZN(n1718), 
	.B2(n1719), 
	.B1(n5241), 
	.A2(n532), 
	.A1(n5253));
   OAI221_X1 U1386 (.ZN(n1717), 
	.C2(n819), 
	.C1(n17099), 
	.B2(n1307), 
	.B1(n776), 
	.A(n1720));
   INV_X1 U1387 (.ZN(n1716), 
	.A(n1721));
   OAI22_X1 U1388 (.ZN(U97_Z_0), 
	.B2(n1715), 
	.B1(n1722), 
	.A2(n1713), 
	.A1(n5544));
   AOI211_X1 U1389 (.ZN(n1722), 
	.C2(n1723), 
	.C1(n597), 
	.B(n1725), 
	.A(n1724));
   INV_X1 U1390 (.ZN(n1725), 
	.A(n1720));
   OAI211_X1 U1391 (.ZN(n1724), 
	.C2(n1719), 
	.C1(n16794), 
	.B(n1727), 
	.A(n1726));
   NAND3_X1 U1392 (.ZN(n1727), 
	.A3(n1728), 
	.A2(n16674), 
	.A1(n16817));
   OAI21_X1 U1393 (.ZN(n1726), 
	.B2(n1730), 
	.B1(n1729), 
	.A(n614));
   INV_X1 U1394 (.ZN(n1730), 
	.A(n664));
   NOR3_X1 U1395 (.ZN(n1729), 
	.A3(FE_OFN73_n16806), 
	.A2(n16810), 
	.A1(n776));
   AOI22_X1 U1397 (.ZN(n1731), 
	.B2(n17090), 
	.B1(add_2072_SUM_9_), 
	.A2(n16719), 
	.A1(n17088));
   OAI21_X1 U1398 (.ZN(U811_Z_0), 
	.B2(n1732), 
	.B1(n5120), 
	.A(n1733));
   OAI21_X1 U1399 (.ZN(n1733), 
	.B2(n1735), 
	.B1(n1734), 
	.A(n1732));
   OAI221_X1 U1400 (.ZN(n1735), 
	.C2(n650), 
	.C1(FE_OFN81_n16856), 
	.B2(n1736), 
	.B1(n4967), 
	.A(n1737));
   AOI222_X1 U1401 (.ZN(n1737), 
	.C2(n1740), 
	.C1(n5120), 
	.B2(n16674), 
	.B1(n1739), 
	.A2(n413), 
	.A1(n1738));
   INV_X1 U1403 (.ZN(n1736), 
	.A(n1741));
   NAND4_X1 U1404 (.ZN(n1734), 
	.A4(n1743), 
	.A3(n1742), 
	.A2(n857), 
	.A1(n890));
   AOI21_X1 U1405 (.ZN(n1743), 
	.B2(n1745), 
	.B1(n1744), 
	.A(n1746));
   OAI33_X1 U1406 (.ZN(n1746), 
	.B3(n1184), 
	.B2(n16683), 
	.B1(n941), 
	.A3(FE_OFN632_n16859), 
	.A2(n16845), 
	.A1(n514));
   XOR2_X1 U1407 (.Z(n1744), 
	.B(n1748), 
	.A(n1747));
   NAND2_X1 U1408 (.ZN(n857), 
	.A2(n897), 
	.A1(n543));
   OAI22_X1 U1409 (.ZN(U810_Z_0), 
	.B2(n17082), 
	.B1(FE_OFN130_n1750), 
	.A2(n17078), 
	.A1(FE_PHN2676_n4987));
   OAI22_X1 U1410 (.ZN(U809_Z_0), 
	.B2(n1753), 
	.B1(n4953), 
	.A2(FE_PHN675_n17126), 
	.A1(n1752));
   AOI21_X1 U1411 (.ZN(n1753), 
	.B2(n84), 
	.B1(n1521), 
	.A(FE_PHN674_n17127));
   INV_X1 U1412 (.ZN(n1521), 
	.A(n1525));
   AOI221_X1 U1413 (.ZN(n1752), 
	.C2(n1755), 
	.C1(n88), 
	.B2(n1754), 
	.B1(n86), 
	.A(n1756));
   AND3_X1 U1414 (.ZN(n1756), 
	.A3(n1524), 
	.A2(n1525), 
	.A1(n84));
   INV_X1 U1415 (.ZN(n1524), 
	.A(n1757));
   AOI22_X1 U1416 (.ZN(n1757), 
	.B2(n4947), 
	.B1(U4_DATA1_0), 
	.A2(n1759), 
	.A1(n1758));
   OAI22_X1 U1417 (.ZN(n1758), 
	.B2(n1762), 
	.B1(n4953), 
	.A2(n1761), 
	.A1(n1760));
   INV_X1 U1418 (.ZN(n1761), 
	.A(n1762));
   NAND2_X1 U1419 (.ZN(n1762), 
	.A2(n1764), 
	.A1(n1763));
   AOI21_X1 U1420 (.ZN(n1760), 
	.B2(n1766), 
	.B1(n1765), 
	.A(n1767));
   AOI211_X1 U1421 (.ZN(n1767), 
	.C2(n16833), 
	.C1(n1768), 
	.B(n1769), 
	.A(n1765));
   NOR3_X1 U1422 (.ZN(n1769), 
	.A3(n1771), 
	.A2(FE_OFN628_n16833), 
	.A1(n1770));
   NOR3_X1 U1423 (.ZN(n1771), 
	.A3(n1774), 
	.A2(n1773), 
	.A1(n1772));
   INV_X1 U1424 (.ZN(n1770), 
	.A(n1775));
   AOI22_X1 U1425 (.ZN(n1775), 
	.B2(n1778), 
	.B1(n1774), 
	.A2(n1777), 
	.A1(n1776));
   OAI22_X1 U1426 (.ZN(n1778), 
	.B2(n1773), 
	.B1(n1781), 
	.A2(n1780), 
	.A1(n1779));
   INV_X1 U1427 (.ZN(n1776), 
	.A(n1782));
   OAI22_X1 U1428 (.ZN(n1766), 
	.B2(FE_OFN87_n16848), 
	.B1(n1768), 
	.A2(n1784), 
	.A1(n1783));
   AOI221_X1 U1429 (.ZN(n1768), 
	.C2(n1787), 
	.C1(n1777), 
	.B2(n1786), 
	.B1(n1785), 
	.A(n1788));
   OAI33_X1 U1430 (.ZN(n1788), 
	.B3(n1791), 
	.B2(n1790), 
	.B1(n1780), 
	.A3(n1789), 
	.A2(n1773), 
	.A1(n1774));
   NOR2_X1 U1431 (.ZN(n1785), 
	.A2(n1773), 
	.A1(n1790));
   AOI21_X1 U1432 (.ZN(n1765), 
	.B2(n1763), 
	.B1(n1792), 
	.A(n1764));
   INV_X1 U1433 (.ZN(n1764), 
	.A(n1793));
   OAI21_X1 U1434 (.ZN(n1792), 
	.B2(n1795), 
	.B1(n1794), 
	.A(n529));
   OAI221_X1 U1435 (.ZN(n1525), 
	.C2(n16824), 
	.C1(n1797), 
	.B2(FE_OFN633_n16868), 
	.B1(n1796), 
	.A(n1798));
   INV_X1 U1436 (.ZN(n1798), 
	.A(n1515));
   OAI221_X1 U1437 (.ZN(n1515), 
	.C2(n1580), 
	.C1(n1519), 
	.B2(n849), 
	.B1(n606), 
	.A(n1799));
   OAI21_X1 U1438 (.ZN(n1799), 
	.B2(n1801), 
	.B1(n1800), 
	.A(n16871));
   NOR3_X1 U1439 (.ZN(n1800), 
	.A3(FE_OFN91_n16864), 
	.A2(FE_OFN98_n1104), 
	.A1(n16826));
   AOI211_X1 U1440 (.ZN(n1797), 
	.C2(n529), 
	.C1(n1802), 
	.B(n1804), 
	.A(n1803));
   AOI21_X1 U1441 (.ZN(n1804), 
	.B2(FE_OFN87_n16848), 
	.B1(n1234), 
	.A(n849));
   INV_X1 U1442 (.ZN(n1802), 
	.A(n1210));
   AOI21_X1 U1443 (.ZN(n1796), 
	.B2(n1805), 
	.B1(FE_OFN70_n16867), 
	.A(n1806));
   OAI22_X1 U1444 (.ZN(U806_Z_0), 
	.B2(n17082), 
	.B1(n1807), 
	.A2(n17078), 
	.A1(FE_PHN2488_n4998));
   OAI22_X1 U1445 (.ZN(U805_Z_0), 
	.B2(n17082), 
	.B1(n1808), 
	.A2(n17078), 
	.A1(FE_PHN2451_n4963));
   OAI22_X1 U1446 (.ZN(U804_Z_0), 
	.B2(n17082), 
	.B1(FE_OFN128_n1809), 
	.A2(n17078), 
	.A1(FE_PHN2726_n5022));
   OAI22_X1 U1447 (.ZN(U803_Z_0), 
	.B2(n17082), 
	.B1(n1810), 
	.A2(n17078), 
	.A1(FE_PHN2741_n5040));
   OAI22_X1 U1448 (.ZN(U802_Z_0), 
	.B2(n1811), 
	.B1(n1669), 
	.A2(n980), 
	.A1(n5227));
   OAI22_X2 U1449 (.ZN(U801_Z_0), 
	.B2(n17077), 
	.B1(n1808), 
	.A2(n17074), 
	.A1(n4981));
   OAI22_X1 U1450 (.ZN(U800_Z_0), 
	.B2(n17077), 
	.B1(n1807), 
	.A2(n17074), 
	.A1(n4997));
   OAI22_X1 U1451 (.ZN(U799_Z_0), 
	.B2(n17077), 
	.B1(FE_OFN128_n1809), 
	.A2(n17074), 
	.A1(FE_PHN2735_n5021));
   OAI22_X1 U1452 (.ZN(U798_Z_0), 
	.B2(n17077), 
	.B1(FE_OFN130_n1750), 
	.A2(n17074), 
	.A1(FE_PHN2648_n4986));
   OAI22_X1 U1453 (.ZN(U797_Z_0), 
	.B2(n17077), 
	.B1(n1810), 
	.A2(n17074), 
	.A1(FE_PHN2765_n5039));
   OAI22_X1 U1454 (.ZN(U795_Z_0), 
	.B2(n1815), 
	.B1(n1814), 
	.A2(n1732), 
	.A1(n5027));
   NOR4_X1 U1455 (.ZN(n1815), 
	.A4(n1819), 
	.A3(n1818), 
	.A2(n1817), 
	.A1(n1816));
   AOI21_X1 U1456 (.ZN(n1819), 
	.B2(n1821), 
	.B1(n1820), 
	.A(n788));
   OAI21_X1 U1457 (.ZN(n1817), 
	.B2(n1822), 
	.B1(n16800), 
	.A(n1823));
   OAI211_X1 U1458 (.ZN(n1823), 
	.C2(n1825), 
	.C1(n1824), 
	.B(n1826), 
	.A(n1745));
   OAI221_X1 U1459 (.ZN(n1816), 
	.C2(n1828), 
	.C1(n5025), 
	.B2(n1827), 
	.B1(n4967), 
	.A(n1829));
   AOI22_X1 U1460 (.ZN(n1829), 
	.B2(n16674), 
	.B1(n1830), 
	.A2(n461), 
	.A1(n1741));
   OAI21_X1 U1461 (.ZN(U792_Z_0), 
	.B2(n946), 
	.B1(n1113), 
	.A(n1831));
   NAND4_X1 U1462 (.ZN(n1831), 
	.A4(n253), 
	.A3(n946), 
	.A2(FE_PHN1894_n5149), 
	.A1(n1111));
   INV_X1 U1463 (.ZN(n946), 
	.A(n256));
   NOR4_X1 U1464 (.ZN(n256), 
	.A4(haddr_o[28]), 
	.A3(n1607), 
	.A2(n1811), 
	.A1(n1610));
   AND2_X1 U1467 (.ZN(n1833), 
	.A2(n17090), 
	.A1(add_2072_SUM_26_));
   OR4_X1 U1468 (.ZN(n1607), 
	.A4(n909), 
	.A3(n17090), 
	.A2(n1834), 
	.A1(n978));
   OAI21_X1 U1469 (.ZN(n978), 
	.B2(n1614), 
	.B1(n1669), 
	.A(n1835));
   OAI22_X1 U1470 (.ZN(n1835), 
	.B2(n1836), 
	.B1(n327), 
	.A2(n1612), 
	.A1(n1613));
   INV_X1 U1471 (.ZN(n1836), 
	.A(n683));
   INV_X4 U1472 (.ZN(n1613), 
	.A(n1611));
   NAND3_X1 U1473 (.ZN(n1611), 
	.A3(n1325), 
	.A2(n1838), 
	.A1(n1837));
   NOR3_X1 U1474 (.ZN(n1325), 
	.A3(FE_OFN506_n1834), 
	.A2(lockup_o), 
	.A1(n1839));
   NAND3_X1 U1475 (.ZN(n1834), 
	.A3(n1842), 
	.A2(n1841), 
	.A1(n1840));
   AOI221_X1 U1476 (.ZN(n1842), 
	.C2(n1844), 
	.C1(n1094), 
	.B2(n746), 
	.B1(n1843), 
	.A(n1845));
   NAND3_X1 U1477 (.ZN(n1845), 
	.A3(n1092), 
	.A2(n1846), 
	.A1(n1177));
   OAI21_X1 U1478 (.ZN(n1844), 
	.B2(n1847), 
	.B1(n16680), 
	.A(n522));
   INV_X1 U1479 (.ZN(n1847), 
	.A(n1848));
   NOR2_X1 U1480 (.ZN(n1843), 
	.A2(n911), 
	.A1(FE_OFN458_n860));
   AOI222_X1 U1481 (.ZN(n1841), 
	.C2(n16821), 
	.C1(n1850), 
	.B2(n1849), 
	.B1(n799), 
	.A2(n1848), 
	.A1(n16824));
   OAI211_X1 U1482 (.ZN(n1850), 
	.C2(n1851), 
	.C1(FE_OFN458_n860), 
	.B(n1853), 
	.A(n1852));
   AOI221_X1 U1483 (.ZN(n1853), 
	.C2(n16868), 
	.C1(n1855), 
	.B2(n1854), 
	.B1(n543), 
	.A(n1200));
   NOR3_X1 U1484 (.ZN(n1200), 
	.A3(n813), 
	.A2(n16854), 
	.A1(n16824));
   NOR2_X1 U1485 (.ZN(n1855), 
	.A2(n1784), 
	.A1(n16859));
   OAI21_X1 U1486 (.ZN(n1854), 
	.B2(FE_OFN85_n16839), 
	.B1(n649), 
	.A(n1856));
   INV_X1 U1487 (.ZN(n649), 
	.A(n753));
   OAI21_X1 U1488 (.ZN(n1852), 
	.B2(n16824), 
	.B1(n1213), 
	.A(n1569));
   INV_X1 U1489 (.ZN(n1569), 
	.A(n818));
   INV_X1 U1490 (.ZN(n1213), 
	.A(n556));
   INV_X1 U1491 (.ZN(n1851), 
	.A(n746));
   NOR2_X1 U1492 (.ZN(n746), 
	.A2(n16848), 
	.A1(n859));
   NAND2_X1 U1493 (.ZN(n859), 
	.A2(n610), 
	.A1(n527));
   OAI22_X1 U1494 (.ZN(n1849), 
	.B2(n1307), 
	.B1(FE_OFN107_n585), 
	.A2(FE_OFN104_n715), 
	.A1(n16833));
   OAI211_X1 U1495 (.ZN(n1848), 
	.C2(n1857), 
	.C1(FE_OFN107_n585), 
	.B(n1859), 
	.A(n1858));
   AOI21_X1 U1496 (.ZN(n1859), 
	.B2(n527), 
	.B1(n798), 
	.A(n16826));
   NAND3_X1 U1497 (.ZN(n1858), 
	.A3(n608), 
	.A2(n808), 
	.A1(n728));
   AOI21_X1 U1498 (.ZN(n1840), 
	.B2(n608), 
	.B1(n565), 
	.A(n701));
   OAI21_X1 U1499 (.ZN(n701), 
	.B2(n522), 
	.B1(n673), 
	.A(n1860));
   OAI33_X1 U1502 (.ZN(n1862), 
	.B3(n16828), 
	.B2(n1863), 
	.B1(n532), 
	.A3(n1023), 
	.A2(n16680), 
	.A1(n524));
   AOI21_X1 U1503 (.ZN(n1863), 
	.B2(n502), 
	.B1(FE_OFN466_n998), 
	.A(n1864));
   NOR4_X1 U1504 (.ZN(n1864), 
	.A4(n918), 
	.A3(n617), 
	.A2(n579), 
	.A1(n5228));
   AOI21_X1 U1505 (.ZN(n1861), 
	.B2(n1846), 
	.B1(n1865), 
	.A(n5228));
   NAND4_X1 U1506 (.ZN(n1846), 
	.A4(n16854), 
	.A3(n1574), 
	.A2(n991), 
	.A1(n997));
   INV_X1 U1507 (.ZN(n1865), 
	.A(n1866));
   OAI22_X1 U1508 (.ZN(n1838), 
	.B2(n375), 
	.B1(n16868), 
	.A2(n1326), 
	.A1(n1867));
   NOR2_X1 U1510 (.ZN(n1867), 
	.A2(n1003), 
	.A1(n4973));
   OAI21_X1 U1511 (.ZN(n1003), 
	.B2(n187), 
	.B1(n1007), 
	.A(n1009));
   OAI21_X1 U1513 (.ZN(n1837), 
	.B2(n1001), 
	.B1(n1326), 
	.A(n4973));
   INV_X1 U1514 (.ZN(n1001), 
	.A(n1106));
   NOR2_X1 U1515 (.ZN(n1326), 
	.A2(n1007), 
	.A1(n188));
   AOI21_X1 U1516 (.ZN(n188), 
	.B2(n1868), 
	.B1(FE_OFN81_n16856), 
	.A(n727));
   INV_X1 U1517 (.ZN(n1669), 
	.A(n327));
   OAI22_X1 U1518 (.ZN(n327), 
	.B2(n1622), 
	.B1(n1689), 
	.A2(n16785), 
	.A1(n1632));
   NAND3_X1 U1520 (.ZN(n1610), 
	.A3(SPCPT1_HADDR_29_), 
	.A2(FE_OFN117_HADDR_31_), 
	.A1(haddr_o[30]));
   NAND2_X1 U1522 (.ZN(n1869), 
	.A2(n17090), 
	.A1(add_2072_SUM_27_));
   AOI22_X1 U1523 (.ZN(n1620), 
	.B2(n1628), 
	.B1(n1870), 
	.A2(n17088), 
	.A1(n16693));
   INV_X2 U1525 (.ZN(n1871), 
	.A(n1617));
   OAI22_X1 U1526 (.ZN(n1617), 
	.B2(n1622), 
	.B1(n1872), 
	.A2(n1632), 
	.A1(n27));
   INV_X4 U1527 (.ZN(n27), 
	.A(n16688));
   XOR2_X1 U1528 (.Z(n1618), 
	.B(add_2072_carry[29]), 
	.A(n5006));
   NAND2_X1 U1530 (.ZN(n1874), 
	.A2(n17090), 
	.A1(add_2072_SUM_28_));
   INV_X1 U1532 (.ZN(n1113), 
	.A(hwrite_o));
   OAI21_X1 U1534 (.ZN(n1878), 
	.B2(n1880), 
	.B1(n1879), 
	.A(n195));
   NOR3_X1 U1535 (.ZN(n1879), 
	.A3(n918), 
	.A2(n616), 
	.A1(n860));
   NOR2_X1 U1536 (.ZN(n1877), 
	.A2(n1881), 
	.A1(n742));
   NOR4_X1 U1537 (.ZN(n1881), 
	.A4(n1303), 
	.A3(n653), 
	.A2(n1882), 
	.A1(n16808));
   NOR2_X1 U1538 (.ZN(n742), 
	.A2(n1303), 
	.A1(n995));
   NAND2_X1 U1539 (.ZN(n995), 
	.A2(n16825), 
	.A1(n608));
   INV_X1 U1540 (.ZN(n1875), 
	.A(n1883));
   OAI22_X1 U1541 (.ZN(U791_Z_0), 
	.B2(n1886), 
	.B1(n226), 
	.A2(n1885), 
	.A1(n1884));
   OAI22_X1 U1542 (.ZN(U790_Z_0), 
	.B2(n1886), 
	.B1(n229), 
	.A2(n1884), 
	.A1(FE_PHN2621_n5521));
   OAI22_X1 U1543 (.ZN(U789_Z_0), 
	.B2(n1886), 
	.B1(n245), 
	.A2(n1884), 
	.A1(n5151));
   OAI22_X1 U1544 (.ZN(U788_Z_0), 
	.B2(n1886), 
	.B1(n247), 
	.A2(n1884), 
	.A1(n5150));
   OAI22_X1 U1545 (.ZN(U787_Z_0), 
	.B2(n1886), 
	.B1(n19), 
	.A2(n1884), 
	.A1(n5152));
   OAI22_X1 U1547 (.ZN(U786_Z_0), 
	.B2(n1886), 
	.B1(n1190), 
	.A2(n1884), 
	.A1(n5153));
   OAI22_X1 U1548 (.ZN(U785_Z_0), 
	.B2(n1886), 
	.B1(n1077), 
	.A2(n1884), 
	.A1(n5154));
   OAI22_X1 U1549 (.ZN(U784_Z_0), 
	.B2(n1886), 
	.B1(n1187), 
	.A2(n1884), 
	.A1(n5155));
   INV_X1 U1550 (.ZN(n1884), 
	.A(n1886));
   OAI22_X1 U1552 (.ZN(U783_Z_0), 
	.B2(n1889), 
	.B1(n226), 
	.A2(n1888), 
	.A1(n5518));
   OAI22_X1 U1553 (.ZN(U782_Z_0), 
	.B2(n1889), 
	.B1(n229), 
	.A2(n1888), 
	.A1(n5522));
   OAI22_X1 U1554 (.ZN(U781_Z_0), 
	.B2(n1889), 
	.B1(n245), 
	.A2(n1888), 
	.A1(n5157));
   OAI22_X1 U1555 (.ZN(U780_Z_0), 
	.B2(n1889), 
	.B1(n247), 
	.A2(n1888), 
	.A1(n5156));
   OAI22_X1 U1556 (.ZN(U779_Z_0), 
	.B2(n1889), 
	.B1(n19), 
	.A2(n1888), 
	.A1(n5158));
   OAI22_X1 U1557 (.ZN(U778_Z_0), 
	.B2(n1889), 
	.B1(n1190), 
	.A2(n1888), 
	.A1(FE_PHN2623_n5159));
   OAI22_X1 U1558 (.ZN(U777_Z_0), 
	.B2(n1889), 
	.B1(n1077), 
	.A2(n1888), 
	.A1(n5160));
   OAI22_X1 U1559 (.ZN(U776_Z_0), 
	.B2(n1889), 
	.B1(n1187), 
	.A2(n1888), 
	.A1(FE_PHN2739_n5161));
   INV_X1 U1560 (.ZN(n1888), 
	.A(n1889));
   OAI22_X1 U1562 (.ZN(U775_Z_0), 
	.B2(n1892), 
	.B1(n226), 
	.A2(n1891), 
	.A1(n5519));
   OAI22_X1 U1563 (.ZN(U774_Z_0), 
	.B2(n1892), 
	.B1(n229), 
	.A2(n1891), 
	.A1(n5523));
   OAI22_X1 U1564 (.ZN(U773_Z_0), 
	.B2(n1892), 
	.B1(n245), 
	.A2(n1891), 
	.A1(FE_PHN2730_n5046));
   OAI22_X1 U1565 (.ZN(U772_Z_0), 
	.B2(n1892), 
	.B1(n247), 
	.A2(n1891), 
	.A1(n5023));
   OAI22_X1 U1566 (.ZN(U771_Z_0), 
	.B2(n1892), 
	.B1(n19), 
	.A2(n1891), 
	.A1(n5053));
   OAI22_X1 U1567 (.ZN(U770_Z_0), 
	.B2(n1892), 
	.B1(n1190), 
	.A2(n1891), 
	.A1(n5008));
   OAI22_X1 U1568 (.ZN(U769_Z_0), 
	.B2(n1892), 
	.B1(n1077), 
	.A2(n1891), 
	.A1(n5009));
   OAI22_X1 U1569 (.ZN(U768_Z_0), 
	.B2(n1892), 
	.B1(n1187), 
	.A2(n1891), 
	.A1(FE_PHN2684_n5010));
   INV_X1 U1570 (.ZN(n1891), 
	.A(n1892));
   OAI22_X1 U1572 (.ZN(U767_Z_0), 
	.B2(n1895), 
	.B1(n226), 
	.A2(n1894), 
	.A1(FE_PHN2476_n5548));
   OAI22_X1 U1573 (.ZN(U766_Z_0), 
	.B2(n1895), 
	.B1(n229), 
	.A2(n1894), 
	.A1(n5549));
   OAI22_X1 U1574 (.ZN(U765_Z_0), 
	.B2(n1895), 
	.B1(n245), 
	.A2(n1894), 
	.A1(FE_PHN2691_n5550));
   OAI22_X1 U1575 (.ZN(U764_Z_0), 
	.B2(n1895), 
	.B1(n247), 
	.A2(n1894), 
	.A1(n5547));
   OAI22_X1 U1576 (.ZN(U763_Z_0), 
	.B2(n1895), 
	.B1(n19), 
	.A2(n1896), 
	.A1(n1894));
   OAI22_X1 U1577 (.ZN(U762_Z_0), 
	.B2(n1895), 
	.B1(n1190), 
	.A2(n1894), 
	.A1(n5551));
   OAI22_X1 U1578 (.ZN(U761_Z_0), 
	.B2(n1895), 
	.B1(n1077), 
	.A2(n1894), 
	.A1(n5552));
   OAI22_X1 U1579 (.ZN(U760_Z_0), 
	.B2(n1895), 
	.B1(n1187), 
	.A2(n1894), 
	.A1(FE_PHN2753_n5553));
   INV_X1 U1580 (.ZN(n1894), 
	.A(n1895));
   OAI22_X1 U1582 (.ZN(U756_Z_0), 
	.B2(n1899), 
	.B1(n16809), 
	.A2(n1898), 
	.A1(n1814));
   AOI21_X1 U1583 (.ZN(n1899), 
	.B2(n1900), 
	.B1(n1740), 
	.A(n1814));
   NOR4_X1 U1584 (.ZN(n1898), 
	.A4(n1903), 
	.A3(n1818), 
	.A2(n1902), 
	.A1(n1901));
   NOR3_X1 U1585 (.ZN(n1903), 
	.A3(n16656), 
	.A2(n788), 
	.A1(n1900));
   INV_X1 U1586 (.ZN(n788), 
	.A(n1740));
   INV_X1 U1587 (.ZN(n1818), 
	.A(n1742));
   NAND2_X1 U1588 (.ZN(n1742), 
	.A2(n1904), 
	.A1(n527));
   OAI21_X1 U1589 (.ZN(n1904), 
	.B2(FE_OFN81_n16856), 
	.B1(n5241), 
	.A(n605));
   OAI22_X1 U1590 (.ZN(n1902), 
	.B2(n1906), 
	.B1(n1905), 
	.A2(n1822), 
	.A1(n17099));
   XNOR2_X1 U1591 (.ZN(n1906), 
	.B(n1907), 
	.A(n1826));
   INV_X1 U1592 (.ZN(n1905), 
	.A(n1745));
   INV_X1 U1593 (.ZN(n1822), 
	.A(n1739));
   NAND2_X1 U1594 (.ZN(n1739), 
	.A2(n1909), 
	.A1(n1908));
   OAI221_X1 U1595 (.ZN(n1901), 
	.C2(n1828), 
	.C1(n175), 
	.B2(n1827), 
	.B1(n5026), 
	.A(n1910));
   AOI22_X1 U1596 (.ZN(n1910), 
	.B2(n16798), 
	.B1(n1830), 
	.A2(n454), 
	.A1(n1741));
   INV_X1 U1597 (.ZN(n1830), 
	.A(n772));
   INV_X1 U1599 (.ZN(n1814), 
	.A(n1732));
   OAI21_X1 U1600 (.ZN(U755_Z_0), 
	.B2(n1732), 
	.B1(n5100), 
	.A(n1911));
   OAI21_X1 U1601 (.ZN(n1911), 
	.B2(n1913), 
	.B1(n1912), 
	.A(n1732));
   OAI221_X1 U1602 (.ZN(n1913), 
	.C2(n524), 
	.C1(FE_OFN632_n16859), 
	.B2(n772), 
	.B1(n17099), 
	.A(n1914));
   AOI222_X1 U1603 (.ZN(n1914), 
	.C2(n415), 
	.C1(n1738), 
	.B2(n16657), 
	.B1(n1915), 
	.A2(n16734), 
	.A1(n1741));
   INV_X1 U1605 (.ZN(n1738), 
	.A(n1828));
   OAI21_X1 U1606 (.ZN(n1828), 
	.B2(n1916), 
	.B1(n807), 
	.A(n194));
   NOR2_X1 U1608 (.ZN(n1916), 
	.A2(n745), 
	.A1(n998));
   INV_X1 U1609 (.ZN(n1915), 
	.A(n1909));
   OAI21_X1 U1610 (.ZN(n1909), 
	.B2(n792), 
	.B1(n1917), 
	.A(n16811));
   AND2_X1 U1611 (.ZN(n792), 
	.A2(n16820), 
	.A1(n936));
   NOR2_X1 U1612 (.ZN(n936), 
	.A2(n16868), 
	.A1(n1552));
   NOR2_X1 U1613 (.ZN(n1917), 
	.A2(n478), 
	.A1(n579));
   OAI211_X1 U1614 (.ZN(n1741), 
	.C2(n945), 
	.C1(n851), 
	.B(n1918), 
	.A(n1291));
   AOI21_X1 U1615 (.ZN(n1918), 
	.B2(n16816), 
	.B1(n476), 
	.A(n1919));
   NOR4_X1 U1616 (.ZN(n1919), 
	.A4(n1184), 
	.A3(n1261), 
	.A2(n16659), 
	.A1(n16814));
   AOI22_X1 U1617 (.ZN(n1291), 
	.B2(n482), 
	.B1(n466), 
	.A2(n476), 
	.A1(n1920));
   NOR2_X1 U1618 (.ZN(n482), 
	.A2(n16811), 
	.A1(n819));
   NAND2_X1 U1619 (.ZN(n772), 
	.A2(n466), 
	.A1(n1220));
   OAI221_X1 U1620 (.ZN(n1912), 
	.C2(n1827), 
	.C1(n5241), 
	.B2(n1908), 
	.B1(n680), 
	.A(n1921));
   AOI221_X1 U1621 (.ZN(n1921), 
	.C2(n1745), 
	.C1(n1923), 
	.B2(n1740), 
	.B1(n1922), 
	.A(n799));
   OAI33_X1 U1622 (.ZN(n1745), 
	.B3(n1184), 
	.B2(n16811), 
	.B1(n940), 
	.A3(n443), 
	.A2(n16816), 
	.A1(n1920));
   NAND2_X1 U1623 (.ZN(n940), 
	.A2(n16733), 
	.A1(n822));
   OAI22_X1 U1624 (.ZN(n1923), 
	.B2(n1826), 
	.B1(n1907), 
	.A2(n1925), 
	.A1(n1924));
   NAND2_X1 U1625 (.ZN(n1826), 
	.A2(n1825), 
	.A1(n1824));
   XOR2_X1 U1626 (.Z(n1825), 
	.B(n1927), 
	.A(n1926));
   AND2_X1 U1627 (.ZN(n1824), 
	.A2(n1747), 
	.A1(n1748));
   INV_X1 U1628 (.ZN(n1747), 
	.A(n1928));
   AOI21_X1 U1629 (.ZN(n1748), 
	.B2(n16800), 
	.B1(n1929), 
	.A(n1927));
   XNOR2_X1 U1630 (.ZN(n1907), 
	.B(n1924), 
	.A(n1925));
   NAND2_X1 U1631 (.ZN(n1925), 
	.A2(n1926), 
	.A1(n1927));
   XOR2_X1 U1632 (.Z(n1926), 
	.B(n1931), 
	.A(n1930));
   NOR2_X1 U1633 (.ZN(n1927), 
	.A2(n16799), 
	.A1(n1929));
   OAI21_X1 U1634 (.ZN(n1929), 
	.B2(n16674), 
	.B1(n1932), 
	.A(n1933));
   XOR2_X1 U1635 (.Z(n1924), 
	.B(n1935), 
	.A(n1934));
   AOI22_X1 U1636 (.ZN(n1935), 
	.B2(n1937), 
	.B1(n1936), 
	.A2(n1931), 
	.A1(n1930));
   XOR2_X1 U1637 (.Z(n1931), 
	.B(n1936), 
	.A(n1937));
   XOR2_X1 U1638 (.Z(n1937), 
	.B(n1939), 
	.A(n1938));
   INV_X1 U1639 (.ZN(n1930), 
	.A(n1933));
   NAND2_X1 U1640 (.ZN(n1933), 
	.A2(n16674), 
	.A1(n1932));
   AOI21_X1 U1641 (.ZN(n1932), 
	.B2(n5244), 
	.B1(n1940), 
	.A(n1936));
   NOR2_X1 U1642 (.ZN(n1936), 
	.A2(n5244), 
	.A1(n1940));
   OAI21_X1 U1643 (.ZN(n1940), 
	.B2(n1941), 
	.B1(n781), 
	.A(n1938));
   OAI22_X1 U1644 (.ZN(n1934), 
	.B2(n1943), 
	.B1(n1942), 
	.A2(n1938), 
	.A1(n1939));
   NAND2_X1 U1645 (.ZN(n1938), 
	.A2(n781), 
	.A1(n1941));
   XOR2_X1 U1646 (.Z(n1941), 
	.B(n1944), 
	.A(n16794));
   XNOR2_X1 U1647 (.ZN(n1939), 
	.B(n1942), 
	.A(n1943));
   AOI21_X1 U1648 (.ZN(n1942), 
	.B2(n1945), 
	.B1(n454), 
	.A(n1555));
   NOR2_X1 U1649 (.ZN(n1555), 
	.A2(n5026), 
	.A1(n4967));
   OR2_X1 U1650 (.ZN(n1943), 
	.A2(n16794), 
	.A1(n1944));
   XOR2_X1 U1651 (.Z(n1944), 
	.B(n1945), 
	.A(n5241));
   XNOR2_X1 U1652 (.ZN(n1945), 
	.B(n4967), 
	.A(n461));
   OAI221_X1 U1653 (.ZN(n1740), 
	.C2(n1093), 
	.C1(n16854), 
	.B2(n514), 
	.B1(n860), 
	.A(n1309));
   AOI22_X1 U1654 (.ZN(n1309), 
	.B2(n1946), 
	.B1(n589), 
	.A2(n1573), 
	.A1(n16862));
   INV_X1 U1655 (.ZN(n1093), 
	.A(n1583));
   XOR2_X1 U1656 (.Z(n1922), 
	.B(n795), 
	.A(n794));
   NOR2_X1 U1657 (.ZN(n794), 
	.A2(n16809), 
	.A1(n1900));
   OAI21_X1 U1658 (.ZN(n1827), 
	.B2(n732), 
	.B1(n1540), 
	.A(n631));
   INV_X1 U1659 (.ZN(n631), 
	.A(n1184));
   NAND2_X1 U1660 (.ZN(n1184), 
	.A2(n16802), 
	.A1(n16820));
   NAND2_X1 U1661 (.ZN(n680), 
	.A2(n16657), 
	.A1(n16812));
   OAI21_X1 U1662 (.ZN(n1732), 
	.B2(FE_PHN675_n17126), 
	.B1(n1947), 
	.A(n1948));
   NAND3_X1 U1663 (.ZN(n1948), 
	.A3(n687), 
	.A2(n911), 
	.A1(n827));
   INV_X1 U1664 (.ZN(n687), 
	.A(n1059));
   NAND2_X1 U1665 (.ZN(n1059), 
	.A2(FE_OFN17_n16805), 
	.A1(n17124));
   NOR4_X1 U1666 (.ZN(n1947), 
	.A4(n1299), 
	.A3(n1951), 
	.A2(n1950), 
	.A1(n1949));
   NAND4_X1 U1667 (.ZN(n1299), 
	.A4(n1955), 
	.A3(n1954), 
	.A2(n1953), 
	.A1(n1952));
   NOR4_X1 U1668 (.ZN(n1955), 
	.A4(n1490), 
	.A3(n1573), 
	.A2(n1470), 
	.A1(n1956));
   NOR4_X1 U1669 (.ZN(n1490), 
	.A4(n16854), 
	.A3(FE_OFN107_n585), 
	.A2(n16689), 
	.A1(FE_OFN486_n1579));
   INV_X1 U1670 (.ZN(n1573), 
	.A(n1957));
   NOR2_X1 U1671 (.ZN(n1470), 
	.A2(n16859), 
	.A1(n1465));
   OAI22_X1 U1672 (.ZN(n1956), 
	.B2(n16657), 
	.B1(n497), 
	.A2(FE_OFN21_n503), 
	.A1(n1958));
   AOI221_X1 U1673 (.ZN(n1958), 
	.C2(n1959), 
	.C1(n934), 
	.B2(n16804), 
	.B1(n333), 
	.A(n541));
   NOR2_X1 U1674 (.ZN(n541), 
	.A2(n16812), 
	.A1(n478));
   INV_X1 U1675 (.ZN(n1959), 
	.A(n1960));
   AOI22_X1 U1676 (.ZN(n1960), 
	.B2(n833), 
	.B1(n731), 
	.A2(n505), 
	.A1(n939));
   NOR2_X1 U1677 (.ZN(n833), 
	.A2(n16797), 
	.A1(n16799));
   NOR2_X1 U1678 (.ZN(n939), 
	.A2(n17099), 
	.A1(n669));
   INV_X1 U1679 (.ZN(n934), 
	.A(n941));
   AOI222_X1 U1680 (.ZN(n1954), 
	.C2(n475), 
	.C1(n473), 
	.B2(n1472), 
	.B1(n16794), 
	.A2(n16802), 
	.A1(n1540));
   INV_X1 U1681 (.ZN(n1952), 
	.A(n510));
   OAI211_X1 U1682 (.ZN(n510), 
	.C2(n1214), 
	.C1(n1580), 
	.B(n1962), 
	.A(n1961));
   AOI22_X1 U1683 (.ZN(n1962), 
	.B2(n16659), 
	.B1(n629), 
	.A2(n16837), 
	.A1(n1472));
   NAND3_X1 U1684 (.ZN(n1961), 
	.A3(n708), 
	.A2(n1963), 
	.A1(n16807));
   NAND2_X1 U1685 (.ZN(n1214), 
	.A2(n16870), 
	.A1(n565));
   NOR2_X1 U1686 (.ZN(n1951), 
	.A2(n696), 
	.A1(n1519));
   OAI22_X1 U1687 (.ZN(n1950), 
	.B2(n692), 
	.B1(n1964), 
	.A2(FE_OFN429_n673), 
	.A1(n16820));
   OAI221_X1 U1688 (.ZN(n1949), 
	.C2(n699), 
	.C1(n610), 
	.B2(n607), 
	.B1(n762), 
	.A(n1965));
   NOR3_X1 U1689 (.ZN(n1965), 
	.A3(n1967), 
	.A2(n1491), 
	.A1(n1966));
   NOR3_X1 U1690 (.ZN(n1967), 
	.A3(n1261), 
	.A2(n16816), 
	.A1(n1267));
   NOR4_X1 U1691 (.ZN(n1491), 
	.A4(FE_OFN70_n16867), 
	.A3(n16862), 
	.A2(n797), 
	.A1(n1307));
   AND3_X1 U1692 (.ZN(n1966), 
	.A3(n16837), 
	.A2(FE_OFN450_n808), 
	.A1(n807));
   NOR2_X1 U1693 (.ZN(n807), 
	.A2(n17097), 
	.A1(n641));
   NAND2_X1 U1694 (.ZN(n607), 
	.A2(n16694), 
	.A1(n195));
   OAI22_X1 U1695 (.ZN(U754_Z_0), 
	.B2(n1715), 
	.B1(n1968), 
	.A2(n1713), 
	.A1(n5545));
   NOR2_X1 U1696 (.ZN(n1968), 
	.A2(n1970), 
	.A1(n1969));
   OAI221_X1 U1697 (.ZN(n1970), 
	.C2(n819), 
	.C1(n16800), 
	.B2(n1721), 
	.B1(n5243), 
	.A(n1170));
   OAI221_X1 U1698 (.ZN(n1969), 
	.C2(n532), 
	.C1(n5003), 
	.B2(n1307), 
	.B1(n1971), 
	.A(n1972));
   INV_X1 U1699 (.ZN(n1972), 
	.A(n1973));
   OAI21_X1 U1700 (.ZN(n1973), 
	.B2(n5026), 
	.B1(n1719), 
	.A(n694));
   AOI221_X1 U1701 (.ZN(n1971), 
	.C2(n437), 
	.C1(n1975), 
	.B2(n776), 
	.B1(n1974), 
	.A(n1976));
   OAI22_X1 U1702 (.ZN(U752_Z_0), 
	.B2(n17071), 
	.B1(n1808), 
	.A2(n17068), 
	.A1(FE_PHN2767_n5450));
   OAI22_X1 U1703 (.ZN(U751_Z_0), 
	.B2(n17071), 
	.B1(n1807), 
	.A2(n17068), 
	.A1(FE_PHN2653_n5451));
   OAI22_X1 U1704 (.ZN(U750_Z_0), 
	.B2(n17071), 
	.B1(FE_OFN128_n1809), 
	.A2(n17068), 
	.A1(FE_PHN2708_n5452));
   OAI22_X1 U1705 (.ZN(U749_Z_0), 
	.B2(n17071), 
	.B1(FE_OFN130_n1750), 
	.A2(n17068), 
	.A1(FE_PHN2711_n5453));
   OAI22_X1 U1706 (.ZN(U748_Z_0), 
	.B2(n17071), 
	.B1(n1810), 
	.A2(n17068), 
	.A1(n5454));
   OAI22_X1 U1707 (.ZN(U747_Z_0), 
	.B2(n17067), 
	.B1(n1808), 
	.A2(n17063), 
	.A1(FE_PHN2688_n5421));
   OAI22_X1 U1708 (.ZN(U746_Z_0), 
	.B2(n17067), 
	.B1(n1807), 
	.A2(n17063), 
	.A1(FE_PHN2597_n5422));
   OAI22_X1 U1709 (.ZN(U745_Z_0), 
	.B2(n17067), 
	.B1(FE_OFN128_n1809), 
	.A2(n17063), 
	.A1(n5423));
   OAI22_X1 U1710 (.ZN(U744_Z_0), 
	.B2(n17067), 
	.B1(FE_OFN130_n1750), 
	.A2(n17063), 
	.A1(FE_PHN2696_n5424));
   OAI22_X1 U1711 (.ZN(U743_Z_0), 
	.B2(n17067), 
	.B1(n1810), 
	.A2(n17063), 
	.A1(n5425));
   OAI22_X1 U1712 (.ZN(U742_Z_0), 
	.B2(n17062), 
	.B1(n1808), 
	.A2(n17058), 
	.A1(FE_PHN2725_n5392));
   OAI22_X1 U1713 (.ZN(U741_Z_0), 
	.B2(n17062), 
	.B1(n1807), 
	.A2(n17058), 
	.A1(FE_PHN2655_n5393));
   OAI22_X1 U1714 (.ZN(U740_Z_0), 
	.B2(n17062), 
	.B1(FE_OFN128_n1809), 
	.A2(n17058), 
	.A1(FE_PHN2591_n5394));
   OAI22_X1 U1715 (.ZN(U739_Z_0), 
	.B2(n17062), 
	.B1(FE_OFN130_n1750), 
	.A2(n17058), 
	.A1(FE_PHN2637_n5395));
   OAI22_X1 U1716 (.ZN(U738_Z_0), 
	.B2(n17062), 
	.B1(n1810), 
	.A2(n17058), 
	.A1(FE_PHN2759_n5396));
   OAI22_X1 U1717 (.ZN(U737_Z_0), 
	.B2(n17057), 
	.B1(n1808), 
	.A2(n17053), 
	.A1(FE_PHN2636_n5363));
   OAI22_X1 U1718 (.ZN(U736_Z_0), 
	.B2(n17057), 
	.B1(n1807), 
	.A2(n17053), 
	.A1(FE_PHN2606_n5364));
   OAI22_X1 U1719 (.ZN(U735_Z_0), 
	.B2(n17057), 
	.B1(FE_OFN128_n1809), 
	.A2(n17053), 
	.A1(FE_PHN2572_n5365));
   OAI22_X1 U1720 (.ZN(U734_Z_0), 
	.B2(n17057), 
	.B1(FE_OFN130_n1750), 
	.A2(n17053), 
	.A1(FE_PHN2716_n5366));
   OAI22_X1 U1721 (.ZN(U733_Z_0), 
	.B2(n17057), 
	.B1(n1810), 
	.A2(n17053), 
	.A1(FE_PHN2620_n5367));
   OAI22_X1 U1722 (.ZN(U732_Z_0), 
	.B2(n17052), 
	.B1(n1808), 
	.A2(n17048), 
	.A1(FE_PHN2549_n5334));
   OAI22_X1 U1723 (.ZN(U731_Z_0), 
	.B2(n17052), 
	.B1(n1807), 
	.A2(n17048), 
	.A1(FE_PHN2555_n5335));
   OAI22_X1 U1724 (.ZN(U730_Z_0), 
	.B2(n17052), 
	.B1(FE_OFN128_n1809), 
	.A2(n17048), 
	.A1(FE_PHN2566_n5336));
   OAI22_X1 U1725 (.ZN(U729_Z_0), 
	.B2(n17052), 
	.B1(FE_OFN130_n1750), 
	.A2(n17048), 
	.A1(FE_PHN2504_n5337));
   OAI22_X1 U1726 (.ZN(U728_Z_0), 
	.B2(n17052), 
	.B1(n1810), 
	.A2(n17048), 
	.A1(n5338));
   OAI22_X2 U1727 (.ZN(U727_Z_0), 
	.B2(n17046), 
	.B1(n1808), 
	.A2(n17043), 
	.A1(n5305));
   OAI22_X1 U1728 (.ZN(U726_Z_0), 
	.B2(n17046), 
	.B1(n1807), 
	.A2(n17043), 
	.A1(n5306));
   OAI22_X1 U1729 (.ZN(U725_Z_0), 
	.B2(n17046), 
	.B1(FE_OFN128_n1809), 
	.A2(n17043), 
	.A1(FE_PHN2440_n5307));
   OAI22_X1 U1730 (.ZN(U724_Z_0), 
	.B2(n17046), 
	.B1(FE_OFN130_n1750), 
	.A2(n17043), 
	.A1(FE_PHN2610_n5308));
   OAI22_X1 U1731 (.ZN(U723_Z_0), 
	.B2(n17046), 
	.B1(n1810), 
	.A2(n17043), 
	.A1(FE_PHN2604_n5309));
   OAI22_X1 U1732 (.ZN(U722_Z_0), 
	.B2(n17042), 
	.B1(n1808), 
	.A2(n17038), 
	.A1(FE_PHN2790_n5284));
   OAI22_X1 U1733 (.ZN(U721_Z_0), 
	.B2(n17042), 
	.B1(n1807), 
	.A2(n17038), 
	.A1(n5285));
   OAI22_X1 U1734 (.ZN(U720_Z_0), 
	.B2(n17042), 
	.B1(FE_OFN128_n1809), 
	.A2(n17038), 
	.A1(FE_PHN2460_n5286));
   OAI22_X1 U1735 (.ZN(U719_Z_0), 
	.B2(n17042), 
	.B1(FE_OFN130_n1750), 
	.A2(n17038), 
	.A1(FE_PHN2712_n5287));
   OAI22_X1 U1736 (.ZN(U718_Z_0), 
	.B2(n17042), 
	.B1(n1810), 
	.A2(n17038), 
	.A1(FE_PHN2785_n5288));
   OAI22_X1 U1737 (.ZN(U717_Z_0), 
	.B2(n17037), 
	.B1(n1808), 
	.A2(n17033), 
	.A1(FE_PHN2521_n5263));
   OAI22_X1 U1738 (.ZN(U716_Z_0), 
	.B2(n17037), 
	.B1(n1807), 
	.A2(n17033), 
	.A1(FE_PHN2508_n5264));
   OAI22_X1 U1739 (.ZN(U715_Z_0), 
	.B2(n17037), 
	.B1(FE_OFN128_n1809), 
	.A2(n17033), 
	.A1(FE_PHN2435_n5265));
   OAI22_X1 U1740 (.ZN(U714_Z_0), 
	.B2(n17037), 
	.B1(FE_OFN130_n1750), 
	.A2(n17033), 
	.A1(FE_PHN2625_n5266));
   OAI22_X1 U1741 (.ZN(U713_Z_0), 
	.B2(n17037), 
	.B1(n1810), 
	.A2(n17033), 
	.A1(FE_PHN2796_n5267));
   OAI22_X2 U1742 (.ZN(U712_Z_0), 
	.B2(n17031), 
	.B1(n1808), 
	.A2(n17028), 
	.A1(n4962));
   OAI22_X1 U1743 (.ZN(U711_Z_0), 
	.B2(n17031), 
	.B1(n1807), 
	.A2(n17028), 
	.A1(n4996));
   OAI22_X1 U1744 (.ZN(U710_Z_0), 
	.B2(n17031), 
	.B1(FE_OFN128_n1809), 
	.A2(n17028), 
	.A1(FE_PHN2720_n5020));
   OAI22_X1 U1745 (.ZN(U709_Z_0), 
	.B2(n17031), 
	.B1(FE_OFN130_n1750), 
	.A2(n17028), 
	.A1(FE_PHN2756_n4985));
   OAI22_X1 U1746 (.ZN(U708_Z_0), 
	.B2(n17031), 
	.B1(n1810), 
	.A2(n17028), 
	.A1(n5038));
   OAI22_X1 U1747 (.ZN(U707_Z_0), 
	.B2(n17027), 
	.B1(n1808), 
	.A2(n17023), 
	.A1(FE_PHN2781_n5169));
   OAI22_X1 U1748 (.ZN(U706_Z_0), 
	.B2(n17027), 
	.B1(n1807), 
	.A2(n17023), 
	.A1(FE_PHN2773_n5170));
   OAI22_X1 U1749 (.ZN(U705_Z_0), 
	.B2(n17027), 
	.B1(FE_OFN128_n1809), 
	.A2(n17023), 
	.A1(FE_PHN2713_n5171));
   OAI22_X1 U1750 (.ZN(U704_Z_0), 
	.B2(n17027), 
	.B1(FE_OFN130_n1750), 
	.A2(n17023), 
	.A1(FE_PHN2772_n5172));
   OAI22_X1 U1751 (.ZN(U703_Z_0), 
	.B2(n17027), 
	.B1(n1810), 
	.A2(n17023), 
	.A1(FE_PHN2764_n5173));
   OAI22_X1 U1752 (.ZN(U702_Z_0), 
	.B2(n17022), 
	.B1(n1808), 
	.A2(n17018), 
	.A1(FE_PHN2614_n4979));
   OAI22_X1 U1753 (.ZN(U701_Z_0), 
	.B2(n17022), 
	.B1(n1807), 
	.A2(n17018), 
	.A1(FE_PHN2585_n4995));
   OAI22_X1 U1754 (.ZN(U700_Z_0), 
	.B2(n17022), 
	.B1(FE_OFN128_n1809), 
	.A2(n17018), 
	.A1(FE_PHN2574_n5019));
   OAI22_X1 U1755 (.ZN(U699_Z_0), 
	.B2(n17022), 
	.B1(FE_OFN130_n1750), 
	.A2(n17018), 
	.A1(FE_PHN2501_n4984));
   OAI22_X1 U1756 (.ZN(U698_Z_0), 
	.B2(n17022), 
	.B1(n1810), 
	.A2(n17018), 
	.A1(FE_PHN2502_n5037));
   OAI22_X1 U1757 (.ZN(U697_Z_0), 
	.B2(n17017), 
	.B1(n1808), 
	.A2(n17013), 
	.A1(FE_PHN2493_n5198));
   OAI22_X1 U1758 (.ZN(U696_Z_0), 
	.B2(n17017), 
	.B1(n1807), 
	.A2(n17013), 
	.A1(FE_PHN2612_n5199));
   OAI22_X1 U1759 (.ZN(U695_Z_0), 
	.B2(n17017), 
	.B1(FE_OFN128_n1809), 
	.A2(n17013), 
	.A1(FE_PHN2568_n5200));
   OAI22_X1 U1760 (.ZN(U694_Z_0), 
	.B2(n17017), 
	.B1(FE_OFN130_n1750), 
	.A2(n17013), 
	.A1(FE_PHN2576_n5201));
   INV_X1 U1762 (.ZN(n179), 
	.A(FE_PHN719_n190));
   AOI221_X1 U1763 (.ZN(n190), 
	.C2(n2005), 
	.C1(n2004), 
	.B2(n2003), 
	.B1(n2002), 
	.A(n2006));
   INV_X1 U1764 (.ZN(n2006), 
	.A(n2007));
   AOI221_X1 U1765 (.ZN(n2007), 
	.C2(n2011), 
	.C1(n2010), 
	.B2(n2009), 
	.B1(n2008), 
	.A(FE_OFN509_n2012));
   OAI22_X1 U1766 (.ZN(U693_Z_0), 
	.B2(n17017), 
	.B1(n1810), 
	.A2(n17013), 
	.A1(FE_PHN2584_n5202));
   AOI22_X1 U1768 (.ZN(n2014), 
	.B2(n1354), 
	.B1(n17008), 
	.A2(FE_OFN2_n2015), 
	.A1(add_2073_SUM_1_));
   INV_X1 U1769 (.ZN(n2013), 
	.A(n2017));
   AOI221_X1 U1770 (.ZN(n192), 
	.C2(n2019), 
	.C1(n2002), 
	.B2(n2018), 
	.B1(n2004), 
	.A(n2020));
   INV_X2 U1771 (.ZN(n2020), 
	.A(n2021));
   AOI221_X1 U1772 (.ZN(n2021), 
	.C2(n2011), 
	.C1(n2023), 
	.B2(n2022), 
	.B1(n2008), 
	.A(n2012));
   OAI22_X1 U1773 (.ZN(U692_Z_0), 
	.B2(n2026), 
	.B1(n2025), 
	.A2(n2024), 
	.A1(n5055));
   AOI22_X1 U1774 (.ZN(n2025), 
	.B2(n2029), 
	.B1(vis_pc_o[1]), 
	.A2(n2028), 
	.A1(n2027));
   INV_X1 U1777 (.ZN(n2024), 
	.A(n2026));
   NAND2_X1 U1778 (.ZN(n2026), 
	.A2(n2030), 
	.A1(n17124));
   NAND3_X1 U1779 (.ZN(n2030), 
	.A3(n2031), 
	.A2(n200), 
	.A1(n753));
   NAND4_X1 U1780 (.ZN(n2031), 
	.A4(n16656), 
	.A3(FE_OFN15_n16671), 
	.A2(n2027), 
	.A1(n2032));
   OAI22_X1 U1781 (.ZN(U691_Z_0), 
	.B2(n2035), 
	.B1(n2034), 
	.A2(n2033), 
	.A1(n4968));
   AOI21_X1 U1782 (.ZN(n2034), 
	.B2(n2037), 
	.B1(n2036), 
	.A(n2038));
   OAI33_X1 U1783 (.ZN(n2038), 
	.B3(n16794), 
	.B2(n5026), 
	.B1(n2039), 
	.A3(n16847), 
	.A2(n4967), 
	.A1(n851));
   NAND2_X1 U1784 (.ZN(n2039), 
	.A2(n855), 
	.A1(n4967));
   INV_X1 U1785 (.ZN(n855), 
	.A(n1178));
   NAND2_X1 U1786 (.ZN(n1178), 
	.A2(FE_OFN90_n16849), 
	.A1(n527));
   OAI21_X1 U1787 (.ZN(n2037), 
	.B2(n753), 
	.B1(n5233), 
	.A(n5055));
   OAI221_X1 U1788 (.ZN(n2036), 
	.C2(n16734), 
	.C1(n16828), 
	.B2(n640), 
	.B1(n16847), 
	.A(n2040));
   NOR3_X1 U1789 (.ZN(n2040), 
	.A3(n799), 
	.A2(n2042), 
	.A1(n2041));
   AOI21_X1 U1790 (.ZN(n2041), 
	.B2(n17096), 
	.B1(n451), 
	.A(n16851));
   INV_X1 U1791 (.ZN(n2033), 
	.A(n2035));
   OAI21_X1 U1792 (.ZN(n2035), 
	.B2(n2044), 
	.B1(n2043), 
	.A(n17122));
   OAI221_X1 U1793 (.ZN(n2044), 
	.C2(n713), 
	.C1(n1857), 
	.B2(n522), 
	.B1(n1023), 
	.A(n2045));
   AOI22_X1 U1794 (.ZN(n2045), 
	.B2(n528), 
	.B1(n534), 
	.A2(n565), 
	.A1(n785));
   INV_X1 U1795 (.ZN(n534), 
	.A(n1230));
   NAND2_X1 U1796 (.ZN(n522), 
	.A2(FE_OFN89_n16849), 
	.A1(n528));
   NAND4_X1 U1797 (.ZN(n2043), 
	.A4(n2048), 
	.A3(n2047), 
	.A2(n738), 
	.A1(n2046));
   AOI22_X1 U1798 (.ZN(n2048), 
	.B2(n16734), 
	.B1(n1472), 
	.A2(n17097), 
	.A1(n546));
   NOR2_X1 U1799 (.ZN(n1472), 
	.A2(n17096), 
	.A1(n594));
   NOR2_X1 U1800 (.ZN(n546), 
	.A2(n16859), 
	.A1(n1217));
   NAND3_X1 U1801 (.ZN(n2047), 
	.A3(n728), 
	.A2(n16824), 
	.A1(n527));
   NAND3_X1 U1802 (.ZN(n2046), 
	.A3(n2049), 
	.A2(n1574), 
	.A1(n1097));
   OAI22_X1 U1803 (.ZN(U687_Z_0), 
	.B2(n17005), 
	.B1(FE_OFN128_n1809), 
	.A2(n17001), 
	.A1(FE_PHN2468_n5260));
   OAI22_X1 U1804 (.ZN(U686_Z_0), 
	.B2(n17005), 
	.B1(n1807), 
	.A2(n17001), 
	.A1(FE_PHN2596_n5261));
   OAI22_X1 U1805 (.ZN(U685_Z_0), 
	.B2(n17005), 
	.B1(n1808), 
	.A2(n17001), 
	.A1(FE_PHN2446_n5262));
   OAI22_X1 U1806 (.ZN(U684_Z_0), 
	.B2(n17000), 
	.B1(FE_OFN128_n1809), 
	.A2(n16996), 
	.A1(FE_PHN2546_n5018));
   INV_X2 U1808 (.ZN(n2056), 
	.A(n39));
   AOI221_X1 U1809 (.ZN(n39), 
	.C2(n2002), 
	.C1(n2058), 
	.B2(n2008), 
	.B1(FE_PSN5239_n2057), 
	.A(n2059));
   INV_X2 U1810 (.ZN(n2059), 
	.A(n2060));
   AOI221_X1 U1811 (.ZN(n2060), 
	.C2(n2062), 
	.C1(n2004), 
	.B2(n2061), 
	.B1(n2011), 
	.A(n2012));
   OAI22_X1 U1812 (.ZN(U683_Z_0), 
	.B2(n17000), 
	.B1(n1807), 
	.A2(n16996), 
	.A1(n4994));
   AOI221_X1 U1814 (.ZN(n76), 
	.C2(n2069), 
	.C1(n2068), 
	.B2(n2067), 
	.B1(n2066), 
	.A(n2070));
   INV_X2 U1815 (.ZN(n2070), 
	.A(n2071));
   AOI221_X1 U1816 (.ZN(n2071), 
	.C2(n2075), 
	.C1(n2074), 
	.B2(n2073), 
	.B1(n2072), 
	.A(n2076));
   OAI22_X1 U1817 (.ZN(U682_Z_0), 
	.B2(n17000), 
	.B1(n1808), 
	.A2(n16996), 
	.A1(FE_PHN2751_n4969));
   OAI22_X1 U1819 (.ZN(U681_Z_0), 
	.B2(n17005), 
	.B1(FE_OFN124_n2079), 
	.A2(n17001), 
	.A1(FE_PHN2639_n5643));
   OAI22_X1 U1820 (.ZN(U680_Z_0), 
	.B2(n17000), 
	.B1(FE_OFN124_n2079), 
	.A2(n16996), 
	.A1(n5642));
   OAI22_X1 U1821 (.ZN(U679_Z_0), 
	.B2(n17042), 
	.B1(FE_OFN124_n2079), 
	.A2(n17038), 
	.A1(FE_PHN2757_n5641));
   OAI22_X1 U1822 (.ZN(U678_Z_0), 
	.B2(n17037), 
	.B1(FE_OFN124_n2079), 
	.A2(n17033), 
	.A1(FE_PHN2556_n5640));
   OAI22_X1 U1823 (.ZN(U677_Z_0), 
	.B2(n17031), 
	.B1(FE_OFN124_n2079), 
	.A2(n17028), 
	.A1(n5082));
   OAI22_X1 U1824 (.ZN(U676_Z_0), 
	.B2(n17027), 
	.B1(FE_OFN124_n2079), 
	.A2(n17023), 
	.A1(FE_PHN2762_n5174));
   OAI22_X1 U1825 (.ZN(U675_Z_0), 
	.B2(n17022), 
	.B1(FE_OFN124_n2079), 
	.A2(n17018), 
	.A1(FE_PHN2589_n5081));
   OAI22_X1 U1826 (.ZN(U674_Z_0), 
	.B2(n17017), 
	.B1(FE_OFN124_n2079), 
	.A2(n17013), 
	.A1(FE_PHN2631_n5203));
   OAI22_X1 U1827 (.ZN(U673_Z_0), 
	.B2(n17046), 
	.B1(FE_OFN124_n2079), 
	.A2(n17043), 
	.A1(n5310));
   OAI22_X1 U1828 (.ZN(U672_Z_0), 
	.B2(n17052), 
	.B1(FE_OFN124_n2079), 
	.A2(n17048), 
	.A1(FE_PHN2535_n5339));
   OAI22_X1 U1829 (.ZN(U671_Z_0), 
	.B2(n17057), 
	.B1(FE_OFN124_n2079), 
	.A2(n17053), 
	.A1(FE_PHN2559_n5368));
   OAI22_X1 U1830 (.ZN(U670_Z_0), 
	.B2(n17062), 
	.B1(FE_OFN124_n2079), 
	.A2(n17058), 
	.A1(FE_PHN2715_n5397));
   OAI22_X1 U1831 (.ZN(U669_Z_0), 
	.B2(n17067), 
	.B1(FE_OFN124_n2079), 
	.A2(n17063), 
	.A1(FE_PHN2745_n5426));
   OAI22_X1 U1832 (.ZN(U668_Z_0), 
	.B2(n17071), 
	.B1(FE_OFN124_n2079), 
	.A2(n17068), 
	.A1(FE_PHN2760_n5455));
   OAI22_X1 U1833 (.ZN(U667_Z_0), 
	.B2(n17077), 
	.B1(FE_OFN124_n2079), 
	.A2(n17074), 
	.A1(n5080));
   OAI22_X1 U1834 (.ZN(U666_Z_0), 
	.B2(n17082), 
	.B1(FE_OFN124_n2079), 
	.A2(n17078), 
	.A1(FE_PHN2570_n5479));
   INV_X1 U1836 (.ZN(n2081), 
	.A(n2082));
   AOI221_X1 U1837 (.ZN(n2082), 
	.C2(FE_OFN2_n2015), 
	.C1(add_2073_SUM_31_), 
	.B2(n2083), 
	.B1(n17008), 
	.A(n2084));
   OAI22_X1 U1838 (.ZN(U665_Z_0), 
	.B2(n2087), 
	.B1(n2086), 
	.A2(n2085), 
	.A1(n4954));
   AOI222_X1 U1839 (.ZN(n2086), 
	.C2(n117), 
	.C1(n86), 
	.B2(n84), 
	.B1(n1528), 
	.A2(n2083), 
	.A1(n88));
   OAI221_X1 U1840 (.ZN(n117), 
	.C2(n2091), 
	.C1(n2090), 
	.B2(n2089), 
	.B1(n2088), 
	.A(n2092));
   AOI221_X1 U1841 (.ZN(n2092), 
	.C2(n2094), 
	.C1(n2067), 
	.B2(n2093), 
	.B1(n2074), 
	.A(n2076));
   INV_X1 U1842 (.ZN(n1528), 
	.A(n2095));
   OAI22_X1 U1843 (.ZN(n2095), 
	.B2(n1759), 
	.B1(n2097), 
	.A2(n2096), 
	.A1(n4947));
   NOR4_X1 U1844 (.ZN(n2097), 
	.A4(n2101), 
	.A3(n2100), 
	.A2(n2099), 
	.A1(n2098));
   NAND4_X1 U1845 (.ZN(n2101), 
	.A4(n2105), 
	.A3(n2104), 
	.A2(n2103), 
	.A1(n2102));
   AND4_X1 U1846 (.ZN(n2105), 
	.A4(n2109), 
	.A3(n2108), 
	.A2(n2107), 
	.A1(n2106));
   INV_X1 U1847 (.ZN(n2108), 
	.A(n2110));
   AND2_X1 U1848 (.ZN(n2106), 
	.A2(n2112), 
	.A1(n2111));
   AND3_X1 U1849 (.ZN(n2104), 
	.A3(n2115), 
	.A2(n2114), 
	.A1(n2113));
   NAND4_X1 U1850 (.ZN(n2100), 
	.A4(n2118), 
	.A3(n2117), 
	.A2(n2063), 
	.A1(n2116));
   AOI211_X1 U1851 (.ZN(n2118), 
	.C2(n2120), 
	.C1(n16994), 
	.B(n2080), 
	.A(n2121));
   OAI221_X1 U1852 (.ZN(n2080), 
	.C2(n2123), 
	.C1(n4954), 
	.B2(n2122), 
	.B1(n1677), 
	.A(n2124));
   INV_X1 U1853 (.ZN(n2123), 
	.A(n2125));
   AOI22_X1 U1854 (.ZN(n2122), 
	.B2(n2128), 
	.B1(n2127), 
	.A2(n2126), 
	.A1(U180_Z_0));
   INV_X1 U1855 (.ZN(n2128), 
	.A(U180_Z_0));
   OAI221_X1 U1856 (.ZN(n2121), 
	.C2(n2132), 
	.C1(n2131), 
	.B2(n2130), 
	.B1(n16992), 
	.A(n2133));
   OAI21_X1 U1857 (.ZN(n2133), 
	.B2(n2135), 
	.B1(n2134), 
	.A(FE_OFN208_n2015));
   NAND4_X1 U1858 (.ZN(n2135), 
	.A4(n2139), 
	.A3(n2138), 
	.A2(n2137), 
	.A1(n2136));
   NOR4_X1 U1859 (.ZN(n2139), 
	.A4(n16719), 
	.A3(n16653), 
	.A2(n16679), 
	.A1(n16658));
   NOR3_X1 U1860 (.ZN(n2138), 
	.A3(n16672), 
	.A2(add_2073_SUM_1_), 
	.A1(n16710));
   INV_X1 U1861 (.ZN(n2137), 
	.A(n16711));
   INV_X1 U1862 (.ZN(n2136), 
	.A(n16715));
   NAND4_X1 U1863 (.ZN(n2134), 
	.A4(n2142), 
	.A3(n2141), 
	.A2(n2140), 
	.A1(n1655));
   NOR3_X1 U1864 (.ZN(n2142), 
	.A3(n16663), 
	.A2(add_2073_SUM_31_), 
	.A1(n2143));
   OR3_X1 U1865 (.ZN(n2143), 
	.A3(n16682), 
	.A2(n16722), 
	.A1(add_2073_SUM_7_));
   NOR3_X1 U1866 (.ZN(n2141), 
	.A3(n16702), 
	.A2(n16655), 
	.A1(n16668));
   INV_X1 U1867 (.ZN(n2140), 
	.A(n16706));
   INV_X1 U1868 (.ZN(n1655), 
	.A(n16709));
   AOI211_X1 U1869 (.ZN(n2132), 
	.C2(n2144), 
	.C1(n5818), 
	.B(n2146), 
	.A(n2145));
   INV_X1 U1870 (.ZN(n2146), 
	.A(n2147));
   AOI22_X1 U1871 (.ZN(n2147), 
	.B2(n5807), 
	.B1(n1665), 
	.A2(n5819), 
	.A1(n2148));
   OAI221_X1 U1872 (.ZN(n2145), 
	.C2(n2150), 
	.C1(n1691), 
	.B2(n2149), 
	.B1(n1654), 
	.A(n2151));
   AOI22_X1 U1873 (.ZN(n2151), 
	.B2(n1651), 
	.B1(n5815), 
	.A2(n1645), 
	.A1(n4952));
   AOI211_X1 U1874 (.ZN(n2130), 
	.C2(n2144), 
	.C1(n2152), 
	.B(n2154), 
	.A(n2153));
   OAI22_X1 U1875 (.ZN(n2154), 
	.B2(n5807), 
	.B1(n1694), 
	.A2(n5819), 
	.A1(n1625));
   OAI221_X1 U1876 (.ZN(n2153), 
	.C2(n5815), 
	.C1(n1687), 
	.B2(n4952), 
	.B1(n1682), 
	.A(n2155));
   AOI22_X1 U1877 (.ZN(n2155), 
	.B2(n1658), 
	.B1(n2150), 
	.A2(n2156), 
	.A1(n2149));
   INV_X1 U1878 (.ZN(n2150), 
	.A(n5811));
   INV_X1 U1879 (.ZN(n2149), 
	.A(n5813));
   INV_X1 U1880 (.ZN(n2152), 
	.A(n5818));
   NAND4_X1 U1881 (.ZN(n2120), 
	.A4(n2160), 
	.A3(n2159), 
	.A2(n2158), 
	.A1(n2157));
   AOI222_X1 U1882 (.ZN(n2160), 
	.C2(n5817), 
	.C1(n1630), 
	.B2(n4952), 
	.B1(n1682), 
	.A2(n5816), 
	.A1(n1686));
   INV_X1 U1883 (.ZN(n1630), 
	.A(n2161));
   AOI222_X1 U1884 (.ZN(n2159), 
	.C2(n5814), 
	.C1(n1688), 
	.B2(n5815), 
	.B1(n1687), 
	.A2(n5813), 
	.A1(n1654));
   AOI222_X1 U1885 (.ZN(n2158), 
	.C2(n5811), 
	.C1(n1691), 
	.B2(n5812), 
	.B1(n1690), 
	.A2(n5810), 
	.A1(n1692));
   AOI222_X1 U1886 (.ZN(n2157), 
	.C2(n5819), 
	.C1(n1625), 
	.B2(n5807), 
	.B1(n1694), 
	.A2(n5818), 
	.A1(n1661));
   NOR3_X1 U1887 (.ZN(n2117), 
	.A3(n2017), 
	.A2(n2054), 
	.A1(n2001));
   OAI221_X1 U1888 (.ZN(n2017), 
	.C2(n2164), 
	.C1(n186), 
	.B2(n2163), 
	.B1(n2162), 
	.A(n2165));
   NOR3_X1 U1889 (.ZN(n2165), 
	.A3(n2167), 
	.A2(n2055), 
	.A1(n2166));
   NOR4_X1 U1890 (.ZN(n2167), 
	.A4(n2168), 
	.A3(n1045), 
	.A2(n16656), 
	.A1(n16810));
   NOR3_X1 U1891 (.ZN(n2166), 
	.A3(n1689), 
	.A2(n16992), 
	.A1(add_2082_B_1_));
   INV_X1 U1892 (.ZN(n2163), 
	.A(add_2082_B_1_));
   XOR2_X1 U1893 (.Z(add_2082_B_1_), 
	.B(n2170), 
	.A(n2169));
   AOI22_X1 U1894 (.ZN(n2170), 
	.B2(n2173), 
	.B1(n2172), 
	.A2(n1354), 
	.A1(n16988));
   AOI22_X2 U1895 (.ZN(n2162), 
	.B2(n2126), 
	.B1(n2174), 
	.A2(n16994), 
	.A1(n1689));
   INV_X4 U1896 (.ZN(n1689), 
	.A(n2174));
   NAND2_X4 U1897 (.ZN(n2174), 
	.A2(n2176), 
	.A1(n2175));
   AOI221_X2 U1898 (.ZN(n2176), 
	.C2(vis_r14_o[0]), 
	.C1(n16984), 
	.B2(vis_r11_o[0]), 
	.B1(n16985), 
	.A(n2181));
   OAI22_X1 U1899 (.ZN(n2181), 
	.B2(FE_PSN5237_n2184), 
	.B1(n2183), 
	.A2(n2182), 
	.A1(n5267));
   AOI221_X2 U1901 (.ZN(n2175), 
	.C2(n2188), 
	.C1(n16976), 
	.B2(vis_r9_o[0]), 
	.B1(n16979), 
	.A(n2189));
   OAI22_X1 U1902 (.ZN(n2189), 
	.B2(n2191), 
	.B1(n5338), 
	.A2(n2190), 
	.A1(n5396));
   OAI211_X1 U1903 (.ZN(n2054), 
	.C2(n2193), 
	.C1(n2192), 
	.B(n2195), 
	.A(n2194));
   AOI22_X1 U1904 (.ZN(n2195), 
	.B2(FE_OFN2_n2015), 
	.B1(n16726), 
	.A2(n2196), 
	.A1(n17008));
   NAND3_X1 U1905 (.ZN(n2194), 
	.A3(n2193), 
	.A2(n2127), 
	.A1(n1627));
   INV_X1 U1906 (.ZN(n2193), 
	.A(n5821));
   XOR2_X1 U1907 (.Z(n5821), 
	.B(n2197), 
	.A(n16990));
   AOI221_X1 U1908 (.ZN(n2197), 
	.C2(n2196), 
	.C1(n16988), 
	.B2(n16674), 
	.B1(n2198), 
	.A(n2199));
   OAI22_X1 U1909 (.ZN(n2199), 
	.B2(n2201), 
	.B1(n5258), 
	.A2(n2200), 
	.A1(n5256));
   AOI22_X1 U1910 (.ZN(n2192), 
	.B2(n2126), 
	.B1(n1627), 
	.A2(n16994), 
	.A1(n1672));
   INV_X1 U1911 (.ZN(n1672), 
	.A(n1627));
   NAND4_X1 U1912 (.ZN(n1627), 
	.A4(n2205), 
	.A3(n2204), 
	.A2(n2203), 
	.A1(n2202));
   AOI222_X1 U1913 (.ZN(n2205), 
	.C2(vis_psp_o[5]), 
	.C1(n16968), 
	.B2(n2209), 
	.B1(n16972), 
	.A2(vis_msp_o[5]), 
	.A1(n16973));
   AOI222_X1 U1914 (.ZN(n2204), 
	.C2(vis_r11_o[7]), 
	.C1(n16985), 
	.B2(vis_r12_o[7]), 
	.B1(FE_OFN109_n16964), 
	.A2(vis_r14_o[7]), 
	.A1(n16982));
   AOI222_X1 U1915 (.ZN(n2203), 
	.C2(vis_r8_o[7]), 
	.C1(n16959), 
	.B2(vis_r10_o[7]), 
	.B1(n16962), 
	.A2(vis_r9_o[7]), 
	.A1(n16979));
   AOI22_X1 U1916 (.ZN(n2202), 
	.B2(n1152), 
	.B1(n16955), 
	.A2(n2221), 
	.A1(n16976));
   OAI211_X1 U1917 (.ZN(n2001), 
	.C2(n2224), 
	.C1(n2223), 
	.B(n2226), 
	.A(n2225));
   AOI222_X1 U1918 (.ZN(n2226), 
	.C2(n2028), 
	.C1(n17008), 
	.B2(vis_ipsr_o[1]), 
	.B1(n2227), 
	.A2(FE_OFN2_n2015), 
	.A1(n16732));
   AOI21_X1 U1919 (.ZN(n2225), 
	.B2(n2224), 
	.B1(n2228), 
	.A(n2229));
   NOR4_X1 U1920 (.ZN(n2229), 
	.A4(n2168), 
	.A3(n16810), 
	.A2(n5055), 
	.A1(n16809));
   NOR2_X1 U1921 (.ZN(n2228), 
	.A2(n1679), 
	.A1(n16992));
   INV_X1 U1922 (.ZN(n2224), 
	.A(n5822));
   XOR2_X1 U1923 (.Z(n5822), 
	.B(n2230), 
	.A(n16990));
   AOI222_X1 U1924 (.ZN(n2230), 
	.C2(n2173), 
	.C1(n2231), 
	.B2(n451), 
	.B1(n2198), 
	.A2(n2028), 
	.A1(n16988));
   AOI22_X1 U1925 (.ZN(n2223), 
	.B2(n2126), 
	.B1(n2232), 
	.A2(n16994), 
	.A1(n1679));
   INV_X4 U1926 (.ZN(n1679), 
	.A(n2232));
   AOI221_X1 U1927 (.ZN(n2063), 
	.C2(n2125), 
	.C1(vis_apsr_o[0]), 
	.B2(n17008), 
	.B1(n89), 
	.A(n2055));
   INV_X1 U1928 (.ZN(n2116), 
	.A(n2233));
   NAND4_X1 U1929 (.ZN(n2099), 
	.A4(n2237), 
	.A3(n2236), 
	.A2(n2235), 
	.A1(n2234));
   NOR3_X1 U1930 (.ZN(n2237), 
	.A3(n2240), 
	.A2(n2239), 
	.A1(n2238));
   AOI21_X1 U1931 (.ZN(n2240), 
	.B2(n2242), 
	.B1(n2241), 
	.A(n2243));
   NOR4_X1 U1932 (.ZN(n2242), 
	.A4(n2247), 
	.A3(n2246), 
	.A2(n2245), 
	.A1(n2244));
   OR3_X1 U1933 (.ZN(n2245), 
	.A3(n2249), 
	.A2(n2248), 
	.A1(n2083));
   OR4_X1 U1934 (.ZN(n2244), 
	.A4(n2252), 
	.A3(n17), 
	.A2(n2251), 
	.A1(n2250));
   OR2_X1 U1935 (.ZN(n2252), 
	.A2(n2254), 
	.A1(n2253));
   NOR4_X1 U1936 (.ZN(n2241), 
	.A4(n2258), 
	.A3(n2257), 
	.A2(n2256), 
	.A1(n2255));
   OR3_X1 U1937 (.ZN(n2256), 
	.A3(n21), 
	.A2(n20), 
	.A1(n22));
   OR4_X1 U1938 (.ZN(n2255), 
	.A4(n2261), 
	.A3(n1354), 
	.A2(n2260), 
	.A1(n2259));
   INV_X1 U1939 (.ZN(n2239), 
	.A(n2064));
   NAND2_X1 U1940 (.ZN(n2064), 
	.A2(FE_OFN2_n2015), 
	.A1(n16695));
   NAND3_X1 U1941 (.ZN(n2238), 
	.A3(n2263), 
	.A2(n2065), 
	.A1(n2262));
   OAI221_X1 U1942 (.ZN(n2065), 
	.C2(n1832), 
	.C1(n16994), 
	.B2(n2264), 
	.B1(U189_Z_0), 
	.A(n2265));
   NAND3_X1 U1943 (.ZN(n2265), 
	.A3(n2131), 
	.A2(n1832), 
	.A1(U189_Z_0));
   NOR2_X1 U1944 (.ZN(n2264), 
	.A2(n16992), 
	.A1(n1680));
   INV_X1 U1945 (.ZN(n1680), 
	.A(FE_OFN504_n1832));
   NAND4_X1 U1946 (.ZN(n1832), 
	.A4(n2269), 
	.A3(n2268), 
	.A2(n2267), 
	.A1(n2266));
   AOI222_X1 U1947 (.ZN(n2269), 
	.C2(vis_psp_o[26]), 
	.C1(n16967), 
	.B2(n2271), 
	.B1(n16972), 
	.A2(vis_msp_o[26]), 
	.A1(n16973));
   AOI222_X1 U1949 (.ZN(n2268), 
	.C2(vis_r11_o[28]), 
	.C1(n16985), 
	.B2(vis_r12_o[28]), 
	.B1(FE_OFN109_n16964), 
	.A2(vis_r14_o[28]), 
	.A1(n16982));
   AOI222_X1 U1952 (.ZN(n2267), 
	.C2(vis_r8_o[28]), 
	.C1(n16958), 
	.B2(vis_r10_o[28]), 
	.B1(n16961), 
	.A2(vis_r9_o[28]), 
	.A1(n16979));
   AOI22_X1 U1954 (.ZN(n2266), 
	.B2(n2280), 
	.B1(n16954), 
	.A2(n2279), 
	.A1(n16976));
   AND3_X1 U1955 (.ZN(n2236), 
	.A3(n2283), 
	.A2(n2282), 
	.A1(n2281));
   NAND4_X1 U1956 (.ZN(n2098), 
	.A4(n2287), 
	.A3(n2286), 
	.A2(n2285), 
	.A1(n2284));
   NOR4_X1 U1957 (.ZN(n2287), 
	.A4(n2290), 
	.A3(n2289), 
	.A2(n2084), 
	.A1(n2288));
   INV_X1 U1958 (.ZN(n2290), 
	.A(n2291));
   AND3_X1 U1959 (.ZN(n2084), 
	.A3(n1677), 
	.A2(U180_Z_0), 
	.A1(n16994));
   AND4_X1 U1960 (.ZN(n1677), 
	.A4(n2295), 
	.A3(n2294), 
	.A2(n2293), 
	.A1(n2292));
   AOI222_X1 U1961 (.ZN(n2295), 
	.C2(vis_psp_o[28]), 
	.C1(n16967), 
	.B2(n2297), 
	.B1(n16972), 
	.A2(vis_msp_o[28]), 
	.A1(n16973));
   AOI222_X1 U1963 (.ZN(n2294), 
	.C2(vis_r11_o[30]), 
	.C1(n16985), 
	.B2(vis_r12_o[30]), 
	.B1(n16965), 
	.A2(vis_r14_o[30]), 
	.A1(n16982));
   AOI222_X1 U1966 (.ZN(n2293), 
	.C2(vis_r8_o[30]), 
	.C1(n16958), 
	.B2(vis_r10_o[30]), 
	.B1(n16961), 
	.A2(vis_r9_o[30]), 
	.A1(n16979));
   AOI22_X1 U1968 (.ZN(n2292), 
	.B2(n881), 
	.B1(n16954), 
	.A2(n874), 
	.A1(n16976));
   NAND3_X1 U1969 (.ZN(n2288), 
	.A3(n2307), 
	.A2(n2306), 
	.A1(n2305));
   NOR3_X1 U1970 (.ZN(n2286), 
	.A3(n2310), 
	.A2(n2309), 
	.A1(n2308));
   AOI221_X1 U1971 (.ZN(n2096), 
	.C2(n2314), 
	.C1(n2313), 
	.B2(n2312), 
	.B1(n2311), 
	.A(n2315));
   OAI221_X1 U1972 (.ZN(n2315), 
	.C2(n2319), 
	.C1(n2318), 
	.B2(n2317), 
	.B1(n2316), 
	.A(n2320));
   OAI33_X1 U1973 (.ZN(n2320), 
	.B3(n2326), 
	.B2(n2325), 
	.B1(n2324), 
	.A3(n2323), 
	.A2(n2322), 
	.A1(n2321));
   NAND3_X1 U1974 (.ZN(n2324), 
	.A3(n2327), 
	.A2(n1789), 
	.A1(n1781));
   OAI33_X1 U1975 (.ZN(n2327), 
	.B3(n2333), 
	.B2(n2332), 
	.B1(n2331), 
	.A3(n2330), 
	.A2(n2329), 
	.A1(n2328));
   OR3_X1 U1976 (.ZN(n2331), 
	.A3(n2336), 
	.A2(n16788), 
	.A1(n2334));
   OR3_X1 U1977 (.ZN(n2328), 
	.A3(n2339), 
	.A2(FE_OFN529_n2338), 
	.A1(n2337));
   AOI21_X1 U1978 (.ZN(n2319), 
	.B2(n2341), 
	.B1(n2340), 
	.A(n2342));
   NOR3_X1 U1979 (.ZN(n2318), 
	.A3(n2345), 
	.A2(n2344), 
	.A1(n2343));
   NAND3_X1 U1980 (.ZN(n2343), 
	.A3(n2347), 
	.A2(n2346), 
	.A1(n1779));
   OAI33_X1 U1981 (.ZN(n2347), 
	.B3(n2353), 
	.B2(n2352), 
	.B1(n2351), 
	.A3(n2350), 
	.A2(n2349), 
	.A1(n2348));
   OR3_X1 U1982 (.ZN(n2351), 
	.A3(n2355), 
	.A2(n16788), 
	.A1(n2354));
   OR3_X1 U1983 (.ZN(n2348), 
	.A3(n2357), 
	.A2(n2356), 
	.A1(n2337));
   NOR4_X1 U1984 (.ZN(n2317), 
	.A4(n2360), 
	.A3(n2359), 
	.A2(n2340), 
	.A1(n2358));
   NOR4_X1 U1985 (.ZN(n2316), 
	.A4(n2364), 
	.A3(n2363), 
	.A2(n2362), 
	.A1(n2361));
   OAI22_X1 U1986 (.ZN(n2362), 
	.B2(n2368), 
	.B1(n2367), 
	.A2(n2366), 
	.A1(n2365));
   NOR2_X1 U1987 (.ZN(n2367), 
	.A2(n2369), 
	.A1(n2337));
   INV_X1 U1988 (.ZN(n2366), 
	.A(n2370));
   INV_X1 U1989 (.ZN(n2365), 
	.A(n2371));
   NAND4_X1 U1990 (.ZN(n2361), 
	.A4(n2375), 
	.A3(n2374), 
	.A2(n2373), 
	.A1(n2372));
   OAI21_X1 U1991 (.ZN(n2314), 
	.B2(n2342), 
	.B1(n2340), 
	.A(n2376));
   INV_X1 U1992 (.ZN(n2342), 
	.A(n2377));
   NAND4_X1 U1993 (.ZN(n2312), 
	.A4(n2381), 
	.A3(n2380), 
	.A2(n2379), 
	.A1(n2378));
   OAI33_X1 U1994 (.ZN(n2381), 
	.B3(n2353), 
	.B2(n2352), 
	.B1(n2383), 
	.A3(n2330), 
	.A2(FE_OFN523_n2329), 
	.A1(n2382));
   OR3_X1 U1995 (.ZN(n2383), 
	.A3(n2385), 
	.A2(n2384), 
	.A1(n2337));
   OR3_X1 U1996 (.ZN(n2382), 
	.A3(n2387), 
	.A2(n16788), 
	.A1(n2386));
   AND2_X1 U1997 (.ZN(n2380), 
	.A2(n1772), 
	.A1(n1791));
   INV_X1 U1998 (.ZN(n2379), 
	.A(n2388));
   OAI21_X1 U1999 (.ZN(n2311), 
	.B2(n2390), 
	.B1(n2389), 
	.A(n2377));
   OAI22_X1 U2000 (.ZN(U664_Z_0), 
	.B2(n17005), 
	.B1(FE_OFN132_n2391), 
	.A2(n17001), 
	.A1(FE_PHN2577_n5079));
   OAI22_X1 U2001 (.ZN(U663_Z_0), 
	.B2(n17000), 
	.B1(FE_OFN132_n2391), 
	.A2(n16996), 
	.A1(n5078));
   OAI22_X1 U2002 (.ZN(U662_Z_0), 
	.B2(n17042), 
	.B1(FE_OFN132_n2391), 
	.A2(n17038), 
	.A1(FE_PHN2650_n5289));
   OAI22_X1 U2003 (.ZN(U661_Z_0), 
	.B2(n17037), 
	.B1(FE_OFN132_n2391), 
	.A2(n17033), 
	.A1(FE_PHN2551_n5268));
   OAI22_X1 U2004 (.ZN(U660_Z_0), 
	.B2(n17031), 
	.B1(FE_OFN132_n2391), 
	.A2(n17028), 
	.A1(n5077));
   OAI22_X1 U2005 (.ZN(U659_Z_0), 
	.B2(n17027), 
	.B1(FE_OFN132_n2391), 
	.A2(n17023), 
	.A1(FE_PHN2687_n5175));
   OAI22_X1 U2006 (.ZN(U658_Z_0), 
	.B2(n17022), 
	.B1(FE_OFN132_n2391), 
	.A2(n17018), 
	.A1(FE_PHN2607_n5076));
   OAI22_X1 U2007 (.ZN(U657_Z_0), 
	.B2(n17017), 
	.B1(FE_OFN132_n2391), 
	.A2(n17013), 
	.A1(FE_PHN2437_n5204));
   OAI22_X1 U2008 (.ZN(U656_Z_0), 
	.B2(n17046), 
	.B1(FE_OFN132_n2391), 
	.A2(n17043), 
	.A1(n5311));
   OAI22_X1 U2009 (.ZN(U655_Z_0), 
	.B2(n17052), 
	.B1(FE_OFN132_n2391), 
	.A2(n17048), 
	.A1(FE_PHN2439_n5340));
   OAI22_X1 U2010 (.ZN(U654_Z_0), 
	.B2(n17057), 
	.B1(FE_OFN132_n2391), 
	.A2(n17053), 
	.A1(FE_PHN2557_n5369));
   OAI22_X1 U2011 (.ZN(U653_Z_0), 
	.B2(n17062), 
	.B1(FE_OFN132_n2391), 
	.A2(n17058), 
	.A1(FE_PHN2692_n5398));
   OAI22_X1 U2012 (.ZN(U652_Z_0), 
	.B2(n17067), 
	.B1(FE_OFN132_n2391), 
	.A2(n17063), 
	.A1(FE_PHN2710_n5427));
   OAI22_X1 U2013 (.ZN(U651_Z_0), 
	.B2(n17071), 
	.B1(FE_OFN132_n2391), 
	.A2(n17068), 
	.A1(n5456));
   OAI22_X1 U2014 (.ZN(U650_Z_0), 
	.B2(n17077), 
	.B1(FE_OFN132_n2391), 
	.A2(n17074), 
	.A1(FE_PHN2778_n5075));
   OAI22_X1 U2015 (.ZN(U649_Z_0), 
	.B2(n17082), 
	.B1(FE_OFN132_n2391), 
	.A2(n17078), 
	.A1(FE_PHN2506_n5480));
   OAI211_X1 U2017 (.ZN(n2233), 
	.C2(n2393), 
	.C1(n2392), 
	.B(n2395), 
	.A(n2394));
   AOI222_X1 U2018 (.ZN(n2395), 
	.C2(FE_OFN2_n2015), 
	.C1(n16693), 
	.B2(n1755), 
	.B1(n17008), 
	.A2(vis_apsr_o[1]), 
	.A1(n2125));
   AOI21_X1 U2020 (.ZN(n2394), 
	.B2(n1870), 
	.B1(n2396), 
	.A(n2055));
   NOR2_X1 U2021 (.ZN(n2396), 
	.A2(n16992), 
	.A1(U158_Z_0));
   AOI22_X1 U2022 (.ZN(n2393), 
	.B2(n2126), 
	.B1(n1870), 
	.A2(n16994), 
	.A1(n1678));
   INV_X1 U2023 (.ZN(n1678), 
	.A(n1870));
   NAND4_X1 U2024 (.ZN(n1870), 
	.A4(n2400), 
	.A3(n2399), 
	.A2(n2398), 
	.A1(n2397));
   AOI222_X1 U2025 (.ZN(n2400), 
	.C2(vis_psp_o[27]), 
	.C1(n16967), 
	.B2(n2402), 
	.B1(n16972), 
	.A2(vis_msp_o[27]), 
	.A1(n16974));
   AOI222_X1 U2027 (.ZN(n2399), 
	.C2(vis_r11_o[29]), 
	.C1(n16985), 
	.B2(vis_r12_o[29]), 
	.B1(n16965), 
	.A2(vis_r14_o[29]), 
	.A1(n16982));
   AOI222_X1 U2030 (.ZN(n2398), 
	.C2(vis_r8_o[29]), 
	.C1(n16958), 
	.B2(vis_r10_o[29]), 
	.B1(n16961), 
	.A2(vis_r9_o[29]), 
	.A1(n16979));
   AOI22_X1 U2032 (.ZN(n2397), 
	.B2(n2279), 
	.B1(n16954), 
	.A2(n881), 
	.A1(n16976));
   INV_X1 U2035 (.ZN(n2392), 
	.A(U158_Z_0));
   INV_X1 U2036 (.ZN(n1754), 
	.A(FE_PHN768_n72));
   AOI221_X1 U2037 (.ZN(n72), 
	.C2(n2074), 
	.C1(n2411), 
	.B2(n2067), 
	.B1(n2410), 
	.A(n2412));
   INV_X2 U2038 (.ZN(n2412), 
	.A(n2413));
   AOI221_X1 U2039 (.ZN(n2413), 
	.C2(n2069), 
	.C1(FE_PHN748_n2415), 
	.B2(n2414), 
	.B1(n2072), 
	.A(n2076));
   OAI22_X1 U2040 (.ZN(U648_Z_0), 
	.B2(n17005), 
	.B1(FE_OFN126_n2416), 
	.A2(n17001), 
	.A1(FE_PHN2534_n5630));
   OAI22_X1 U2041 (.ZN(U647_Z_0), 
	.B2(n17000), 
	.B1(FE_OFN126_n2416), 
	.A2(n16996), 
	.A1(FE_PHN2630_n5629));
   OAI22_X1 U2042 (.ZN(U646_Z_0), 
	.B2(n17042), 
	.B1(FE_OFN126_n2416), 
	.A2(n17038), 
	.A1(n5628));
   OAI22_X1 U2043 (.ZN(U645_Z_0), 
	.B2(n17037), 
	.B1(FE_OFN126_n2416), 
	.A2(n17033), 
	.A1(FE_PHN2462_n5627));
   OAI22_X1 U2044 (.ZN(U644_Z_0), 
	.B2(n17031), 
	.B1(FE_OFN126_n2416), 
	.A2(n17028), 
	.A1(n5113));
   OAI22_X1 U2045 (.ZN(U643_Z_0), 
	.B2(n17027), 
	.B1(FE_OFN126_n2416), 
	.A2(n17023), 
	.A1(FE_PHN2633_n5176));
   OAI22_X1 U2046 (.ZN(U642_Z_0), 
	.B2(n17022), 
	.B1(FE_OFN126_n2416), 
	.A2(n17018), 
	.A1(FE_PHN2609_n5112));
   OAI22_X1 U2047 (.ZN(U641_Z_0), 
	.B2(n17017), 
	.B1(FE_OFN126_n2416), 
	.A2(n17013), 
	.A1(FE_PHN2616_n5205));
   OAI22_X1 U2048 (.ZN(U640_Z_0), 
	.B2(n17046), 
	.B1(FE_OFN126_n2416), 
	.A2(n17043), 
	.A1(FE_PHN2748_n5312));
   OAI22_X1 U2049 (.ZN(U639_Z_0), 
	.B2(n17052), 
	.B1(FE_OFN126_n2416), 
	.A2(n17048), 
	.A1(FE_PHN2450_n5341));
   OAI22_X1 U2050 (.ZN(U638_Z_0), 
	.B2(n17057), 
	.B1(FE_OFN126_n2416), 
	.A2(n17053), 
	.A1(FE_PHN2449_n5370));
   OAI22_X1 U2051 (.ZN(U637_Z_0), 
	.B2(n17062), 
	.B1(FE_OFN126_n2416), 
	.A2(n17058), 
	.A1(FE_PHN2657_n5399));
   OAI22_X1 U2052 (.ZN(U636_Z_0), 
	.B2(n17067), 
	.B1(FE_OFN126_n2416), 
	.A2(n17063), 
	.A1(FE_PHN2746_n5428));
   OAI22_X1 U2053 (.ZN(U635_Z_0), 
	.B2(n17071), 
	.B1(FE_OFN126_n2416), 
	.A2(n17068), 
	.A1(FE_PHN2801_n5457));
   OAI22_X1 U2054 (.ZN(U634_Z_0), 
	.B2(n17077), 
	.B1(FE_OFN126_n2416), 
	.A2(n17074), 
	.A1(n5111));
   OAI22_X1 U2055 (.ZN(U633_Z_0), 
	.B2(n17082), 
	.B1(FE_OFN126_n2416), 
	.A2(n17078), 
	.A1(FE_PHN2617_n5481));
   OAI221_X1 U2057 (.ZN(n99), 
	.C2(n2419), 
	.C1(n2089), 
	.B2(n2418), 
	.B1(n2417), 
	.A(n2420));
   AOI221_X1 U2058 (.ZN(n2420), 
	.C2(n2069), 
	.C1(n2422), 
	.B2(FE_PHN728_n2421), 
	.B1(n2074), 
	.A(n2076));
   OAI211_X1 U2059 (.ZN(n2110), 
	.C2(n2424), 
	.C1(n2423), 
	.B(n2426), 
	.A(n2425));
   AOI22_X1 U2060 (.ZN(n2426), 
	.B2(FE_OFN2_n2015), 
	.B1(n16698), 
	.A2(n2427), 
	.A1(n17008));
   NAND3_X1 U2061 (.ZN(n2425), 
	.A3(n1644), 
	.A2(n2423), 
	.A1(n2127));
   AOI22_X1 U2062 (.ZN(n2424), 
	.B2(n2126), 
	.B1(n1644), 
	.A2(n16994), 
	.A1(n1681));
   INV_X1 U2063 (.ZN(n1681), 
	.A(n1644));
   NAND4_X1 U2064 (.ZN(n1644), 
	.A4(n2431), 
	.A3(n2430), 
	.A2(n2429), 
	.A1(n2428));
   AOI222_X1 U2065 (.ZN(n2431), 
	.C2(vis_psp_o[25]), 
	.C1(n16967), 
	.B2(n2433), 
	.B1(n16972), 
	.A2(vis_msp_o[25]), 
	.A1(n16973));
   AOI222_X1 U2067 (.ZN(n2430), 
	.C2(vis_r11_o[27]), 
	.C1(n16985), 
	.B2(vis_r12_o[27]), 
	.B1(FE_OFN109_n16964), 
	.A2(vis_r14_o[27]), 
	.A1(n16982));
   AOI222_X1 U2070 (.ZN(n2429), 
	.C2(vis_r8_o[27]), 
	.C1(n16958), 
	.B2(vis_r10_o[27]), 
	.B1(n16961), 
	.A2(vis_r9_o[27]), 
	.A1(n16979));
   AOI22_X1 U2072 (.ZN(n2428), 
	.B2(n2441), 
	.B1(n16954), 
	.A2(n2280), 
	.A1(n16976));
   INV_X1 U2074 (.ZN(n2423), 
	.A(U175_Z_0));
   OAI22_X1 U2075 (.ZN(U632_Z_0), 
	.B2(n17005), 
	.B1(n2442), 
	.A2(n17001), 
	.A1(n4993));
   OAI22_X1 U2076 (.ZN(U631_Z_0), 
	.B2(n17000), 
	.B1(n2442), 
	.A2(n16996), 
	.A1(FE_PHN3624_n4992));
   OAI22_X1 U2077 (.ZN(U630_Z_0), 
	.B2(n17042), 
	.B1(n2442), 
	.A2(n17038), 
	.A1(n5290));
   OAI22_X1 U2078 (.ZN(U629_Z_0), 
	.B2(n17037), 
	.B1(n2442), 
	.A2(n17033), 
	.A1(FE_PHN3593_n5269));
   OAI22_X1 U2079 (.ZN(U628_Z_0), 
	.B2(n17031), 
	.B1(n2442), 
	.A2(n17028), 
	.A1(n4991));
   OAI22_X1 U2080 (.ZN(U627_Z_0), 
	.B2(n17027), 
	.B1(n2442), 
	.A2(n17023), 
	.A1(n5177));
   OAI22_X1 U2081 (.ZN(U626_Z_0), 
	.B2(n17022), 
	.B1(n2442), 
	.A2(n17018), 
	.A1(FE_PHN3584_n4990));
   OAI22_X1 U2082 (.ZN(U625_Z_0), 
	.B2(n17017), 
	.B1(n2442), 
	.A2(n17013), 
	.A1(FE_PHN3556_n5206));
   OAI22_X1 U2083 (.ZN(U624_Z_0), 
	.B2(n17046), 
	.B1(n2442), 
	.A2(n17043), 
	.A1(n5313));
   OAI22_X1 U2084 (.ZN(U623_Z_0), 
	.B2(n17052), 
	.B1(n2442), 
	.A2(n17048), 
	.A1(FE_PHN3567_n5342));
   OAI22_X1 U2085 (.ZN(U622_Z_0), 
	.B2(n17057), 
	.B1(n2442), 
	.A2(n17053), 
	.A1(FE_PHN3562_n5371));
   OAI22_X1 U2086 (.ZN(U621_Z_0), 
	.B2(n17062), 
	.B1(n2442), 
	.A2(n17058), 
	.A1(FE_PHN3629_n5400));
   OAI22_X1 U2087 (.ZN(U620_Z_0), 
	.B2(n17067), 
	.B1(n2442), 
	.A2(n17063), 
	.A1(FE_PHN3637_n5429));
   OAI22_X1 U2088 (.ZN(U619_Z_0), 
	.B2(n17071), 
	.B1(n2442), 
	.A2(n17068), 
	.A1(n5458));
   OAI22_X1 U2089 (.ZN(U618_Z_0), 
	.B2(n17077), 
	.B1(n2442), 
	.A2(n17074), 
	.A1(FE_PHN3633_n4989));
   OAI22_X1 U2090 (.ZN(U617_Z_0), 
	.B2(n17082), 
	.B1(n2442), 
	.A2(n17078), 
	.A1(FE_PHN3563_n5482));
   AOI221_X1 U2092 (.ZN(n2444), 
	.C2(FE_OFN2_n2015), 
	.C1(n16663), 
	.B2(n2260), 
	.B1(n17008), 
	.A(n2055));
   OAI221_X1 U2093 (.ZN(n2443), 
	.C2(n1645), 
	.C1(n16994), 
	.B2(n2445), 
	.B1(n4952), 
	.A(n2446));
   NAND3_X1 U2094 (.ZN(n2446), 
	.A3(n4952), 
	.A2(n1645), 
	.A1(n2131));
   NOR2_X1 U2095 (.ZN(n2445), 
	.A2(n16992), 
	.A1(n1682));
   INV_X1 U2096 (.ZN(n1682), 
	.A(n1645));
   NAND4_X2 U2097 (.ZN(n1645), 
	.A4(n2450), 
	.A3(n2449), 
	.A2(n2448), 
	.A1(n2447));
   AOI222_X1 U2098 (.ZN(n2450), 
	.C2(vis_psp_o[24]), 
	.C1(n16967), 
	.B2(n2452), 
	.B1(n16972), 
	.A2(vis_msp_o[24]), 
	.A1(n16973));
   AOI222_X1 U2100 (.ZN(n2449), 
	.C2(vis_r11_o[26]), 
	.C1(n16985), 
	.B2(vis_r12_o[26]), 
	.B1(FE_OFN109_n16964), 
	.A2(vis_r14_o[26]), 
	.A1(n16982));
   AOI222_X1 U2103 (.ZN(n2448), 
	.C2(vis_r8_o[26]), 
	.C1(n16958), 
	.B2(vis_r10_o[26]), 
	.B1(n16961), 
	.A2(vis_r9_o[26]), 
	.A1(n16980));
   AOI22_X1 U2105 (.ZN(n2447), 
	.B2(n2460), 
	.B1(n16954), 
	.A2(n2441), 
	.A1(n16976));
   INV_X1 U2108 (.ZN(n2463), 
	.A(n2260));
   AOI221_X1 U2109 (.ZN(n100), 
	.C2(n2074), 
	.C1(FE_PHN679_n2465), 
	.B2(n2069), 
	.B1(n2464), 
	.A(n2466));
   INV_X1 U2110 (.ZN(n2466), 
	.A(n2467));
   AOI221_X1 U2111 (.ZN(n2467), 
	.C2(n2067), 
	.C1(n2469), 
	.B2(n2072), 
	.B1(n2468), 
	.A(n2076));
   OAI22_X1 U2112 (.ZN(U614_Z_0), 
	.B2(n17005), 
	.B1(n2470), 
	.A2(n17001), 
	.A1(FE_PHN2445_n5016));
   OAI22_X1 U2113 (.ZN(U613_Z_0), 
	.B2(n17000), 
	.B1(n2470), 
	.A2(n16996), 
	.A1(FE_PHN2750_n5015));
   OAI22_X1 U2114 (.ZN(U612_Z_0), 
	.B2(n17042), 
	.B1(n2470), 
	.A2(n17038), 
	.A1(n5291));
   OAI22_X1 U2115 (.ZN(U611_Z_0), 
	.B2(n17037), 
	.B1(n2470), 
	.A2(n17033), 
	.A1(FE_PHN2613_n5270));
   OAI22_X1 U2116 (.ZN(U610_Z_0), 
	.B2(n17031), 
	.B1(n2470), 
	.A2(n17028), 
	.A1(n5014));
   OAI22_X1 U2117 (.ZN(U609_Z_0), 
	.B2(n17027), 
	.B1(n2470), 
	.A2(n17023), 
	.A1(FE_PHN2770_n5178));
   OAI22_X1 U2118 (.ZN(U608_Z_0), 
	.B2(n17022), 
	.B1(n2470), 
	.A2(n17018), 
	.A1(FE_PHN2627_n5013));
   OAI22_X1 U2119 (.ZN(U607_Z_0), 
	.B2(n17017), 
	.B1(n2470), 
	.A2(n17013), 
	.A1(FE_PHN2635_n5207));
   OAI22_X1 U2120 (.ZN(U606_Z_0), 
	.B2(n17046), 
	.B1(n2470), 
	.A2(n17043), 
	.A1(n5314));
   OAI22_X1 U2121 (.ZN(U605_Z_0), 
	.B2(n17052), 
	.B1(n2470), 
	.A2(n17048), 
	.A1(FE_PHN2603_n5343));
   OAI22_X1 U2122 (.ZN(U604_Z_0), 
	.B2(n17057), 
	.B1(n2470), 
	.A2(n17053), 
	.A1(FE_PHN2563_n5372));
   OAI22_X1 U2123 (.ZN(U603_Z_0), 
	.B2(n17062), 
	.B1(n2470), 
	.A2(n17058), 
	.A1(FE_PHN2695_n5401));
   OAI22_X1 U2124 (.ZN(U602_Z_0), 
	.B2(n17067), 
	.B1(n2470), 
	.A2(n17063), 
	.A1(FE_PHN2701_n5430));
   OAI22_X1 U2125 (.ZN(U601_Z_0), 
	.B2(n17071), 
	.B1(n2470), 
	.A2(n17068), 
	.A1(FE_PHN2707_n5459));
   OAI22_X1 U2126 (.ZN(U600_Z_0), 
	.B2(n17077), 
	.B1(n2470), 
	.A2(n17074), 
	.A1(FE_PHN2722_n5012));
   OAI22_X1 U2127 (.ZN(U599_Z_0), 
	.B2(n17082), 
	.B1(n2470), 
	.A2(n17078), 
	.A1(FE_PHN2622_n5483));
   AOI221_X1 U2129 (.ZN(n2471), 
	.C2(n2248), 
	.C1(n17008), 
	.B2(FE_OFN2_n2015), 
	.B1(n16655), 
	.A(n108));
   OAI221_X1 U2130 (.ZN(n108), 
	.C2(n2089), 
	.C1(n2473), 
	.B2(n2472), 
	.B1(n2417), 
	.A(n2474));
   AOI221_X1 U2131 (.ZN(n2474), 
	.C2(n2069), 
	.C1(n2005), 
	.B2(n2003), 
	.B1(n2074), 
	.A(n2076));
   NAND3_X1 U2132 (.ZN(n2234), 
	.A3(n1683), 
	.A2(n4951), 
	.A1(n16994));
   INV_X1 U2133 (.ZN(n1683), 
	.A(n1647));
   NAND2_X1 U2134 (.ZN(n2291), 
	.A2(n1647), 
	.A1(n2475));
   NAND4_X1 U2135 (.ZN(n1647), 
	.A4(n2479), 
	.A3(n2478), 
	.A2(n2477), 
	.A1(n2476));
   AOI222_X1 U2136 (.ZN(n2479), 
	.C2(vis_r9_o[25]), 
	.C1(n16979), 
	.B2(n16954), 
	.B1(n2481), 
	.A2(vis_r8_o[25]), 
	.A1(n16958));
   AOI222_X1 U2138 (.ZN(n2478), 
	.C2(vis_r14_o[25]), 
	.C1(n16984), 
	.B2(n2484), 
	.B1(n16972), 
	.A2(vis_r11_o[25]), 
	.A1(n16985));
   AOI222_X1 U2141 (.ZN(n2477), 
	.C2(vis_msp_o[23]), 
	.C1(n16975), 
	.B2(vis_r10_o[25]), 
	.B1(n16961), 
	.A2(vis_psp_o[23]), 
	.A1(n16967));
   AOI22_X1 U2143 (.ZN(n2476), 
	.B2(n2460), 
	.B1(n16976), 
	.A2(vis_r12_o[25]), 
	.A1(n16966));
   OAI22_X1 U2145 (.ZN(n2475), 
	.B2(n2490), 
	.B1(n2131), 
	.A2(n4951), 
	.A1(n16992));
   INV_X1 U2146 (.ZN(n4951), 
	.A(n2490));
   OAI22_X1 U2147 (.ZN(n2490), 
	.B2(n2493), 
	.B1(n2248), 
	.A2(n2492), 
	.A1(n2491));
   INV_X1 U2148 (.ZN(n2491), 
	.A(n2248));
   OAI22_X1 U2149 (.ZN(U598_Z_0), 
	.B2(n17005), 
	.B1(n2494), 
	.A2(n17001), 
	.A1(FE_PHN3553_n5647));
   OAI22_X1 U2150 (.ZN(U597_Z_0), 
	.B2(n17000), 
	.B1(n2494), 
	.A2(n16996), 
	.A1(n5646));
   OAI22_X1 U2151 (.ZN(U596_Z_0), 
	.B2(n17042), 
	.B1(n2494), 
	.A2(n17038), 
	.A1(FE_PHN3635_n5645));
   OAI22_X1 U2152 (.ZN(U595_Z_0), 
	.B2(n17037), 
	.B1(n2494), 
	.A2(n17033), 
	.A1(n5644));
   OAI22_X1 U2153 (.ZN(U594_Z_0), 
	.B2(n17031), 
	.B1(n2494), 
	.A2(n17028), 
	.A1(n4972));
   OAI22_X1 U2154 (.ZN(U593_Z_0), 
	.B2(n17027), 
	.B1(n2494), 
	.A2(n17023), 
	.A1(FE_PHN3642_n5179));
   OAI22_X1 U2155 (.ZN(U592_Z_0), 
	.B2(n17022), 
	.B1(n2494), 
	.A2(n17018), 
	.A1(FE_PHN3583_n4980));
   OAI22_X1 U2156 (.ZN(U591_Z_0), 
	.B2(n17017), 
	.B1(n2494), 
	.A2(n17013), 
	.A1(n5208));
   OAI22_X1 U2157 (.ZN(U590_Z_0), 
	.B2(n17046), 
	.B1(n2494), 
	.A2(n17043), 
	.A1(n5315));
   OAI22_X1 U2158 (.ZN(U589_Z_0), 
	.B2(n17052), 
	.B1(n2494), 
	.A2(n17048), 
	.A1(n5344));
   OAI22_X1 U2159 (.ZN(U588_Z_0), 
	.B2(n17057), 
	.B1(n2494), 
	.A2(n17053), 
	.A1(FE_PHN3559_n5373));
   OAI22_X1 U2160 (.ZN(U587_Z_0), 
	.B2(n17062), 
	.B1(n2494), 
	.A2(n17058), 
	.A1(FE_PHN3605_n5402));
   OAI22_X1 U2161 (.ZN(U586_Z_0), 
	.B2(n17067), 
	.B1(n2494), 
	.A2(n17063), 
	.A1(n5431));
   OAI22_X1 U2162 (.ZN(U585_Z_0), 
	.B2(n17071), 
	.B1(n2494), 
	.A2(n17068), 
	.A1(n5460));
   OAI22_X1 U2163 (.ZN(U584_Z_0), 
	.B2(n17077), 
	.B1(n2494), 
	.A2(n17074), 
	.A1(FE_PHN4831_n4982));
   OAI22_X1 U2164 (.ZN(U583_Z_0), 
	.B2(n17082), 
	.B1(n2494), 
	.A2(n17078), 
	.A1(n5484));
   AOI221_X1 U2166 (.ZN(n2109), 
	.C2(n17008), 
	.C1(FE_OFN537_n2496), 
	.B2(n16701), 
	.B1(n2495), 
	.A(n2497));
   INV_X1 U2167 (.ZN(n2497), 
	.A(n2498));
   AOI211_X1 U2168 (.ZN(n2498), 
	.C2(U163_Z_0), 
	.C1(n2499), 
	.B(n2500), 
	.A(n2055));
   NOR3_X1 U2169 (.ZN(n2500), 
	.A3(n16992), 
	.A2(U163_Z_0), 
	.A1(n1684));
   OAI22_X1 U2170 (.ZN(n2499), 
	.B2(n1648), 
	.B1(FE_OFN538_n2501), 
	.A2(n1684), 
	.A1(n2131));
   INV_X1 U2171 (.ZN(n1684), 
	.A(n1648));
   NAND4_X1 U2172 (.ZN(n1648), 
	.A4(n2505), 
	.A3(n2504), 
	.A2(n2503), 
	.A1(n2502));
   AOI222_X1 U2173 (.ZN(n2505), 
	.C2(vis_psp_o[22]), 
	.C1(n16967), 
	.B2(n2507), 
	.B1(n16972), 
	.A2(vis_msp_o[22]), 
	.A1(n16973));
   AOI222_X1 U2175 (.ZN(n2504), 
	.C2(vis_r11_o[24]), 
	.C1(n16986), 
	.B2(vis_r12_o[24]), 
	.B1(FE_OFN109_n16964), 
	.A2(vis_r14_o[24]), 
	.A1(n16983));
   AOI222_X1 U2178 (.ZN(n2503), 
	.C2(vis_r8_o[24]), 
	.C1(n16958), 
	.B2(vis_r10_o[24]), 
	.B1(n16961), 
	.A2(vis_r9_o[24]), 
	.A1(n16979));
   AOI22_X1 U2180 (.ZN(n2502), 
	.B2(n2515), 
	.B1(n16954), 
	.A2(n2481), 
	.A1(n16977));
   INV_X1 U2182 (.ZN(n109), 
	.A(FE_PHN752_n1337));
   OAI221_X1 U2183 (.ZN(n1337), 
	.C2(n2091), 
	.C1(n2517), 
	.B2(n2089), 
	.B1(FE_PHN685_n2516), 
	.A(n2518));
   AOI221_X1 U2184 (.ZN(n2518), 
	.C2(n2067), 
	.C1(n2023), 
	.B2(n2019), 
	.B1(n2074), 
	.A(n2076));
   INV_X1 U2185 (.ZN(n2091), 
	.A(n2069));
   INV_X1 U2186 (.ZN(n2089), 
	.A(n2072));
   OAI22_X1 U2187 (.ZN(U582_Z_0), 
	.B2(n17005), 
	.B1(n2519), 
	.A2(n17001), 
	.A1(FE_PHN2615_n5045));
   OAI22_X1 U2188 (.ZN(U581_Z_0), 
	.B2(n17000), 
	.B1(n2519), 
	.A2(n16996), 
	.A1(FE_PHN2526_n5044));
   OAI22_X1 U2189 (.ZN(U580_Z_0), 
	.B2(n17042), 
	.B1(n2519), 
	.A2(n17038), 
	.A1(FE_PHN2524_n5292));
   OAI22_X1 U2190 (.ZN(U579_Z_0), 
	.B2(n17037), 
	.B1(n2519), 
	.A2(n17033), 
	.A1(FE_PHN2580_n5271));
   OAI22_X1 U2191 (.ZN(U578_Z_0), 
	.B2(n17031), 
	.B1(FE_OFN539_n2519), 
	.A2(n17028), 
	.A1(FE_PHN2689_n5043));
   OAI22_X1 U2192 (.ZN(U577_Z_0), 
	.B2(n17027), 
	.B1(n2519), 
	.A2(n17023), 
	.A1(FE_PHN2643_n5180));
   OAI22_X1 U2193 (.ZN(U576_Z_0), 
	.B2(n17022), 
	.B1(n2519), 
	.A2(n17018), 
	.A1(FE_PHN2495_n5042));
   OAI22_X1 U2194 (.ZN(U575_Z_0), 
	.B2(n17017), 
	.B1(n2519), 
	.A2(n17013), 
	.A1(FE_PHN2536_n5209));
   OAI22_X1 U2195 (.ZN(U574_Z_0), 
	.B2(n17046), 
	.B1(n2519), 
	.A2(n17043), 
	.A1(FE_PHN2554_n5316));
   OAI22_X1 U2196 (.ZN(U573_Z_0), 
	.B2(n17052), 
	.B1(n2519), 
	.A2(n17048), 
	.A1(FE_PHN2454_n5345));
   OAI22_X1 U2197 (.ZN(U572_Z_0), 
	.B2(n17057), 
	.B1(n2519), 
	.A2(n17053), 
	.A1(FE_PHN2587_n5374));
   OAI22_X1 U2198 (.ZN(U571_Z_0), 
	.B2(n17062), 
	.B1(n2519), 
	.A2(n17058), 
	.A1(FE_PHN2582_n5403));
   OAI22_X1 U2199 (.ZN(U570_Z_0), 
	.B2(n17067), 
	.B1(FE_OFN539_n2519), 
	.A2(n17063), 
	.A1(FE_PHN2705_n5432));
   OAI22_X1 U2200 (.ZN(U569_Z_0), 
	.B2(n17071), 
	.B1(FE_OFN539_n2519), 
	.A2(n17068), 
	.A1(FE_PHN2755_n5461));
   OAI22_X1 U2201 (.ZN(U568_Z_0), 
	.B2(n17077), 
	.B1(FE_OFN539_n2519), 
	.A2(n17074), 
	.A1(FE_PHN2680_n5041));
   OAI22_X1 U2202 (.ZN(U567_Z_0), 
	.B2(n17082), 
	.B1(FE_OFN539_n2519), 
	.A2(n17078), 
	.A1(FE_PHN2723_n5485));
   OR3_X1 U2204 (.ZN(n2521), 
	.A3(n2524), 
	.A2(n2523), 
	.A1(n2522));
   NOR3_X1 U2205 (.ZN(n2524), 
	.A3(n2525), 
	.A2(n2501), 
	.A1(n2161));
   INV_X1 U2206 (.ZN(n2523), 
	.A(n2235));
   OAI221_X1 U2207 (.ZN(n2235), 
	.C2(n2127), 
	.C1(n5817), 
	.B2(n2525), 
	.B1(n2126), 
	.A(n2161));
   NAND4_X1 U2208 (.ZN(n2161), 
	.A4(n2529), 
	.A3(n2528), 
	.A2(n2527), 
	.A1(n2526));
   AOI222_X1 U2209 (.ZN(n2529), 
	.C2(vis_psp_o[4]), 
	.C1(n16967), 
	.B2(n2531), 
	.B1(n16972), 
	.A2(vis_msp_o[4]), 
	.A1(n16973));
   AOI222_X1 U2210 (.ZN(n2528), 
	.C2(vis_r11_o[6]), 
	.C1(n16985), 
	.B2(vis_r12_o[6]), 
	.B1(FE_OFN109_n16964), 
	.A2(vis_r14_o[6]), 
	.A1(n16982));
   AOI222_X1 U2211 (.ZN(n2527), 
	.C2(vis_r8_o[6]), 
	.C1(n16958), 
	.B2(vis_r10_o[6]), 
	.B1(n16961), 
	.A2(vis_r9_o[6]), 
	.A1(n16979));
   AOI22_X1 U2212 (.ZN(n2526), 
	.B2(n2539), 
	.B1(n16954), 
	.A2(n1152), 
	.A1(n16977));
   INV_X1 U2213 (.ZN(n2525), 
	.A(n5817));
   XOR2_X1 U2214 (.Z(n5817), 
	.B(n2540), 
	.A(n16990));
   AOI221_X1 U2215 (.ZN(n2540), 
	.C2(n2250), 
	.C1(n16988), 
	.B2(FE_OFN15_n16671), 
	.B1(n2541), 
	.A(n2542));
   OAI22_X1 U2216 (.ZN(n2542), 
	.B2(n2201), 
	.B1(n5257), 
	.A2(n2543), 
	.A1(n5244));
   INV_X1 U2217 (.ZN(n2541), 
	.A(n2200));
   AOI21_X1 U2218 (.ZN(n2522), 
	.B2(n16782), 
	.B1(n2124), 
	.A(n2544));
   INV_X1 U2220 (.ZN(n2520), 
	.A(n148));
   AOI221_X1 U2221 (.ZN(n148), 
	.C2(n2546), 
	.C1(n2008), 
	.B2(n2545), 
	.B1(n2004), 
	.A(n2547));
   INV_X1 U2222 (.ZN(n2547), 
	.A(n2548));
   AOI221_X1 U2223 (.ZN(n2548), 
	.C2(n2011), 
	.C1(n2094), 
	.B2(n2002), 
	.B1(n2093), 
	.A(n2012));
   OAI22_X1 U2224 (.ZN(U566_Z_0), 
	.B2(n17005), 
	.B1(n2549), 
	.A2(n17001), 
	.A1(n5095));
   OAI22_X1 U2225 (.ZN(U565_Z_0), 
	.B2(n17000), 
	.B1(n2549), 
	.A2(n16996), 
	.A1(FE_PHN3601_n5094));
   OAI22_X1 U2226 (.ZN(U564_Z_0), 
	.B2(n17042), 
	.B1(n2549), 
	.A2(n17038), 
	.A1(FE_PHN3586_n5293));
   OAI22_X1 U2227 (.ZN(U563_Z_0), 
	.B2(n17037), 
	.B1(n2549), 
	.A2(n17033), 
	.A1(n5272));
   OAI22_X1 U2228 (.ZN(U562_Z_0), 
	.B2(n17031), 
	.B1(n2549), 
	.A2(n17028), 
	.A1(FE_PHN2664_n5093));
   OAI22_X1 U2229 (.ZN(U561_Z_0), 
	.B2(n17027), 
	.B1(n2549), 
	.A2(n17023), 
	.A1(FE_PHN2719_n5181));
   OAI22_X1 U2230 (.ZN(U560_Z_0), 
	.B2(n17022), 
	.B1(n2549), 
	.A2(n17018), 
	.A1(FE_PHN2473_n5092));
   OAI22_X1 U2231 (.ZN(U559_Z_0), 
	.B2(n17017), 
	.B1(n2549), 
	.A2(n17013), 
	.A1(FE_PHN2441_n5210));
   OAI22_X1 U2232 (.ZN(U558_Z_0), 
	.B2(n17046), 
	.B1(n2549), 
	.A2(n17043), 
	.A1(FE_PHN2545_n5317));
   OAI22_X1 U2233 (.ZN(U557_Z_0), 
	.B2(n17052), 
	.B1(n2549), 
	.A2(n17048), 
	.A1(n5346));
   OAI22_X1 U2234 (.ZN(U556_Z_0), 
	.B2(n17057), 
	.B1(n2549), 
	.A2(n17053), 
	.A1(FE_PHN3564_n5375));
   OAI22_X1 U2235 (.ZN(U555_Z_0), 
	.B2(n17062), 
	.B1(n2549), 
	.A2(n17058), 
	.A1(FE_PHN3565_n5404));
   OAI22_X1 U2236 (.ZN(U554_Z_0), 
	.B2(n17067), 
	.B1(n2549), 
	.A2(n17063), 
	.A1(FE_PHN2721_n5433));
   OAI22_X1 U2237 (.ZN(U553_Z_0), 
	.B2(n17071), 
	.B1(n2549), 
	.A2(n17068), 
	.A1(FE_PHN2699_n5462));
   OAI22_X1 U2238 (.ZN(U552_Z_0), 
	.B2(n17077), 
	.B1(n2549), 
	.A2(n17074), 
	.A1(FE_PHN2673_n5091));
   OAI22_X1 U2239 (.ZN(U551_Z_0), 
	.B2(n17082), 
	.B1(n2549), 
	.A2(n17078), 
	.A1(FE_PHN2744_n5486));
   OAI221_X1 U2241 (.ZN(n2281), 
	.C2(n1634), 
	.C1(n16994), 
	.B2(n5802), 
	.B1(n2550), 
	.A(n2551));
   NAND3_X1 U2242 (.ZN(n2551), 
	.A3(n5802), 
	.A2(n1634), 
	.A1(n2131));
   XOR2_X1 U2243 (.Z(n5802), 
	.B(n16991), 
	.A(n2552));
   OAI221_X1 U2244 (.ZN(n2552), 
	.C2(n2554), 
	.C1(n5100), 
	.B2(n2201), 
	.B1(n5256), 
	.A(n2555));
   AOI22_X1 U2245 (.ZN(n2555), 
	.B2(n781), 
	.B1(n2198), 
	.A2(n2556), 
	.A1(n16988));
   NOR2_X1 U2246 (.ZN(n2550), 
	.A2(n16992), 
	.A1(n1673));
   INV_X1 U2247 (.ZN(n1673), 
	.A(n1634));
   NAND4_X1 U2248 (.ZN(n1634), 
	.A4(n2560), 
	.A3(n2559), 
	.A2(n2558), 
	.A1(n2557));
   AOI222_X1 U2249 (.ZN(n2560), 
	.C2(vis_psp_o[3]), 
	.C1(n16967), 
	.B2(n2562), 
	.B1(n16971), 
	.A2(vis_msp_o[3]), 
	.A1(n16973));
   AOI222_X1 U2250 (.ZN(n2559), 
	.C2(vis_r11_o[5]), 
	.C1(n16986), 
	.B2(vis_r12_o[5]), 
	.B1(FE_OFN109_n16964), 
	.A2(vis_r14_o[5]), 
	.A1(n16982));
   AOI222_X1 U2251 (.ZN(n2558), 
	.C2(vis_r8_o[5]), 
	.C1(n16958), 
	.B2(vis_r10_o[5]), 
	.B1(n16962), 
	.A2(vis_r9_o[5]), 
	.A1(n16979));
   AOI22_X1 U2252 (.ZN(n2557), 
	.B2(n2570), 
	.B1(n16954), 
	.A2(n2539), 
	.A1(n16977));
   NAND2_X1 U2253 (.ZN(n2263), 
	.A2(FE_OFN2_n2015), 
	.A1(n16731));
   AOI221_X1 U2254 (.ZN(n2107), 
	.C2(n17008), 
	.C1(n2556), 
	.B2(n2227), 
	.B1(vis_ipsr_o[5]), 
	.A(n2055));
   AOI221_X1 U2255 (.ZN(n152), 
	.C2(n2004), 
	.C1(FE_PHN748_n2415), 
	.B2(n2011), 
	.B1(n2410), 
	.A(n2571));
   INV_X1 U2256 (.ZN(n2571), 
	.A(n2572));
   AOI221_X1 U2257 (.ZN(n2572), 
	.C2(n2002), 
	.C1(n2411), 
	.B2(n2414), 
	.B1(n2008), 
	.A(n2012));
   OAI22_X1 U2258 (.ZN(U550_Z_0), 
	.B2(n17005), 
	.B1(n2573), 
	.A2(n17001), 
	.A1(FE_PHN2578_n5125));
   OAI22_X1 U2259 (.ZN(U549_Z_0), 
	.B2(n17000), 
	.B1(n2573), 
	.A2(n16996), 
	.A1(FE_PHN2509_n5124));
   OAI22_X1 U2260 (.ZN(U548_Z_0), 
	.B2(n17042), 
	.B1(n2573), 
	.A2(n17038), 
	.A1(FE_PHN2490_n5294));
   OAI22_X1 U2261 (.ZN(U547_Z_0), 
	.B2(n17037), 
	.B1(n2573), 
	.A2(n17033), 
	.A1(FE_PHN2619_n5273));
   OAI22_X1 U2262 (.ZN(U546_Z_0), 
	.B2(n17031), 
	.B1(n2573), 
	.A2(n17028), 
	.A1(FE_PHN2679_n5123));
   OAI22_X1 U2263 (.ZN(U545_Z_0), 
	.B2(n17027), 
	.B1(n2573), 
	.A2(n17023), 
	.A1(FE_PHN2649_n5182));
   OAI22_X1 U2264 (.ZN(U544_Z_0), 
	.B2(n17022), 
	.B1(n2573), 
	.A2(n17018), 
	.A1(FE_PHN2472_n5122));
   OAI22_X1 U2265 (.ZN(U543_Z_0), 
	.B2(n17017), 
	.B1(n2573), 
	.A2(n17013), 
	.A1(FE_PHN2537_n5211));
   OAI22_X1 U2266 (.ZN(U542_Z_0), 
	.B2(n17046), 
	.B1(n2573), 
	.A2(n17043), 
	.A1(FE_PHN2464_n5318));
   OAI22_X1 U2267 (.ZN(U541_Z_0), 
	.B2(n17052), 
	.B1(n2573), 
	.A2(n17048), 
	.A1(FE_PHN2539_n5347));
   OAI22_X1 U2268 (.ZN(U540_Z_0), 
	.B2(n17057), 
	.B1(n2573), 
	.A2(n17053), 
	.A1(FE_PHN2532_n5376));
   OAI22_X1 U2269 (.ZN(U539_Z_0), 
	.B2(n17062), 
	.B1(n2573), 
	.A2(n17058), 
	.A1(FE_PHN2573_n5405));
   OAI22_X1 U2270 (.ZN(U538_Z_0), 
	.B2(n17067), 
	.B1(n2573), 
	.A2(n17063), 
	.A1(FE_PHN2669_n5434));
   OAI22_X1 U2271 (.ZN(U537_Z_0), 
	.B2(n17071), 
	.B1(n2573), 
	.A2(n17068), 
	.A1(FE_PHN2729_n5463));
   OAI22_X1 U2272 (.ZN(U536_Z_0), 
	.B2(n17077), 
	.B1(n2573), 
	.A2(n17074), 
	.A1(FE_PHN2742_n5121));
   OAI22_X1 U2273 (.ZN(U535_Z_0), 
	.B2(n17082), 
	.B1(n2573), 
	.A2(n17078), 
	.A1(FE_PHN2782_n5487));
   OAI221_X1 U2275 (.ZN(n2283), 
	.C2(n1636), 
	.C1(n16994), 
	.B2(n5801), 
	.B1(n2574), 
	.A(n2575));
   NAND3_X1 U2276 (.ZN(n2575), 
	.A3(n5801), 
	.A2(n1636), 
	.A1(n2131));
   XOR2_X1 U2277 (.Z(n5801), 
	.B(n2576), 
	.A(n16990));
   AOI221_X1 U2278 (.ZN(n2576), 
	.C2(n2578), 
	.C1(n16988), 
	.B2(n2577), 
	.B1(n16656), 
	.A(n2579));
   OAI22_X1 U2279 (.ZN(n2579), 
	.B2(n2201), 
	.B1(n16810), 
	.A2(n2543), 
	.A1(n16794));
   NOR2_X1 U2280 (.ZN(n2574), 
	.A2(n16992), 
	.A1(n1674));
   INV_X1 U2281 (.ZN(n1674), 
	.A(n1636));
   NAND4_X1 U2282 (.ZN(n1636), 
	.A4(n2583), 
	.A3(n2582), 
	.A2(n2581), 
	.A1(n2580));
   AOI222_X1 U2283 (.ZN(n2583), 
	.C2(vis_psp_o[2]), 
	.C1(n16967), 
	.B2(n2585), 
	.B1(n16971), 
	.A2(vis_msp_o[2]), 
	.A1(n16973));
   AOI222_X1 U2284 (.ZN(n2582), 
	.C2(vis_r11_o[4]), 
	.C1(n16986), 
	.B2(vis_r12_o[4]), 
	.B1(n16965), 
	.A2(vis_r14_o[4]), 
	.A1(n16982));
   AOI222_X1 U2285 (.ZN(n2581), 
	.C2(vis_r8_o[4]), 
	.C1(n16959), 
	.B2(vis_r10_o[4]), 
	.B1(n16962), 
	.A2(vis_r9_o[4]), 
	.A1(n16979));
   AOI22_X1 U2286 (.ZN(n2580), 
	.B2(n2593), 
	.B1(n16954), 
	.A2(n2570), 
	.A1(n16977));
   NAND2_X1 U2287 (.ZN(n2262), 
	.A2(FE_OFN2_n2015), 
	.A1(n16730));
   AOI221_X1 U2288 (.ZN(n2112), 
	.C2(n17008), 
	.C1(n2578), 
	.B2(n2227), 
	.B1(vis_ipsr_o[4]), 
	.A(n2055));
   AOI221_X1 U2289 (.ZN(n160), 
	.C2(n2004), 
	.C1(n2068), 
	.B2(n2011), 
	.B1(n2066), 
	.A(n2594));
   INV_X1 U2290 (.ZN(n2594), 
	.A(n2595));
   AOI221_X1 U2291 (.ZN(n2595), 
	.C2(n2075), 
	.C1(n2002), 
	.B2(n2073), 
	.B1(n2008), 
	.A(n2012));
   INV_X1 U2292 (.ZN(n2073), 
	.A(n2596));
   OAI22_X1 U2293 (.ZN(U534_Z_0), 
	.B2(n17005), 
	.B1(n2597), 
	.A2(n17001), 
	.A1(FE_PHN3581_n5032));
   OAI22_X1 U2294 (.ZN(U533_Z_0), 
	.B2(n17000), 
	.B1(n2597), 
	.A2(n16996), 
	.A1(FE_PHN3566_n5031));
   OAI22_X1 U2295 (.ZN(U532_Z_0), 
	.B2(n17042), 
	.B1(n2597), 
	.A2(n17038), 
	.A1(FE_PHN3577_n5295));
   OAI22_X1 U2296 (.ZN(U531_Z_0), 
	.B2(n17037), 
	.B1(n2597), 
	.A2(n17033), 
	.A1(FE_PHN3557_n5274));
   OAI22_X1 U2297 (.ZN(U530_Z_0), 
	.B2(n17031), 
	.B1(n2597), 
	.A2(n17028), 
	.A1(FE_PHN2685_n5030));
   OAI22_X1 U2298 (.ZN(U529_Z_0), 
	.B2(n17027), 
	.B1(n2597), 
	.A2(n17023), 
	.A1(FE_PHN2667_n5183));
   OAI22_X1 U2299 (.ZN(U528_Z_0), 
	.B2(n17022), 
	.B1(n2597), 
	.A2(n17018), 
	.A1(n5029));
   OAI22_X1 U2300 (.ZN(U527_Z_0), 
	.B2(n17017), 
	.B1(n2597), 
	.A2(n17013), 
	.A1(FE_PHN2520_n5212));
   OAI22_X1 U2301 (.ZN(U526_Z_0), 
	.B2(n17046), 
	.B1(n2597), 
	.A2(n17043), 
	.A1(FE_PHN2564_n5319));
   OAI22_X1 U2302 (.ZN(U525_Z_0), 
	.B2(n17052), 
	.B1(n2597), 
	.A2(n17048), 
	.A1(FE_PHN2628_n5348));
   OAI22_X1 U2303 (.ZN(U524_Z_0), 
	.B2(n17057), 
	.B1(n2597), 
	.A2(n17053), 
	.A1(FE_PHN3599_n5377));
   OAI22_X1 U2304 (.ZN(U523_Z_0), 
	.B2(n17062), 
	.B1(n2597), 
	.A2(n17058), 
	.A1(FE_PHN3578_n5406));
   OAI22_X1 U2305 (.ZN(U522_Z_0), 
	.B2(n17067), 
	.B1(n2597), 
	.A2(n17063), 
	.A1(FE_PHN2659_n5435));
   OAI22_X1 U2306 (.ZN(U521_Z_0), 
	.B2(n17071), 
	.B1(n2597), 
	.A2(n17068), 
	.A1(FE_PHN2734_n5464));
   OAI22_X1 U2307 (.ZN(U520_Z_0), 
	.B2(n17077), 
	.B1(n2597), 
	.A2(n17074), 
	.A1(FE_PHN2634_n5028));
   OAI22_X1 U2308 (.ZN(U519_Z_0), 
	.B2(n17082), 
	.B1(n2597), 
	.A2(n17078), 
	.A1(n5488));
   AOI222_X1 U2310 (.ZN(n2598), 
	.C2(n2055), 
	.C1(n2032), 
	.B2(FE_OFN2_n2015), 
	.B1(n16682), 
	.A2(n2257), 
	.A1(n17008));
   INV_X1 U2311 (.ZN(n2032), 
	.A(n2599));
   INV_X1 U2312 (.ZN(n2111), 
	.A(n2600));
   OAI221_X1 U2313 (.ZN(n2600), 
	.C2(n2164), 
	.C1(n170), 
	.B2(n2602), 
	.B1(n2601), 
	.A(n2603));
   NAND3_X1 U2314 (.ZN(n2603), 
	.A3(n2602), 
	.A2(n2127), 
	.A1(n2604));
   INV_X1 U2315 (.ZN(n2164), 
	.A(n2227));
   INV_X1 U2316 (.ZN(n2602), 
	.A(add_2082_B_4_));
   XOR2_X1 U2317 (.Z(add_2082_B_4_), 
	.B(n16991), 
	.A(n2605));
   OAI221_X1 U2318 (.ZN(n2605), 
	.C2(n2554), 
	.C1(n5027), 
	.B2(n2201), 
	.B1(n5100), 
	.A(n2606));
   AOI22_X1 U2319 (.ZN(n2606), 
	.B2(n454), 
	.B1(n2198), 
	.A2(n2257), 
	.A1(n16989));
   AOI22_X1 U2320 (.ZN(n2601), 
	.B2(n2126), 
	.B1(n2604), 
	.A2(n16994), 
	.A1(n1638));
   INV_X4 U2321 (.ZN(n1638), 
	.A(n2604));
   NAND4_X2 U2322 (.ZN(n2604), 
	.A4(n2610), 
	.A3(n2609), 
	.A2(n2608), 
	.A1(n2607));
   AOI222_X1 U2323 (.ZN(n2610), 
	.C2(vis_psp_o[1]), 
	.C1(n16968), 
	.B2(n2612), 
	.B1(n16971), 
	.A2(vis_msp_o[1]), 
	.A1(n16973));
   AOI222_X1 U2324 (.ZN(n2609), 
	.C2(vis_r11_o[3]), 
	.C1(n16986), 
	.B2(vis_r12_o[3]), 
	.B1(n16965), 
	.A2(vis_r14_o[3]), 
	.A1(n16982));
   AOI222_X1 U2325 (.ZN(n2608), 
	.C2(vis_r8_o[3]), 
	.C1(n16959), 
	.B2(vis_r10_o[3]), 
	.B1(n16962), 
	.A2(vis_r9_o[3]), 
	.A1(n16979));
   AOI22_X1 U2326 (.ZN(n2607), 
	.B2(n2620), 
	.B1(n16955), 
	.A2(n2593), 
	.A1(n16977));
   AOI221_X1 U2327 (.ZN(n166), 
	.C2(n2004), 
	.C1(n2422), 
	.B2(n2002), 
	.B1(FE_PHN728_n2421), 
	.A(n2621));
   INV_X1 U2328 (.ZN(n2621), 
	.A(n2622));
   AOI221_X1 U2329 (.ZN(n2622), 
	.C2(n2011), 
	.C1(FE_PHN859_n2624), 
	.B2(n2008), 
	.B1(n2623), 
	.A(FE_OFN509_n2012));
   OAI22_X1 U2330 (.ZN(U518_Z_0), 
	.B2(n1811), 
	.B1(n683), 
	.A2(n980), 
	.A1(n5102));
   OAI222_X1 U2334 (.ZN(n2627), 
	.C2(n782), 
	.C1(FE_OFN81_n16856), 
	.B2(n1027), 
	.B1(n16837), 
	.A2(n2628), 
	.A1(n16957));
   OAI221_X1 U2335 (.ZN(n2626), 
	.C2(n1857), 
	.C1(n16826), 
	.B2(n16828), 
	.B1(n2629), 
	.A(n2630));
   NAND3_X1 U2336 (.ZN(n2630), 
	.A3(n2631), 
	.A2(n16851), 
	.A1(FE_OFN75_n16806));
   AOI21_X1 U2337 (.ZN(n2629), 
	.B2(n565), 
	.B1(n1564), 
	.A(n1606));
   NAND3_X2 U2338 (.ZN(n2232), 
	.A3(n2634), 
	.A2(n2633), 
	.A1(n2632));
   AOI221_X2 U2339 (.ZN(n2634), 
	.C2(n2188), 
	.C1(n16956), 
	.B2(n2635), 
	.B1(n16976), 
	.A(n2636));
   OAI22_X1 U2340 (.ZN(n2636), 
	.B2(n2190), 
	.B1(n5395), 
	.A2(n2637), 
	.A1(n5366));
   AOI222_X1 U2342 (.ZN(n2633), 
	.C2(vis_r12_o[1]), 
	.C1(n16964), 
	.B2(n2639), 
	.B1(n16971), 
	.A2(vis_r11_o[1]), 
	.A1(n16985));
   AOI22_X1 U2343 (.ZN(n2632), 
	.B2(vis_r10_o[1]), 
	.B1(n16963), 
	.A2(vis_r14_o[1]), 
	.A1(n16984));
   AOI222_X1 U2348 (.ZN(n2645), 
	.C2(n16828), 
	.C1(n2646), 
	.B2(n16954), 
	.B1(n2628), 
	.A2(n16836), 
	.A1(n1806));
   INV_X1 U2349 (.ZN(n1806), 
	.A(n919));
   NAND4_X1 U2350 (.ZN(n2643), 
	.A4(n2647), 
	.A3(n673), 
	.A2(FE_OFN72_n16867), 
	.A1(n1103));
   AOI21_X1 U2351 (.ZN(n2647), 
	.B2(n502), 
	.B1(n1561), 
	.A(n611));
   INV_X1 U2352 (.ZN(n502), 
	.A(n1218));
   XOR2_X1 U2353 (.Z(n2625), 
	.B(n1106), 
	.A(n4973));
   OAI21_X1 U2354 (.ZN(n1106), 
	.B2(n187), 
	.B1(n1007), 
	.A(n1008));
   AOI21_X1 U2356 (.ZN(n187), 
	.B2(n1563), 
	.B1(n16845), 
	.A(n943));
   INV_X1 U2357 (.ZN(n943), 
	.A(n1217));
   NAND2_X1 U2358 (.ZN(n1217), 
	.A2(n16728), 
	.A1(n483));
   INV_X1 U2359 (.ZN(n1563), 
	.A(n846));
   NAND2_X1 U2360 (.ZN(n846), 
	.A2(FE_OFN85_n16839), 
	.A1(n16868));
   AND3_X1 U2361 (.ZN(n1007), 
	.A3(n2650), 
	.A2(n2649), 
	.A1(n2648));
   NOR4_X1 U2362 (.ZN(n2650), 
	.A4(n2654), 
	.A3(n2653), 
	.A2(n2652), 
	.A1(n2651));
   NOR4_X1 U2363 (.ZN(n2654), 
	.A4(n604), 
	.A3(n1519), 
	.A2(n16820), 
	.A1(n16836));
   NOR4_X1 U2364 (.ZN(n2653), 
	.A4(n498), 
	.A3(FE_OFN98_n1104), 
	.A2(n16859), 
	.A1(FE_OFN100_n1086));
   NAND2_X1 U2365 (.ZN(n498), 
	.A2(n16821), 
	.A1(FE_OFN79_n16834));
   INV_X1 U2366 (.ZN(n2652), 
	.A(n2655));
   OAI211_X1 U2367 (.ZN(n2655), 
	.C2(n542), 
	.C1(n998), 
	.B(FE_OFN104_n715), 
	.A(n566));
   OAI33_X1 U2368 (.ZN(n2651), 
	.B3(FE_OFN17_n16805), 
	.B2(n16833), 
	.B1(n648), 
	.A3(n917), 
	.A2(n1218), 
	.A1(n532));
   AOI22_X1 U2369 (.ZN(n2649), 
	.B2(n2657), 
	.B1(n757), 
	.A2(n596), 
	.A1(n2656));
   NAND4_X1 U2370 (.ZN(n2657), 
	.A4(n1579), 
	.A3(n1856), 
	.A2(n918), 
	.A1(FE_OFN70_n16867));
   NAND2_X1 U2371 (.ZN(n2656), 
	.A2(n2659), 
	.A1(n2658));
   NAND3_X1 U2372 (.ZN(n2659), 
	.A3(n1095), 
	.A2(n1574), 
	.A1(n991));
   AOI22_X1 U2373 (.ZN(n2648), 
	.B2(n2662), 
	.B1(n2661), 
	.A2(n16826), 
	.A1(n2660));
   NAND4_X1 U2374 (.ZN(n2660), 
	.A4(n2664), 
	.A3(n2663), 
	.A2(n694), 
	.A1(n1857));
   AOI221_X1 U2375 (.ZN(n2664), 
	.C2(n16808), 
	.C1(n527), 
	.B2(n16728), 
	.B1(n897), 
	.A(n2665));
   OAI22_X1 U2376 (.ZN(n2665), 
	.B2(n616), 
	.B1(n556), 
	.A2(n745), 
	.A1(n605));
   AOI21_X1 U2377 (.ZN(n2663), 
	.B2(n596), 
	.B1(n2666), 
	.A(n2667));
   NOR3_X1 U2378 (.ZN(n2667), 
	.A3(FE_OFN107_n585), 
	.A2(n16845), 
	.A1(n16808));
   OAI21_X1 U2380 (.ZN(n2666), 
	.B2(n16828), 
	.B1(n2668), 
	.A(n2669));
   NAND3_X1 U2381 (.ZN(n2669), 
	.A3(n16804), 
	.A2(n1574), 
	.A1(n592));
   AOI222_X1 U2382 (.ZN(n2668), 
	.C2(n1468), 
	.C1(n2672), 
	.B2(n466), 
	.B1(n2671), 
	.A2(n2670), 
	.A1(n592));
   NOR2_X1 U2383 (.ZN(n2671), 
	.A2(n1469), 
	.A1(FE_OFN631_n16851));
   INV_X1 U2384 (.ZN(n2670), 
	.A(n2673));
   NOR4_X1 U2387 (.ZN(n2677), 
	.A4(n2681), 
	.A3(n2680), 
	.A2(n2679), 
	.A1(n2678));
   NOR4_X1 U2388 (.ZN(n2681), 
	.A4(n762), 
	.A3(n917), 
	.A2(FE_OFN100_n1086), 
	.A1(n16694));
   INV_X1 U2389 (.ZN(n2680), 
	.A(n1177));
   AND3_X1 U2390 (.ZN(n2679), 
	.A3(n809), 
	.A2(n1094), 
	.A1(n1561));
   NOR2_X1 U2391 (.ZN(n1561), 
	.A2(n16851), 
	.A1(n16826));
   OAI33_X1 U2392 (.ZN(n2678), 
	.B3(n16808), 
	.B2(n16859), 
	.B1(n524), 
	.A3(n616), 
	.A2(n16836), 
	.A1(n713));
   AOI21_X1 U2393 (.ZN(n2676), 
	.B2(n16864), 
	.B1(n2682), 
	.A(n2683));
   OAI33_X1 U2394 (.ZN(n2683), 
	.B3(FE_OFN627_n16828), 
	.B2(n16845), 
	.B1(FE_OFN465_n945), 
	.A3(FE_OFN103_n715), 
	.A2(n16821), 
	.A1(n696));
   OAI211_X1 U2395 (.ZN(n2682), 
	.C2(n1857), 
	.C1(n16824), 
	.B(n1279), 
	.A(n2684));
   NAND3_X1 U2396 (.ZN(n1279), 
	.A3(n5165), 
	.A2(n16824), 
	.A1(n809));
   INV_X1 U2397 (.ZN(n2684), 
	.A(n609));
   NAND2_X1 U2398 (.ZN(n1857), 
	.A2(n1574), 
	.A1(n563));
   NAND2_X1 U2399 (.ZN(n2675), 
	.A2(FE_OFN469_n1034), 
	.A1(n660));
   INV_X1 U2400 (.ZN(n980), 
	.A(n1811));
   NAND2_X1 U2401 (.ZN(n1811), 
	.A2(hprot_o[0]), 
	.A1(n17124));
   NOR4_X1 U2403 (.ZN(n2686), 
	.A4(n2688), 
	.A3(n615), 
	.A2(n1272), 
	.A1(n2687));
   INV_X1 U2404 (.ZN(n2688), 
	.A(n1025));
   NAND3_X1 U2405 (.ZN(n1025), 
	.A3(n660), 
	.A2(n16824), 
	.A1(n827));
   NOR2_X1 U2406 (.ZN(n660), 
	.A2(FE_OFN634_n16871), 
	.A1(n558));
   INV_X1 U2407 (.ZN(n615), 
	.A(n646));
   NAND2_X1 U2408 (.ZN(n646), 
	.A2(n590), 
	.A1(n798));
   NOR3_X1 U2409 (.ZN(n1272), 
	.A3(n808), 
	.A2(n745), 
	.A1(FE_OFN422_n641));
   OAI33_X1 U2410 (.ZN(n2687), 
	.B3(n640), 
	.B2(n16859), 
	.B1(n2689), 
	.A3(n16826), 
	.A2(n16833), 
	.A1(n650));
   AOI222_X1 U2411 (.ZN(n2685), 
	.C2(n991), 
	.C1(n609), 
	.B2(n506), 
	.B1(n2690), 
	.A2(FE_OFN82_n16856), 
	.A1(n1037));
   NOR2_X1 U2412 (.ZN(n609), 
	.A2(n558), 
	.A1(n1307));
   NOR2_X1 U2413 (.ZN(n2690), 
	.A2(n808), 
	.A1(n16848));
   NOR3_X1 U2415 (.ZN(n1037), 
	.A3(n699), 
	.A2(n1467), 
	.A1(n16821));
   INV_X1 U2416 (.ZN(n2674), 
	.A(n2691));
   OAI211_X1 U2417 (.ZN(n2691), 
	.C2(n499), 
	.C1(n16833), 
	.B(n1476), 
	.A(n1024));
   AND2_X1 U2418 (.ZN(n1476), 
	.A2(n1957), 
	.A1(n2692));
   OAI21_X1 U2419 (.ZN(n2692), 
	.B2(n1306), 
	.B1(n506), 
	.A(n526));
   NOR2_X1 U2420 (.ZN(n1306), 
	.A2(n696), 
	.A1(n610));
   NAND2_X1 U2421 (.ZN(n1024), 
	.A2(n590), 
	.A1(n695));
   INV_X1 U2422 (.ZN(n590), 
	.A(n650));
   NOR2_X1 U2423 (.ZN(n695), 
	.A2(FE_OFN82_n16856), 
	.A1(n16859));
   INV_X1 U2424 (.ZN(n1876), 
	.A(n2693));
   OAI33_X1 U2425 (.ZN(n2693), 
	.B3(FE_OFN103_n715), 
	.B2(n16833), 
	.B1(n558), 
	.A3(n1882), 
	.A2(n16826), 
	.A1(n1517));
   NAND2_X1 U2426 (.ZN(n558), 
	.A2(n592), 
	.A1(n16680));
   OAI22_X1 U2427 (.ZN(U517_Z_0), 
	.B2(n17005), 
	.B1(n2694), 
	.A2(n17001), 
	.A1(FE_PHN2496_n5052));
   OAI22_X1 U2428 (.ZN(U516_Z_0), 
	.B2(n17000), 
	.B1(n2694), 
	.A2(n16996), 
	.A1(FE_PHN2690_n5051));
   OAI22_X1 U2429 (.ZN(U515_Z_0), 
	.B2(n17042), 
	.B1(n2694), 
	.A2(n17038), 
	.A1(FE_PHN2758_n5296));
   OAI22_X1 U2430 (.ZN(U514_Z_0), 
	.B2(n17037), 
	.B1(n2694), 
	.A2(n17033), 
	.A1(FE_PHN2447_n5275));
   OAI22_X1 U2431 (.ZN(U513_Z_0), 
	.B2(n17031), 
	.B1(n2694), 
	.A2(n17028), 
	.A1(n5050));
   OAI22_X1 U2432 (.ZN(U512_Z_0), 
	.B2(n17027), 
	.B1(n2694), 
	.A2(n17023), 
	.A1(FE_PHN2697_n5184));
   OAI22_X1 U2433 (.ZN(U511_Z_0), 
	.B2(n17022), 
	.B1(n2694), 
	.A2(n17018), 
	.A1(FE_PHN2586_n5049));
   OAI22_X1 U2434 (.ZN(U510_Z_0), 
	.B2(n17017), 
	.B1(n2694), 
	.A2(n17013), 
	.A1(FE_PHN2548_n5213));
   OAI22_X1 U2435 (.ZN(U509_Z_0), 
	.B2(n17046), 
	.B1(n2694), 
	.A2(n17043), 
	.A1(n5320));
   OAI22_X1 U2436 (.ZN(U508_Z_0), 
	.B2(n17052), 
	.B1(n2694), 
	.A2(FE_OFN656_n17048), 
	.A1(FE_PHN2533_n5349));
   OAI22_X1 U2437 (.ZN(U507_Z_0), 
	.B2(n17057), 
	.B1(n2694), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2522_n5378));
   OAI22_X1 U2438 (.ZN(U506_Z_0), 
	.B2(n17062), 
	.B1(n2694), 
	.A2(n17058), 
	.A1(n5407));
   OAI22_X1 U2439 (.ZN(U505_Z_0), 
	.B2(n17067), 
	.B1(n2694), 
	.A2(n17063), 
	.A1(FE_PHN2611_n5436));
   OAI22_X1 U2440 (.ZN(U504_Z_0), 
	.B2(n17071), 
	.B1(n2694), 
	.A2(n17068), 
	.A1(n5465));
   OAI22_X1 U2441 (.ZN(U503_Z_0), 
	.B2(FE_OFN666_n17077), 
	.B1(n2694), 
	.A2(n17074), 
	.A1(n5048));
   OAI22_X1 U2442 (.ZN(U502_Z_0), 
	.B2(n17082), 
	.B1(n2694), 
	.A2(n17078), 
	.A1(FE_PHN2494_n5489));
   AOI221_X1 U2444 (.ZN(n2697), 
	.C2(FE_OFN208_n2015), 
	.C1(n16702), 
	.B2(n2251), 
	.B1(n17008), 
	.A(n2698));
   INV_X1 U2445 (.ZN(n2698), 
	.A(n2282));
   OAI221_X1 U2446 (.ZN(n2282), 
	.C2(n2127), 
	.C1(n5816), 
	.B2(n2699), 
	.B1(n2126), 
	.A(n1650));
   INV_X1 U2447 (.ZN(n2699), 
	.A(n5816));
   NAND3_X1 U2448 (.ZN(n2695), 
	.A3(n1686), 
	.A2(n16994), 
	.A1(n5816));
   INV_X1 U2449 (.ZN(n1686), 
	.A(n1650));
   NAND4_X1 U2450 (.ZN(n1650), 
	.A4(n2703), 
	.A3(n2702), 
	.A2(n2701), 
	.A1(n2700));
   AOI222_X1 U2451 (.ZN(n2703), 
	.C2(vis_psp_o[20]), 
	.C1(n16968), 
	.B2(n2705), 
	.B1(n16971), 
	.A2(vis_msp_o[20]), 
	.A1(n16973));
   AOI222_X1 U2453 (.ZN(n2702), 
	.C2(vis_r11_o[22]), 
	.C1(n16986), 
	.B2(vis_r12_o[22]), 
	.B1(n16965), 
	.A2(vis_r14_o[22]), 
	.A1(n16982));
   AOI222_X1 U2456 (.ZN(n2701), 
	.C2(vis_r8_o[22]), 
	.C1(n16959), 
	.B2(vis_r10_o[22]), 
	.B1(n16962), 
	.A2(vis_r9_o[22]), 
	.A1(n16980));
   AOI22_X1 U2458 (.ZN(n2700), 
	.B2(n2714), 
	.B1(n16955), 
	.A2(n2713), 
	.A1(n16977));
   XOR2_X1 U2459 (.Z(n5816), 
	.B(n2715), 
	.A(n16990));
   AOI221_X1 U2460 (.ZN(n2715), 
	.C2(n2251), 
	.C1(n16988), 
	.B2(n16813), 
	.B1(n2716), 
	.A(n2717));
   NAND2_X1 U2461 (.ZN(n2717), 
	.A2(n2719), 
	.A1(n2718));
   NAND3_X1 U2462 (.ZN(n2718), 
	.A3(n16812), 
	.A2(n2198), 
	.A1(n5254));
   AOI221_X1 U2463 (.ZN(n61), 
	.C2(n2093), 
	.C1(n2721), 
	.B2(n2094), 
	.B1(n2720), 
	.A(n2722));
   OAI22_X1 U2464 (.ZN(n2722), 
	.B2(n2724), 
	.B1(n2088), 
	.A2(n2090), 
	.A1(n2723));
   OAI22_X1 U2465 (.ZN(U501_Z_0), 
	.B2(n17005), 
	.B1(n2725), 
	.A2(n17001), 
	.A1(FE_PHN2608_n5624));
   OAI22_X1 U2466 (.ZN(U500_Z_0), 
	.B2(n17000), 
	.B1(n2725), 
	.A2(n16996), 
	.A1(n5623));
   OAI22_X1 U2467 (.ZN(U499_Z_0), 
	.B2(n17042), 
	.B1(n2725), 
	.A2(n17038), 
	.A1(FE_PHN2783_n5622));
   OAI22_X1 U2468 (.ZN(U498_Z_0), 
	.B2(n17037), 
	.B1(n2725), 
	.A2(FE_OFN652_n17033), 
	.A1(FE_PHN2544_n5621));
   OAI22_X1 U2469 (.ZN(U497_Z_0), 
	.B2(n17031), 
	.B1(n2725), 
	.A2(n17028), 
	.A1(n5117));
   OAI22_X1 U2470 (.ZN(U496_Z_0), 
	.B2(n17027), 
	.B1(n2725), 
	.A2(n17023), 
	.A1(n5185));
   OAI22_X1 U2471 (.ZN(U495_Z_0), 
	.B2(n17022), 
	.B1(n2725), 
	.A2(n17018), 
	.A1(FE_PHN2479_n5116));
   OAI22_X1 U2472 (.ZN(U494_Z_0), 
	.B2(n17017), 
	.B1(n2725), 
	.A2(n17013), 
	.A1(FE_PHN2474_n5214));
   OAI22_X1 U2473 (.ZN(U493_Z_0), 
	.B2(n17046), 
	.B1(n2725), 
	.A2(n17043), 
	.A1(n5321));
   OAI22_X1 U2474 (.ZN(U492_Z_0), 
	.B2(n17052), 
	.B1(n2725), 
	.A2(FE_OFN656_n17048), 
	.A1(FE_PHN2498_n5350));
   OAI22_X1 U2475 (.ZN(U491_Z_0), 
	.B2(n17057), 
	.B1(n2725), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2485_n5379));
   OAI22_X1 U2476 (.ZN(U490_Z_0), 
	.B2(n17062), 
	.B1(n2725), 
	.A2(FE_OFN663_n17058), 
	.A1(n5408));
   OAI22_X1 U2477 (.ZN(U489_Z_0), 
	.B2(n17067), 
	.B1(n2725), 
	.A2(n17063), 
	.A1(FE_PHN2747_n5437));
   OAI22_X1 U2478 (.ZN(U488_Z_0), 
	.B2(n17071), 
	.B1(n2725), 
	.A2(n17068), 
	.A1(FE_PHN2694_n5466));
   OAI22_X1 U2479 (.ZN(U487_Z_0), 
	.B2(FE_OFN666_n17077), 
	.B1(n2725), 
	.A2(n17074), 
	.A1(FE_PHN2728_n5115));
   OAI22_X1 U2480 (.ZN(U486_Z_0), 
	.B2(n17082), 
	.B1(n2725), 
	.A2(n17078), 
	.A1(FE_PHN2461_n5490));
   AOI222_X1 U2482 (.ZN(n2726), 
	.C2(FE_OFN208_n2015), 
	.C1(n16668), 
	.B2(n2728), 
	.B1(n2727), 
	.A2(n21), 
	.A1(n17008));
   NAND3_X1 U2483 (.ZN(n2728), 
	.A3(n5815), 
	.A2(n1651), 
	.A1(n2131));
   OAI21_X1 U2484 (.ZN(n2727), 
	.B2(n1687), 
	.B1(n16992), 
	.A(n2729));
   OAI21_X1 U2485 (.ZN(n2729), 
	.B2(n1651), 
	.B1(n16994), 
	.A(n5815));
   AOI221_X1 U2487 (.ZN(n2730), 
	.C2(n2731), 
	.C1(n2198), 
	.B2(n21), 
	.B1(n16989), 
	.A(n2732));
   INV_X1 U2488 (.ZN(n1687), 
	.A(n1651));
   NAND4_X1 U2489 (.ZN(n1651), 
	.A4(n2736), 
	.A3(n2735), 
	.A2(n2734), 
	.A1(n2733));
   AOI222_X1 U2490 (.ZN(n2736), 
	.C2(vis_psp_o[19]), 
	.C1(n16968), 
	.B2(n2738), 
	.B1(n16971), 
	.A2(vis_msp_o[19]), 
	.A1(n16974));
   AOI222_X1 U2492 (.ZN(n2735), 
	.C2(vis_r11_o[21]), 
	.C1(n16986), 
	.B2(vis_r12_o[21]), 
	.B1(n16965), 
	.A2(vis_r14_o[21]), 
	.A1(n16983));
   AOI222_X1 U2495 (.ZN(n2734), 
	.C2(vis_r8_o[21]), 
	.C1(n16959), 
	.B2(vis_r10_o[21]), 
	.B1(n16962), 
	.A2(vis_r9_o[21]), 
	.A1(n16980));
   AOI22_X1 U2497 (.ZN(n2733), 
	.B2(n2746), 
	.B1(n16955), 
	.A2(n2714), 
	.A1(FE_OFN646_n16977));
   AOI221_X1 U2499 (.ZN(n58), 
	.C2(n2411), 
	.C1(n2721), 
	.B2(n2410), 
	.B1(n2720), 
	.A(n2747));
   INV_X1 U2500 (.ZN(n2747), 
	.A(n2748));
   AOI22_X1 U2501 (.ZN(n2748), 
	.B2(n2749), 
	.B1(n2414), 
	.A2(FE_PHN748_n2415), 
	.A1(n2074));
   OAI22_X1 U2502 (.ZN(U483_Z_0), 
	.B2(n17005), 
	.B1(n2750), 
	.A2(n17001), 
	.A1(FE_PHN2515_n5617));
   OAI22_X1 U2503 (.ZN(U482_Z_0), 
	.B2(n17000), 
	.B1(n2750), 
	.A2(n16996), 
	.A1(FE_PHN2733_n5616));
   OAI22_X1 U2504 (.ZN(U481_Z_0), 
	.B2(n17042), 
	.B1(n2750), 
	.A2(n17038), 
	.A1(n5615));
   OAI22_X1 U2505 (.ZN(U480_Z_0), 
	.B2(n17037), 
	.B1(n2750), 
	.A2(FE_OFN652_n17033), 
	.A1(FE_PHN2448_n5614));
   OAI22_X1 U2506 (.ZN(U479_Z_0), 
	.B2(n17031), 
	.B1(n2750), 
	.A2(n17028), 
	.A1(n5613));
   OAI22_X1 U2507 (.ZN(U478_Z_0), 
	.B2(n17027), 
	.B1(n2750), 
	.A2(n17023), 
	.A1(FE_PHN2780_n5612));
   OAI22_X1 U2508 (.ZN(U477_Z_0), 
	.B2(n17022), 
	.B1(n2750), 
	.A2(n17018), 
	.A1(FE_PHN2492_n5611));
   OAI22_X1 U2509 (.ZN(U476_Z_0), 
	.B2(n17017), 
	.B1(n2750), 
	.A2(n17013), 
	.A1(FE_PHN2514_n5610));
   OAI22_X1 U2510 (.ZN(U475_Z_0), 
	.B2(n17046), 
	.B1(n2750), 
	.A2(n17043), 
	.A1(n5609));
   OAI22_X1 U2511 (.ZN(U474_Z_0), 
	.B2(n17052), 
	.B1(n2750), 
	.A2(FE_OFN656_n17048), 
	.A1(FE_PHN2459_n5608));
   OAI22_X1 U2512 (.ZN(U473_Z_0), 
	.B2(n17057), 
	.B1(n2750), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2487_n5607));
   OAI22_X1 U2513 (.ZN(U472_Z_0), 
	.B2(n17062), 
	.B1(n2750), 
	.A2(FE_OFN663_n17058), 
	.A1(FE_PHN2678_n5606));
   OAI22_X1 U2514 (.ZN(U471_Z_0), 
	.B2(n17067), 
	.B1(n2750), 
	.A2(n17063), 
	.A1(n5605));
   OAI22_X1 U2515 (.ZN(U470_Z_0), 
	.B2(n17071), 
	.B1(n2750), 
	.A2(n17068), 
	.A1(FE_PHN2779_n5604));
   OAI22_X1 U2516 (.ZN(U469_Z_0), 
	.B2(FE_OFN666_n17077), 
	.B1(n2750), 
	.A2(n17074), 
	.A1(FE_PHN2787_n5603));
   OAI22_X1 U2517 (.ZN(U468_Z_0), 
	.B2(n17082), 
	.B1(n2750), 
	.A2(n17078), 
	.A1(FE_PHN2497_n5602));
   AOI221_X1 U2519 (.ZN(n2753), 
	.C2(FE_OFN208_n2015), 
	.C1(n16706), 
	.B2(n20), 
	.B1(n17008), 
	.A(n2754));
   INV_X1 U2520 (.ZN(n2754), 
	.A(n2284));
   OAI221_X1 U2521 (.ZN(n2284), 
	.C2(n2127), 
	.C1(n5814), 
	.B2(n2755), 
	.B1(n2126), 
	.A(n1653));
   INV_X1 U2522 (.ZN(n2755), 
	.A(n5814));
   INV_X1 U2523 (.ZN(n2752), 
	.A(n55));
   OAI221_X1 U2524 (.ZN(n55), 
	.C2(n2596), 
	.C1(n2724), 
	.B2(n2757), 
	.B1(n2756), 
	.A(n2758));
   AOI22_X1 U2525 (.ZN(n2758), 
	.B2(n2721), 
	.B1(n2075), 
	.A2(n2068), 
	.A1(n2074));
   NAND3_X1 U2526 (.ZN(n2751), 
	.A3(n1688), 
	.A2(n16994), 
	.A1(n5814));
   INV_X1 U2527 (.ZN(n1688), 
	.A(n1653));
   NAND4_X1 U2528 (.ZN(n1653), 
	.A4(n2762), 
	.A3(n2761), 
	.A2(n2760), 
	.A1(n2759));
   AOI222_X1 U2529 (.ZN(n2762), 
	.C2(vis_psp_o[18]), 
	.C1(n16968), 
	.B2(n2764), 
	.B1(n16971), 
	.A2(vis_msp_o[18]), 
	.A1(n16974));
   AOI222_X1 U2531 (.ZN(n2761), 
	.C2(vis_r11_o[20]), 
	.C1(n16986), 
	.B2(vis_r12_o[20]), 
	.B1(n16965), 
	.A2(vis_r14_o[20]), 
	.A1(n16983));
   AOI222_X1 U2534 (.ZN(n2760), 
	.C2(vis_r8_o[20]), 
	.C1(n16959), 
	.B2(vis_r10_o[20]), 
	.B1(n16962), 
	.A2(vis_r9_o[20]), 
	.A1(n16980));
   AOI22_X1 U2536 (.ZN(n2759), 
	.B2(n2772), 
	.B1(n16955), 
	.A2(n2746), 
	.A1(FE_OFN646_n16977));
   XOR2_X1 U2538 (.Z(n5814), 
	.B(n2773), 
	.A(n16990));
   AOI221_X1 U2539 (.ZN(n2773), 
	.C2(n2774), 
	.C1(n2198), 
	.B2(n20), 
	.B1(n16989), 
	.A(n2732));
   OAI22_X1 U2540 (.ZN(U467_Z_0), 
	.B2(n17005), 
	.B1(n2775), 
	.A2(n17001), 
	.A1(FE_PHN2593_n5638));
   OAI22_X1 U2541 (.ZN(U466_Z_0), 
	.B2(n17000), 
	.B1(n2775), 
	.A2(n16996), 
	.A1(n5637));
   OAI22_X1 U2542 (.ZN(U465_Z_0), 
	.B2(n17042), 
	.B1(n2775), 
	.A2(n17038), 
	.A1(FE_PHN2732_n5636));
   OAI22_X1 U2543 (.ZN(U464_Z_0), 
	.B2(n17037), 
	.B1(n2775), 
	.A2(FE_OFN652_n17033), 
	.A1(FE_PHN2457_n5635));
   OAI22_X1 U2544 (.ZN(U463_Z_0), 
	.B2(n17031), 
	.B1(n2775), 
	.A2(n17028), 
	.A1(n5090));
   OAI22_X1 U2545 (.ZN(U462_Z_0), 
	.B2(n17027), 
	.B1(n2775), 
	.A2(n17023), 
	.A1(FE_PHN2766_n5186));
   OAI22_X1 U2546 (.ZN(U461_Z_0), 
	.B2(n17022), 
	.B1(n2775), 
	.A2(n17018), 
	.A1(FE_PHN2471_n5089));
   OAI22_X1 U2547 (.ZN(U460_Z_0), 
	.B2(n17017), 
	.B1(n2775), 
	.A2(n17013), 
	.A1(FE_PHN2475_n5215));
   OAI22_X1 U2548 (.ZN(U459_Z_0), 
	.B2(n17046), 
	.B1(n2775), 
	.A2(n17043), 
	.A1(n5322));
   OAI22_X1 U2549 (.ZN(U458_Z_0), 
	.B2(n17052), 
	.B1(n2775), 
	.A2(FE_OFN656_n17048), 
	.A1(FE_PHN2469_n5351));
   OAI22_X1 U2550 (.ZN(U457_Z_0), 
	.B2(n17057), 
	.B1(n2775), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2477_n5380));
   OAI22_X1 U2551 (.ZN(U456_Z_0), 
	.B2(n17062), 
	.B1(n2775), 
	.A2(FE_OFN663_n17058), 
	.A1(FE_PHN2629_n5409));
   OAI22_X1 U2552 (.ZN(U455_Z_0), 
	.B2(n17067), 
	.B1(n2775), 
	.A2(n17063), 
	.A1(FE_PHN2717_n5438));
   OAI22_X1 U2553 (.ZN(U454_Z_0), 
	.B2(n17071), 
	.B1(n2775), 
	.A2(n17068), 
	.A1(n5467));
   OAI22_X1 U2554 (.ZN(U453_Z_0), 
	.B2(FE_OFN666_n17077), 
	.B1(n2775), 
	.A2(n17074), 
	.A1(n5088));
   OAI22_X1 U2555 (.ZN(U452_Z_0), 
	.B2(n17082), 
	.B1(n2775), 
	.A2(n17078), 
	.A1(FE_PHN2542_n5491));
   AOI222_X1 U2557 (.ZN(n2777), 
	.C2(FE_OFN208_n2015), 
	.C1(n16709), 
	.B2(n2779), 
	.B1(n2778), 
	.A2(n22), 
	.A1(n17008));
   NAND3_X1 U2558 (.ZN(n2779), 
	.A3(n5813), 
	.A2(n2156), 
	.A1(n2131));
   OAI21_X1 U2559 (.ZN(n2778), 
	.B2(n1654), 
	.B1(n16992), 
	.A(n2780));
   OAI21_X1 U2560 (.ZN(n2780), 
	.B2(n2156), 
	.B1(n16994), 
	.A(n5813));
   XOR2_X1 U2561 (.Z(n5813), 
	.B(n2781), 
	.A(n16990));
   AOI221_X1 U2562 (.ZN(n2781), 
	.C2(n486), 
	.C1(n2198), 
	.B2(n22), 
	.B1(n16989), 
	.A(n2732));
   INV_X1 U2563 (.ZN(n1654), 
	.A(n2156));
   NAND4_X1 U2564 (.ZN(n2156), 
	.A4(n2785), 
	.A3(n2784), 
	.A2(n2783), 
	.A1(n2782));
   AOI222_X1 U2565 (.ZN(n2785), 
	.C2(vis_psp_o[17]), 
	.C1(n16968), 
	.B2(n2787), 
	.B1(n16971), 
	.A2(vis_msp_o[17]), 
	.A1(n16974));
   AOI222_X1 U2567 (.ZN(n2784), 
	.C2(vis_r11_o[19]), 
	.C1(n16986), 
	.B2(vis_r12_o[19]), 
	.B1(n16965), 
	.A2(vis_r14_o[19]), 
	.A1(n16983));
   AOI222_X1 U2570 (.ZN(n2783), 
	.C2(vis_r8_o[19]), 
	.C1(n16959), 
	.B2(vis_r10_o[19]), 
	.B1(n16962), 
	.A2(vis_r9_o[19]), 
	.A1(n16980));
   AOI22_X1 U2572 (.ZN(n2782), 
	.B2(n2795), 
	.B1(n16955), 
	.A2(n2772), 
	.A1(FE_OFN646_n16977));
   INV_X1 U2574 (.ZN(n2776), 
	.A(n70));
   OAI221_X1 U2575 (.ZN(n70), 
	.C2(n2419), 
	.C1(n2724), 
	.B2(n2418), 
	.B1(n2756), 
	.A(n2796));
   AOI22_X1 U2576 (.ZN(n2796), 
	.B2(n2721), 
	.B1(FE_PHN728_n2421), 
	.A2(n2422), 
	.A1(n2074));
   OAI22_X1 U2577 (.ZN(U449_Z_0), 
	.B2(n17005), 
	.B1(n2797), 
	.A2(n17001), 
	.A1(FE_PHN2491_n5066));
   OAI22_X1 U2578 (.ZN(U448_Z_0), 
	.B2(n17000), 
	.B1(n2797), 
	.A2(n16996), 
	.A1(n5065));
   OAI22_X1 U2579 (.ZN(U447_Z_0), 
	.B2(n17042), 
	.B1(n2797), 
	.A2(n17038), 
	.A1(FE_PHN2791_n5297));
   OAI22_X1 U2580 (.ZN(U446_Z_0), 
	.B2(n17037), 
	.B1(n2797), 
	.A2(FE_OFN652_n17033), 
	.A1(FE_PHN2486_n5276));
   OAI22_X1 U2581 (.ZN(U445_Z_0), 
	.B2(n17031), 
	.B1(n2797), 
	.A2(n17028), 
	.A1(n5064));
   OAI22_X1 U2582 (.ZN(U444_Z_0), 
	.B2(n17027), 
	.B1(n2797), 
	.A2(n17023), 
	.A1(FE_PHN2752_n5187));
   OAI22_X1 U2583 (.ZN(U443_Z_0), 
	.B2(n17022), 
	.B1(n2797), 
	.A2(n17018), 
	.A1(FE_PHN2540_n5063));
   OAI22_X1 U2584 (.ZN(U442_Z_0), 
	.B2(n17017), 
	.B1(n2797), 
	.A2(n17013), 
	.A1(FE_PHN2500_n5216));
   OAI22_X1 U2585 (.ZN(U441_Z_0), 
	.B2(n17046), 
	.B1(n2797), 
	.A2(n17043), 
	.A1(n5323));
   OAI22_X1 U2586 (.ZN(U440_Z_0), 
	.B2(n17052), 
	.B1(n2797), 
	.A2(FE_OFN656_n17048), 
	.A1(FE_PHN2482_n5352));
   OAI22_X1 U2587 (.ZN(U439_Z_0), 
	.B2(n17057), 
	.B1(n2797), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2525_n5381));
   OAI22_X1 U2588 (.ZN(U438_Z_0), 
	.B2(n17062), 
	.B1(n2797), 
	.A2(FE_OFN663_n17058), 
	.A1(FE_PHN2665_n5410));
   OAI22_X1 U2589 (.ZN(U437_Z_0), 
	.B2(n17067), 
	.B1(n2797), 
	.A2(n17063), 
	.A1(FE_PHN2698_n5439));
   OAI22_X1 U2590 (.ZN(U436_Z_0), 
	.B2(n17071), 
	.B1(n2797), 
	.A2(n17068), 
	.A1(FE_PHN2771_n5468));
   OAI22_X1 U2591 (.ZN(U435_Z_0), 
	.B2(FE_OFN666_n17077), 
	.B1(n2797), 
	.A2(n17074), 
	.A1(FE_PHN2788_n5062));
   OAI22_X1 U2592 (.ZN(U434_Z_0), 
	.B2(n17082), 
	.B1(n2797), 
	.A2(n17078), 
	.A1(FE_PHN2467_n5492));
   AOI221_X1 U2594 (.ZN(n2799), 
	.C2(FE_OFN208_n2015), 
	.C1(n16672), 
	.B2(n2249), 
	.B1(n17008), 
	.A(n2289));
   AND2_X1 U2595 (.ZN(n2289), 
	.A2(n1657), 
	.A1(n2800));
   OAI22_X1 U2596 (.ZN(n2800), 
	.B2(n2801), 
	.B1(n2131), 
	.A2(n5812), 
	.A1(n16992));
   INV_X1 U2597 (.ZN(n2801), 
	.A(n5812));
   AOI221_X1 U2598 (.ZN(n64), 
	.C2(n2469), 
	.C1(n2720), 
	.B2(n2074), 
	.B1(n2464), 
	.A(n2802));
   INV_X1 U2599 (.ZN(n2802), 
	.A(n2803));
   AOI22_X1 U2600 (.ZN(n2803), 
	.B2(n2721), 
	.B1(FE_PHN679_n2465), 
	.A2(n2749), 
	.A1(n2468));
   NAND3_X1 U2601 (.ZN(n2798), 
	.A3(n1690), 
	.A2(n16994), 
	.A1(n5812));
   INV_X1 U2602 (.ZN(n1690), 
	.A(n1657));
   NAND4_X1 U2603 (.ZN(n1657), 
	.A4(n2807), 
	.A3(n2806), 
	.A2(n2805), 
	.A1(n2804));
   AOI222_X1 U2604 (.ZN(n2807), 
	.C2(vis_psp_o[16]), 
	.C1(n16968), 
	.B2(n2809), 
	.B1(n16971), 
	.A2(vis_msp_o[16]), 
	.A1(n16974));
   AOI222_X1 U2606 (.ZN(n2806), 
	.C2(vis_r11_o[18]), 
	.C1(n16986), 
	.B2(vis_r12_o[18]), 
	.B1(n16965), 
	.A2(vis_r14_o[18]), 
	.A1(n16983));
   AOI222_X1 U2609 (.ZN(n2805), 
	.C2(vis_r8_o[18]), 
	.C1(n16959), 
	.B2(vis_r10_o[18]), 
	.B1(n16962), 
	.A2(vis_r9_o[18]), 
	.A1(n16980));
   AOI22_X1 U2611 (.ZN(n2804), 
	.B2(n2817), 
	.B1(n16955), 
	.A2(n2795), 
	.A1(FE_OFN646_n16977));
   XOR2_X1 U2613 (.Z(n5812), 
	.B(n2818), 
	.A(n16990));
   AOI221_X1 U2614 (.ZN(n2818), 
	.C2(n2819), 
	.C1(n2198), 
	.B2(n2249), 
	.B1(n16989), 
	.A(n2732));
   OAI22_X1 U2615 (.ZN(U433_Z_0), 
	.B2(n17005), 
	.B1(n2820), 
	.A2(n17001), 
	.A1(FE_PHN2489_n5087));
   OAI22_X1 U2616 (.ZN(U432_Z_0), 
	.B2(n17000), 
	.B1(n2820), 
	.A2(n16996), 
	.A1(FE_PHN2727_n5086));
   OAI22_X1 U2617 (.ZN(U431_Z_0), 
	.B2(n17042), 
	.B1(n2820), 
	.A2(n17038), 
	.A1(FE_PHN2652_n5298));
   OAI22_X1 U2618 (.ZN(U430_Z_0), 
	.B2(n17037), 
	.B1(n2820), 
	.A2(FE_OFN652_n17033), 
	.A1(FE_PHN2481_n5277));
   OAI22_X1 U2619 (.ZN(U429_Z_0), 
	.B2(n17031), 
	.B1(n2820), 
	.A2(n17028), 
	.A1(n5085));
   OAI22_X1 U2620 (.ZN(U428_Z_0), 
	.B2(n17027), 
	.B1(n2820), 
	.A2(n17023), 
	.A1(n5188));
   OAI22_X1 U2621 (.ZN(U427_Z_0), 
	.B2(n17022), 
	.B1(n2820), 
	.A2(n17018), 
	.A1(FE_PHN2507_n5084));
   OAI22_X1 U2622 (.ZN(U426_Z_0), 
	.B2(n17017), 
	.B1(n2820), 
	.A2(n17013), 
	.A1(FE_PHN2543_n5217));
   OAI22_X1 U2623 (.ZN(U425_Z_0), 
	.B2(n17046), 
	.B1(n2820), 
	.A2(n17043), 
	.A1(n5324));
   OAI22_X1 U2624 (.ZN(U424_Z_0), 
	.B2(n17052), 
	.B1(n2820), 
	.A2(FE_OFN656_n17048), 
	.A1(FE_PHN2458_n5353));
   OAI22_X1 U2625 (.ZN(U423_Z_0), 
	.B2(n17057), 
	.B1(n2820), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2470_n5382));
   OAI22_X1 U2626 (.ZN(U422_Z_0), 
	.B2(n17062), 
	.B1(n2820), 
	.A2(FE_OFN663_n17058), 
	.A1(FE_PHN2654_n5411));
   OAI22_X1 U2627 (.ZN(U421_Z_0), 
	.B2(n17067), 
	.B1(n2820), 
	.A2(n17063), 
	.A1(FE_PHN2646_n5440));
   OAI22_X1 U2628 (.ZN(U420_Z_0), 
	.B2(n17071), 
	.B1(n2820), 
	.A2(n17068), 
	.A1(FE_PHN2738_n5469));
   OAI22_X1 U2629 (.ZN(U419_Z_0), 
	.B2(FE_OFN666_n17077), 
	.B1(n2820), 
	.A2(n17074), 
	.A1(FE_PHN2774_n5083));
   OAI22_X1 U2630 (.ZN(U418_Z_0), 
	.B2(n17082), 
	.B1(n2820), 
	.A2(n17078), 
	.A1(FE_PHN2466_n5493));
   AOI222_X1 U2632 (.ZN(n2822), 
	.C2(FE_OFN208_n2015), 
	.C1(n16710), 
	.B2(n2824), 
	.B1(n2823), 
	.A2(n2258), 
	.A1(n17008));
   NAND3_X1 U2633 (.ZN(n2824), 
	.A3(n5811), 
	.A2(n1658), 
	.A1(n2131));
   OAI21_X1 U2634 (.ZN(n2823), 
	.B2(n1691), 
	.B1(n16992), 
	.A(n2825));
   OAI21_X1 U2635 (.ZN(n2825), 
	.B2(n1658), 
	.B1(n16994), 
	.A(n5811));
   XOR2_X1 U2636 (.Z(n5811), 
	.B(n2826), 
	.A(n16990));
   AOI221_X1 U2637 (.ZN(n2826), 
	.C2(n2827), 
	.C1(n2198), 
	.B2(n2258), 
	.B1(n16989), 
	.A(n2732));
   INV_X1 U2638 (.ZN(n1691), 
	.A(n1658));
   NAND4_X1 U2639 (.ZN(n1658), 
	.A4(n2831), 
	.A3(n2830), 
	.A2(n2829), 
	.A1(n2828));
   AOI222_X1 U2640 (.ZN(n2831), 
	.C2(vis_psp_o[15]), 
	.C1(n16968), 
	.B2(n2833), 
	.B1(n16971), 
	.A2(vis_msp_o[15]), 
	.A1(n16974));
   AOI222_X1 U2642 (.ZN(n2830), 
	.C2(vis_r11_o[17]), 
	.C1(n16986), 
	.B2(vis_r12_o[17]), 
	.B1(n16965), 
	.A2(vis_r14_o[17]), 
	.A1(n16983));
   AOI222_X1 U2645 (.ZN(n2829), 
	.C2(vis_r8_o[17]), 
	.C1(n16959), 
	.B2(vis_r10_o[17]), 
	.B1(n16962), 
	.A2(vis_r9_o[17]), 
	.A1(n16980));
   AOI22_X1 U2647 (.ZN(n2828), 
	.B2(n2841), 
	.B1(n16955), 
	.A2(n2817), 
	.A1(FE_OFN646_n16977));
   INV_X1 U2649 (.ZN(n2821), 
	.A(n66));
   OAI221_X1 U2650 (.ZN(n66), 
	.C2(n2473), 
	.C1(n2724), 
	.B2(n2472), 
	.B1(n2756), 
	.A(n2842));
   AOI22_X1 U2651 (.ZN(n2842), 
	.B2(n2721), 
	.B1(n2003), 
	.A2(n2005), 
	.A1(n2074));
   OAI22_X1 U2652 (.ZN(U415_Z_0), 
	.B2(n17005), 
	.B1(n2843), 
	.A2(n17001), 
	.A1(FE_PHN2438_n5073));
   OAI22_X1 U2653 (.ZN(U414_Z_0), 
	.B2(n17000), 
	.B1(n2843), 
	.A2(n16996), 
	.A1(FE_PHN2786_n5072));
   OAI22_X1 U2654 (.ZN(U413_Z_0), 
	.B2(n17042), 
	.B1(n2843), 
	.A2(n17038), 
	.A1(FE_PHN2769_n5299));
   OAI22_X1 U2655 (.ZN(U412_Z_0), 
	.B2(n17037), 
	.B1(n2843), 
	.A2(FE_OFN652_n17033), 
	.A1(FE_PHN2562_n5278));
   OAI22_X1 U2656 (.ZN(U411_Z_0), 
	.B2(n17031), 
	.B1(n2843), 
	.A2(n17028), 
	.A1(n5071));
   OAI22_X1 U2657 (.ZN(U410_Z_0), 
	.B2(n17027), 
	.B1(n2843), 
	.A2(n17023), 
	.A1(FE_PHN2647_n5189));
   OAI22_X1 U2658 (.ZN(U409_Z_0), 
	.B2(n17022), 
	.B1(n2843), 
	.A2(n17018), 
	.A1(FE_PHN2583_n5070));
   OAI22_X1 U2659 (.ZN(U408_Z_0), 
	.B2(FE_OFN648_n17017), 
	.B1(n2843), 
	.A2(n17013), 
	.A1(FE_PHN2553_n5218));
   OAI22_X1 U2660 (.ZN(U407_Z_0), 
	.B2(n17046), 
	.B1(n2843), 
	.A2(n17043), 
	.A1(n5325));
   OAI22_X1 U2661 (.ZN(U406_Z_0), 
	.B2(n17052), 
	.B1(n2843), 
	.A2(FE_OFN656_n17048), 
	.A1(FE_PHN2463_n5354));
   OAI22_X1 U2662 (.ZN(U405_Z_0), 
	.B2(n17057), 
	.B1(n2843), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2547_n5383));
   OAI22_X1 U2663 (.ZN(U404_Z_0), 
	.B2(n17062), 
	.B1(n2843), 
	.A2(FE_OFN663_n17058), 
	.A1(FE_PHN2651_n5412));
   OAI22_X1 U2664 (.ZN(U403_Z_0), 
	.B2(n17067), 
	.B1(n2843), 
	.A2(n17063), 
	.A1(FE_PHN2641_n5441));
   OAI22_X1 U2665 (.ZN(U402_Z_0), 
	.B2(n17071), 
	.B1(n2843), 
	.A2(n17068), 
	.A1(FE_PHN2775_n5470));
   OAI22_X1 U2666 (.ZN(U401_Z_0), 
	.B2(FE_OFN666_n17077), 
	.B1(n2843), 
	.A2(n17074), 
	.A1(FE_PHN2700_n5069));
   OAI22_X1 U2667 (.ZN(U400_Z_0), 
	.B2(n17082), 
	.B1(n2843), 
	.A2(n17078), 
	.A1(FE_PHN2480_n5494));
   AOI221_X1 U2669 (.ZN(n2846), 
	.C2(FE_OFN208_n2015), 
	.C1(n16711), 
	.B2(n17), 
	.B1(n17008), 
	.A(n2847));
   INV_X1 U2670 (.ZN(n2847), 
	.A(n2307));
   NAND2_X1 U2671 (.ZN(n2307), 
	.A2(n1660), 
	.A1(n2848));
   OAI22_X1 U2672 (.ZN(n2848), 
	.B2(n2849), 
	.B1(n2131), 
	.A2(n5810), 
	.A1(n16992));
   INV_X1 U2673 (.ZN(n2849), 
	.A(n5810));
   INV_X1 U2674 (.ZN(n2845), 
	.A(n68));
   OAI221_X1 U2675 (.ZN(n68), 
	.C2(FE_PHN685_n2516), 
	.C1(n2724), 
	.B2(n2723), 
	.B1(n2517), 
	.A(n2850));
   AOI22_X1 U2676 (.ZN(n2850), 
	.B2(n2721), 
	.B1(n2019), 
	.A2(n2720), 
	.A1(n2023));
   INV_X1 U2677 (.ZN(n2724), 
	.A(n2749));
   NAND3_X1 U2678 (.ZN(n2844), 
	.A3(n1692), 
	.A2(n16994), 
	.A1(n5810));
   INV_X1 U2679 (.ZN(n1692), 
	.A(n1660));
   NAND4_X1 U2680 (.ZN(n1660), 
	.A4(n2854), 
	.A3(n2853), 
	.A2(n2852), 
	.A1(n2851));
   AOI222_X1 U2681 (.ZN(n2854), 
	.C2(vis_psp_o[14]), 
	.C1(n16968), 
	.B2(n2856), 
	.B1(n16971), 
	.A2(vis_msp_o[14]), 
	.A1(n16974));
   AOI222_X1 U2683 (.ZN(n2853), 
	.C2(vis_r11_o[16]), 
	.C1(n16986), 
	.B2(vis_r12_o[16]), 
	.B1(n16965), 
	.A2(vis_r14_o[16]), 
	.A1(n16983));
   AOI222_X1 U2686 (.ZN(n2852), 
	.C2(vis_r8_o[16]), 
	.C1(n16959), 
	.B2(vis_r10_o[16]), 
	.B1(n16963), 
	.A2(vis_r9_o[16]), 
	.A1(n16980));
   AOI22_X1 U2688 (.ZN(n2851), 
	.B2(n1163), 
	.B1(n16955), 
	.A2(n2841), 
	.A1(FE_OFN646_n16977));
   XOR2_X1 U2690 (.Z(n5810), 
	.B(n2864), 
	.A(n16990));
   AOI221_X1 U2691 (.ZN(n2864), 
	.C2(n2865), 
	.C1(n2198), 
	.B2(n17), 
	.B1(n16989), 
	.A(n2732));
   NOR2_X1 U2692 (.ZN(n2696), 
	.A2(FE_OFN383_n71), 
	.A1(n2055));
   OAI22_X1 U2693 (.ZN(U399_Z_0), 
	.B2(n17005), 
	.B1(n2866), 
	.A2(n17001), 
	.A1(FE_PHN2581_n5107));
   OAI22_X1 U2694 (.ZN(U398_Z_0), 
	.B2(n17000), 
	.B1(n2866), 
	.A2(n16996), 
	.A1(FE_PHN2666_n5106));
   OAI22_X1 U2695 (.ZN(U397_Z_0), 
	.B2(n17042), 
	.B1(n2866), 
	.A2(n17038), 
	.A1(FE_PHN2718_n5300));
   OAI22_X1 U2696 (.ZN(U396_Z_0), 
	.B2(n17037), 
	.B1(n2866), 
	.A2(n17033), 
	.A1(FE_PHN2527_n5279));
   OAI22_X1 U2697 (.ZN(U395_Z_0), 
	.B2(n17031), 
	.B1(n2866), 
	.A2(n17028), 
	.A1(n5105));
   OAI22_X1 U2698 (.ZN(U394_Z_0), 
	.B2(n17027), 
	.B1(n2866), 
	.A2(n17023), 
	.A1(FE_PHN2693_n5190));
   OAI22_X1 U2699 (.ZN(U393_Z_0), 
	.B2(n17022), 
	.B1(n2866), 
	.A2(n17018), 
	.A1(FE_PHN2511_n5104));
   OAI22_X1 U2700 (.ZN(U392_Z_0), 
	.B2(n17017), 
	.B1(n2866), 
	.A2(n17013), 
	.A1(FE_PHN2592_n5219));
   OAI22_X1 U2701 (.ZN(U391_Z_0), 
	.B2(n17046), 
	.B1(n2866), 
	.A2(n17043), 
	.A1(n5326));
   OAI22_X1 U2702 (.ZN(U390_Z_0), 
	.B2(n17052), 
	.B1(n2866), 
	.A2(n17048), 
	.A1(FE_PHN2571_n5355));
   OAI22_X1 U2703 (.ZN(U389_Z_0), 
	.B2(n17057), 
	.B1(n2866), 
	.A2(n17053), 
	.A1(FE_PHN2605_n5384));
   OAI22_X1 U2704 (.ZN(U388_Z_0), 
	.B2(n17062), 
	.B1(n2866), 
	.A2(n17058), 
	.A1(FE_PHN2601_n5413));
   OAI22_X1 U2705 (.ZN(U387_Z_0), 
	.B2(n17067), 
	.B1(n2866), 
	.A2(n17063), 
	.A1(FE_PHN2714_n5442));
   OAI22_X1 U2706 (.ZN(U386_Z_0), 
	.B2(n17071), 
	.B1(n2866), 
	.A2(n17068), 
	.A1(n5471));
   OAI22_X1 U2707 (.ZN(U385_Z_0), 
	.B2(n17077), 
	.B1(n2866), 
	.A2(n17074), 
	.A1(FE_PHN2736_n5103));
   OAI22_X1 U2708 (.ZN(U384_Z_0), 
	.B2(n17082), 
	.B1(n2866), 
	.A2(n17078), 
	.A1(FE_PHN2442_n5495));
   AOI221_X1 U2710 (.ZN(n2867), 
	.C2(n2253), 
	.C1(n17008), 
	.B2(FE_OFN2_n2015), 
	.B1(n16658), 
	.A(n135));
   OAI221_X1 U2711 (.ZN(n135), 
	.C2(n2088), 
	.C1(n2869), 
	.B2(n2090), 
	.B1(n2868), 
	.A(n2870));
   AOI221_X1 U2712 (.ZN(n2870), 
	.C2(n2872), 
	.C1(n2094), 
	.B2(n2871), 
	.B1(n2093), 
	.A(n2873));
   OAI211_X1 U2713 (.ZN(n2094), 
	.C2(n2875), 
	.C1(n2874), 
	.B(n2877), 
	.A(n2876));
   AOI222_X1 U2714 (.ZN(n2877), 
	.C2(n2881), 
	.C1(n16787), 
	.B2(n2879), 
	.B1(hrdata_i[22]), 
	.A2(n2878), 
	.A1(sub_2068_A_22_));
   AOI22_X1 U2716 (.ZN(n2876), 
	.B2(n2344), 
	.B1(n16645), 
	.A2(n2883), 
	.A1(n2882));
   OAI221_X1 U2717 (.ZN(n2883), 
	.C2(n2886), 
	.C1(n5053), 
	.B2(n2885), 
	.B1(n1896), 
	.A(n2887));
   AOI222_X1 U2718 (.ZN(n2887), 
	.C2(n2890), 
	.C1(n1887), 
	.B2(n2889), 
	.B1(n1191), 
	.A2(n2888), 
	.A1(n1890));
   NAND4_X1 U2720 (.ZN(n2093), 
	.A4(n2894), 
	.A3(n2893), 
	.A2(FE_PHN780_n2892), 
	.A1(n2891));
   AOI221_X1 U2721 (.ZN(n2894), 
	.C2(n2896), 
	.C1(n2882), 
	.B2(n2895), 
	.B1(n407), 
	.A(n2897));
   OAI221_X1 U2722 (.ZN(n2896), 
	.C2(n2899), 
	.C1(n5157), 
	.B2(n2898), 
	.B1(n5151), 
	.A(n2900));
   AOI22_X1 U2723 (.ZN(n2900), 
	.B2(n2902), 
	.B1(n1893), 
	.A2(n2901), 
	.A1(n1897));
   INV_X1 U2724 (.ZN(n407), 
	.A(n426));
   OAI211_X1 U2725 (.ZN(n426), 
	.C2(n1372), 
	.C1(n2903), 
	.B(n2905), 
	.A(n2904));
   NAND3_X1 U2726 (.ZN(n2904), 
	.A3(n2907), 
	.A2(n1372), 
	.A1(n2906));
   OAI22_X1 U2727 (.ZN(n2906), 
	.B2(n2911), 
	.B1(n2910), 
	.A2(n2909), 
	.A1(n2908));
   AOI22_X1 U2728 (.ZN(n2893), 
	.B2(FE_OFN534_n2388), 
	.B1(n16645), 
	.A2(n2352), 
	.A1(n2912));
   AOI222_X1 U2729 (.ZN(n2892), 
	.C2(n2916), 
	.C1(n2915), 
	.B2(n2914), 
	.B1(n2913), 
	.A2(n2879), 
	.A1(hrdata_i[14]));
   AOI22_X1 U2730 (.ZN(n2891), 
	.B2(n2878), 
	.B1(sub_2068_A_14_), 
	.A2(n2917), 
	.A1(n16787));
   INV_X1 U2732 (.ZN(n2088), 
	.A(n2546));
   OAI211_X1 U2733 (.ZN(n2546), 
	.C2(FE_PHN2928_n1145), 
	.C1(n2918), 
	.B(n2920), 
	.A(n2919));
   AOI211_X1 U2734 (.ZN(n2920), 
	.C2(n2922), 
	.C1(n2921), 
	.B(n2897), 
	.A(n2923));
   AOI21_X1 U2735 (.ZN(n2923), 
	.B2(n2925), 
	.B1(n2924), 
	.A(n2926));
   AOI222_X1 U2736 (.ZN(n2925), 
	.C2(n2929), 
	.C1(n1191), 
	.B2(n1189), 
	.B1(n2928), 
	.A2(n2927), 
	.A1(n1887));
   NOR2_X1 U2737 (.ZN(n2928), 
	.A2(n2930), 
	.A1(n5503));
   AOI222_X1 U2738 (.ZN(n2924), 
	.C2(n2933), 
	.C1(n1897), 
	.B2(n2932), 
	.B1(n1890), 
	.A2(n2931), 
	.A1(n1893));
   INV_X1 U2739 (.ZN(n2921), 
	.A(n2373));
   OAI22_X1 U2740 (.ZN(n2373), 
	.B2(n2936), 
	.B1(n2935), 
	.A2(n2934), 
	.A1(n2313));
   INV_X1 U2741 (.ZN(n2936), 
	.A(n2934));
   AOI22_X1 U2742 (.ZN(n2935), 
	.B2(n16788), 
	.B1(n2938), 
	.A2(n2337), 
	.A1(n2937));
   INV_X1 U2743 (.ZN(n2938), 
	.A(FE_OFN525_n2332));
   AOI22_X1 U2744 (.ZN(n2934), 
	.B2(n2942), 
	.B1(n2941), 
	.A2(n2940), 
	.A1(n2939));
   INV_X1 U2745 (.ZN(n1145), 
	.A(hrdata_i[30]));
   INV_X1 U2746 (.ZN(n2090), 
	.A(n2545));
   NAND3_X1 U2747 (.ZN(n2545), 
	.A3(n2945), 
	.A2(n2944), 
	.A1(n2943));
   AOI221_X1 U2748 (.ZN(n2945), 
	.C2(n2878), 
	.C1(sub_2068_A_6_), 
	.B2(n2946), 
	.B1(n16787), 
	.A(n2947));
   OAI22_X1 U2749 (.ZN(n2947), 
	.B2(n2948), 
	.B1(n4798), 
	.A2(n397), 
	.A1(n2918));
   INV_X1 U2750 (.ZN(n397), 
	.A(hrdata_i[6]));
   AOI22_X1 U2752 (.ZN(n2944), 
	.B2(n2325), 
	.B1(n16645), 
	.A2(n2949), 
	.A1(n2882));
   OAI221_X1 U2753 (.ZN(n2949), 
	.C2(n2899), 
	.C1(n5518), 
	.B2(n2898), 
	.B1(n1885), 
	.A(n2950));
   AOI22_X1 U2754 (.ZN(n2950), 
	.B2(n2952), 
	.B1(n1893), 
	.A2(n2951), 
	.A1(n1897));
   AOI22_X1 U2756 (.ZN(n2943), 
	.B2(n2953), 
	.B1(n2913), 
	.A2(n2329), 
	.A1(n2912));
   INV_X1 U2757 (.ZN(n2868), 
	.A(n2954));
   NAND3_X1 U2758 (.ZN(n2285), 
	.A3(n1693), 
	.A2(n16994), 
	.A1(n5809));
   INV_X1 U2759 (.ZN(n1693), 
	.A(n1663));
   NAND2_X1 U2760 (.ZN(n2305), 
	.A2(n1663), 
	.A1(n2955));
   NAND4_X1 U2761 (.ZN(n1663), 
	.A4(n2959), 
	.A3(n2958), 
	.A2(n2957), 
	.A1(n2956));
   AOI222_X1 U2762 (.ZN(n2959), 
	.C2(vis_r9_o[14]), 
	.C1(n16979), 
	.B2(n2961), 
	.B1(n16976), 
	.A2(vis_r8_o[14]), 
	.A1(n16958));
   AOI222_X1 U2764 (.ZN(n2958), 
	.C2(vis_r14_o[14]), 
	.C1(n16984), 
	.B2(n2964), 
	.B1(n16970), 
	.A2(vis_r11_o[14]), 
	.A1(n16985));
   AOI222_X1 U2767 (.ZN(n2957), 
	.C2(vis_msp_o[12]), 
	.C1(n16975), 
	.B2(vis_r10_o[14]), 
	.B1(n16963), 
	.A2(vis_psp_o[12]), 
	.A1(n16967));
   AOI22_X1 U2769 (.ZN(n2956), 
	.B2(n16956), 
	.B1(n2970), 
	.A2(vis_r12_o[14]), 
	.A1(n16966));
   OAI22_X1 U2770 (.ZN(n2955), 
	.B2(n2971), 
	.B1(n2131), 
	.A2(n5809), 
	.A1(n16992));
   INV_X1 U2771 (.ZN(n2971), 
	.A(n5809));
   XOR2_X1 U2772 (.Z(n5809), 
	.B(n2972), 
	.A(n2169));
   AOI221_X1 U2773 (.ZN(n2972), 
	.C2(n795), 
	.C1(n2198), 
	.B2(n2253), 
	.B1(n16989), 
	.A(n2732));
   OAI22_X1 U2774 (.ZN(U383_Z_0), 
	.B2(n17005), 
	.B1(n2973), 
	.A2(n17001), 
	.A1(FE_PHN2510_n5599));
   OAI22_X1 U2775 (.ZN(U382_Z_0), 
	.B2(n17000), 
	.B1(n2973), 
	.A2(n16996), 
	.A1(FE_PHN2749_n5598));
   OAI22_X1 U2776 (.ZN(U381_Z_0), 
	.B2(n17042), 
	.B1(n2973), 
	.A2(n17038), 
	.A1(FE_PHN2743_n5597));
   OAI22_X1 U2777 (.ZN(U380_Z_0), 
	.B2(n17037), 
	.B1(n2973), 
	.A2(n17033), 
	.A1(FE_PHN2618_n5596));
   OAI22_X1 U2778 (.ZN(U379_Z_0), 
	.B2(n17031), 
	.B1(n2973), 
	.A2(n17028), 
	.A1(FE_PHN4896_n5134));
   OAI22_X1 U2779 (.ZN(U378_Z_0), 
	.B2(n17027), 
	.B1(n2973), 
	.A2(n17023), 
	.A1(FE_PHN2683_n5191));
   OAI22_X1 U2780 (.ZN(U377_Z_0), 
	.B2(n17022), 
	.B1(n2973), 
	.A2(n17018), 
	.A1(FE_PHN2530_n5133));
   OAI22_X1 U2781 (.ZN(U376_Z_0), 
	.B2(n17017), 
	.B1(n2973), 
	.A2(n17013), 
	.A1(FE_PHN2517_n5220));
   OAI22_X1 U2782 (.ZN(U375_Z_0), 
	.B2(n17046), 
	.B1(n2973), 
	.A2(n17043), 
	.A1(FE_PHN3609_n5327));
   OAI22_X1 U2783 (.ZN(U374_Z_0), 
	.B2(n17052), 
	.B1(n2973), 
	.A2(n17048), 
	.A1(FE_PHN2541_n5356));
   OAI22_X1 U2784 (.ZN(U373_Z_0), 
	.B2(n17057), 
	.B1(n2973), 
	.A2(n17053), 
	.A1(FE_PHN2505_n5385));
   OAI22_X1 U2785 (.ZN(U372_Z_0), 
	.B2(n17062), 
	.B1(n2973), 
	.A2(n17058), 
	.A1(FE_PHN2642_n5414));
   OAI22_X1 U2786 (.ZN(U371_Z_0), 
	.B2(n17067), 
	.B1(n2973), 
	.A2(n17063), 
	.A1(FE_PHN2594_n5443));
   OAI22_X1 U2787 (.ZN(U370_Z_0), 
	.B2(n17071), 
	.B1(n2973), 
	.A2(n17068), 
	.A1(FE_PHN2761_n5472));
   OAI22_X1 U2788 (.ZN(U369_Z_0), 
	.B2(n17077), 
	.B1(n2973), 
	.A2(n17074), 
	.A1(FE_PHN2662_n5132));
   OAI22_X1 U2789 (.ZN(U368_Z_0), 
	.B2(n17082), 
	.B1(n2973), 
	.A2(n17078), 
	.A1(FE_PHN2456_n5496));
   AOI221_X1 U2791 (.ZN(n2975), 
	.C2(n2259), 
	.C1(n17008), 
	.B2(FE_OFN2_n2015), 
	.B1(n16679), 
	.A(n2976));
   INV_X4 U2792 (.ZN(n2976), 
	.A(FE_OFN384_n118));
   AOI221_X1 U2793 (.ZN(n118), 
	.C2(n2977), 
	.C1(n2414), 
	.B2(FE_PHN748_n2415), 
	.B1(n2954), 
	.A(n2978));
   INV_X2 U2794 (.ZN(n2978), 
	.A(n2979));
   AOI221_X1 U2795 (.ZN(n2979), 
	.C2(n2872), 
	.C1(n2410), 
	.B2(n2871), 
	.B1(n2411), 
	.A(n2873));
   OAI221_X1 U2796 (.ZN(n2410), 
	.C2(n270), 
	.C1(n2981), 
	.B2(n16685), 
	.B1(n5625), 
	.A(FE_PHN935_n2982));
   AOI222_X1 U2797 (.ZN(n2982), 
	.C2(n2357), 
	.C1(n2912), 
	.B2(n2345), 
	.B1(n16645), 
	.A2(n2879), 
	.A1(hrdata_i[21]));
   NAND3_X1 U2799 (.ZN(n2411), 
	.A3(n2985), 
	.A2(n2984), 
	.A1(n2983));
   AOI221_X1 U2800 (.ZN(n2985), 
	.C2(n2878), 
	.C1(sub_2068_A_13_), 
	.B2(n2986), 
	.B1(n16787), 
	.A(n2987));
   OAI22_X1 U2801 (.ZN(n2987), 
	.B2(n2948), 
	.B1(n244), 
	.A2(n382), 
	.A1(n2918));
   INV_X1 U2802 (.ZN(n382), 
	.A(hrdata_i[13]));
   AOI22_X1 U2804 (.ZN(n2984), 
	.B2(n2988), 
	.B1(n16645), 
	.A2(n410), 
	.A1(n2895));
   OAI211_X1 U2805 (.ZN(n410), 
	.C2(n2989), 
	.C1(n1067), 
	.B(n4965), 
	.A(n5229));
   AOI211_X1 U2806 (.ZN(n2989), 
	.C2(n2990), 
	.C1(n2908), 
	.B(n1370), 
	.A(n2991));
   OAI21_X1 U2807 (.ZN(n2991), 
	.B2(n2992), 
	.B1(n2908), 
	.A(n2907));
   AOI22_X1 U2808 (.ZN(n2992), 
	.B2(n2995), 
	.B1(n2909), 
	.A2(n2994), 
	.A1(n2993));
   OAI21_X1 U2809 (.ZN(n2990), 
	.B2(n2910), 
	.B1(n2996), 
	.A(n2997));
   AOI22_X1 U2810 (.ZN(n2983), 
	.B2(n4751), 
	.B1(n2913), 
	.A2(n2353), 
	.A1(n2912));
   OAI221_X1 U2811 (.ZN(n2414), 
	.C2(FE_PHN765_n1144), 
	.C1(n2918), 
	.B2(n2374), 
	.B1(n2998), 
	.A(n2999));
   INV_X1 U2812 (.ZN(n2999), 
	.A(n3000));
   OAI21_X1 U2813 (.ZN(n3000), 
	.B2(n3002), 
	.B1(n3001), 
	.A(n3003));
   INV_X1 U2814 (.ZN(n1144), 
	.A(hrdata_i[29]));
   OAI221_X1 U2815 (.ZN(n2374), 
	.C2(n3004), 
	.C1(n16788), 
	.B2(FE_OFN527_n2336), 
	.B1(n2337), 
	.A(n3002));
   AOI22_X1 U2816 (.ZN(n3002), 
	.B2(n3006), 
	.B1(n2941), 
	.A2(n2940), 
	.A1(n3005));
   NAND2_X1 U2817 (.ZN(n2415), 
	.A2(n3008), 
	.A1(n3007));
   AOI221_X1 U2818 (.ZN(n3008), 
	.C2(n2330), 
	.C1(n2912), 
	.B2(n2326), 
	.B1(n16645), 
	.A(n3009));
   OAI22_X1 U2819 (.ZN(n3009), 
	.B2(n3011), 
	.B1(n5533), 
	.A2(n2948), 
	.A1(n3010));
   AOI222_X1 U2820 (.ZN(n3007), 
	.C2(n3012), 
	.C1(n16787), 
	.B2(n2879), 
	.B1(hrdata_i[5]), 
	.A2(n2878), 
	.A1(sub_2068_A_5_));
   INV_X1 U2822 (.ZN(n2974), 
	.A(n2308));
   NOR3_X1 U2823 (.ZN(n2308), 
	.A3(n1664), 
	.A2(n2501), 
	.A1(n3013));
   NAND2_X1 U2824 (.ZN(n2306), 
	.A2(n1664), 
	.A1(n3014));
   NAND4_X1 U2825 (.ZN(n1664), 
	.A4(n3018), 
	.A3(n3017), 
	.A2(n3016), 
	.A1(n3015));
   AOI222_X1 U2826 (.ZN(n3018), 
	.C2(vis_r9_o[13]), 
	.C1(n16979), 
	.B2(n2970), 
	.B1(n16976), 
	.A2(vis_r8_o[13]), 
	.A1(n16958));
   AOI222_X1 U2829 (.ZN(n3017), 
	.C2(vis_r11_o[13]), 
	.C1(n16987), 
	.B2(n3022), 
	.B1(n16970), 
	.A2(vis_r10_o[13]), 
	.A1(n16961));
   AOI222_X1 U2831 (.ZN(n3016), 
	.C2(vis_r12_o[13]), 
	.C1(FE_OFN109_n16964), 
	.B2(vis_r14_o[13]), 
	.B1(n16984), 
	.A2(vis_msp_o[11]), 
	.A1(n16974));
   AOI22_X1 U2834 (.ZN(n3015), 
	.B2(n16956), 
	.B1(n3028), 
	.A2(vis_psp_o[11]), 
	.A1(n16969));
   OAI22_X1 U2835 (.ZN(n3014), 
	.B2(n3013), 
	.B1(n2131), 
	.A2(n5808), 
	.A1(n16992));
   INV_X1 U2836 (.ZN(n3013), 
	.A(n5808));
   XOR2_X1 U2837 (.Z(n5808), 
	.B(n3029), 
	.A(n2169));
   AOI221_X1 U2838 (.ZN(n3029), 
	.C2(FE_OFN602_n16656), 
	.C1(n2198), 
	.B2(n2259), 
	.B1(n16989), 
	.A(n2732));
   OAI22_X1 U2839 (.ZN(U367_Z_0), 
	.B2(n17005), 
	.B1(n3030), 
	.A2(n17001), 
	.A1(FE_PHN2550_n5131));
   OAI22_X1 U2840 (.ZN(U366_Z_0), 
	.B2(n17000), 
	.B1(n3030), 
	.A2(n16996), 
	.A1(FE_PHN2789_n5130));
   OAI22_X1 U2841 (.ZN(U365_Z_0), 
	.B2(n17042), 
	.B1(n3030), 
	.A2(n17038), 
	.A1(FE_PHN2645_n5301));
   OAI22_X1 U2842 (.ZN(U364_Z_0), 
	.B2(n17037), 
	.B1(n3030), 
	.A2(FE_OFN652_n17033), 
	.A1(FE_PHN2513_n5280));
   OAI22_X1 U2843 (.ZN(U363_Z_0), 
	.B2(n17031), 
	.B1(n3030), 
	.A2(n17028), 
	.A1(n5129));
   OAI22_X1 U2844 (.ZN(U362_Z_0), 
	.B2(FE_OFN651_n17027), 
	.B1(n3030), 
	.A2(n17023), 
	.A1(FE_PHN2670_n5192));
   OAI22_X1 U2845 (.ZN(U361_Z_0), 
	.B2(n17022), 
	.B1(n3030), 
	.A2(n17018), 
	.A1(FE_PHN2579_n5128));
   OAI22_X1 U2846 (.ZN(U360_Z_0), 
	.B2(FE_OFN648_n17017), 
	.B1(n3030), 
	.A2(n17013), 
	.A1(FE_PHN2519_n5221));
   OAI22_X1 U2847 (.ZN(U359_Z_0), 
	.B2(n17046), 
	.B1(n3030), 
	.A2(n17043), 
	.A1(n5328));
   OAI22_X1 U2848 (.ZN(U358_Z_0), 
	.B2(n17052), 
	.B1(n3030), 
	.A2(n17048), 
	.A1(FE_PHN2595_n5357));
   OAI22_X1 U2849 (.ZN(U357_Z_0), 
	.B2(FE_OFN661_n17057), 
	.B1(n3030), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2602_n5386));
   OAI22_X1 U2850 (.ZN(U356_Z_0), 
	.B2(n17062), 
	.B1(n3030), 
	.A2(FE_OFN663_n17058), 
	.A1(FE_PHN2624_n5415));
   OAI22_X1 U2851 (.ZN(U355_Z_0), 
	.B2(n17067), 
	.B1(n3030), 
	.A2(n17063), 
	.A1(FE_PHN2668_n5444));
   OAI22_X1 U2852 (.ZN(U354_Z_0), 
	.B2(n17071), 
	.B1(n3030), 
	.A2(n17068), 
	.A1(FE_PHN2671_n5473));
   OAI22_X1 U2853 (.ZN(U353_Z_0), 
	.B2(n17077), 
	.B1(n3030), 
	.A2(FE_OFN665_n17074), 
	.A1(n5127));
   OAI22_X1 U2854 (.ZN(U352_Z_0), 
	.B2(n17082), 
	.B1(n3030), 
	.A2(n17078), 
	.A1(FE_PHN2503_n5497));
   AOI221_X1 U2856 (.ZN(n3032), 
	.C2(FE_OFN208_n2015), 
	.C1(n16653), 
	.B2(n2247), 
	.B1(n17008), 
	.A(n2055));
   OAI221_X1 U2857 (.ZN(n3031), 
	.C2(n1665), 
	.C1(n16994), 
	.B2(n5807), 
	.B1(n3033), 
	.A(n3034));
   NAND3_X1 U2858 (.ZN(n3034), 
	.A3(n5807), 
	.A2(n1665), 
	.A1(n2131));
   AOI221_X1 U2860 (.ZN(n3035), 
	.C2(n2231), 
	.C1(n2198), 
	.B2(n2247), 
	.B1(n16989), 
	.A(n2732));
   NOR2_X1 U2861 (.ZN(n3033), 
	.A2(n16992), 
	.A1(n1694));
   INV_X1 U2862 (.ZN(n1694), 
	.A(n1665));
   NAND4_X1 U2863 (.ZN(n1665), 
	.A4(n3039), 
	.A3(n3038), 
	.A2(n3037), 
	.A1(n3036));
   AOI222_X1 U2864 (.ZN(n3039), 
	.C2(vis_psp_o[10]), 
	.C1(n16968), 
	.B2(n3041), 
	.B1(n16970), 
	.A2(vis_msp_o[10]), 
	.A1(n16974));
   AOI222_X1 U2866 (.ZN(n3038), 
	.C2(vis_r11_o[12]), 
	.C1(n16987), 
	.B2(vis_r12_o[12]), 
	.B1(n16966), 
	.A2(vis_r14_o[12]), 
	.A1(n16983));
   AOI222_X1 U2869 (.ZN(n3037), 
	.C2(vis_r8_o[12]), 
	.C1(n16959), 
	.B2(vis_r10_o[12]), 
	.B1(n16962), 
	.A2(vis_r9_o[12]), 
	.A1(n16980));
   AOI22_X1 U2871 (.ZN(n3036), 
	.B2(n3049), 
	.B1(n16955), 
	.A2(n3028), 
	.A1(n16976));
   INV_X1 U2873 (.ZN(n136), 
	.A(n3050));
   OAI221_X1 U2874 (.ZN(n3050), 
	.C2(n2869), 
	.C1(n2596), 
	.B2(n3051), 
	.B1(n2757), 
	.A(n3052));
   AOI221_X1 U2875 (.ZN(n3052), 
	.C2(n2954), 
	.C1(n2068), 
	.B2(n2075), 
	.B1(n2871), 
	.A(n2873));
   NAND3_X1 U2876 (.ZN(n2068), 
	.A3(n3055), 
	.A2(n3054), 
	.A1(n3053));
   AOI221_X1 U2877 (.ZN(n3055), 
	.C2(n2878), 
	.C1(sub_2068_A_4_), 
	.B2(n3056), 
	.B1(n16787), 
	.A(n3057));
   OAI22_X1 U2878 (.ZN(n3057), 
	.B2(n2948), 
	.B1(n4800), 
	.A2(FE_PHN870_n420), 
	.A1(n2918));
   INV_X1 U2879 (.ZN(n420), 
	.A(hrdata_i[4]));
   AOI22_X1 U2881 (.ZN(n3054), 
	.B2(n2333), 
	.B1(n16645), 
	.A2(n3059), 
	.A1(n3058));
   AOI22_X1 U2883 (.ZN(n3053), 
	.B2(n3060), 
	.B1(n2913), 
	.A2(n2339), 
	.A1(n2912));
   NAND3_X1 U2884 (.ZN(n2075), 
	.A3(FE_PHN1025_n3063), 
	.A2(n3062), 
	.A1(n3061));
   AOI221_X1 U2885 (.ZN(n3063), 
	.C2(n2878), 
	.C1(sub_2068_A_12_), 
	.B2(n2879), 
	.B1(hrdata_i[12]), 
	.A(n3064));
   OAI22_X1 U2886 (.ZN(n3064), 
	.B2(n2948), 
	.B1(n4795), 
	.A2(n16685), 
	.A1(FE_PHN2428_n5507));
   AOI22_X1 U2887 (.ZN(n3062), 
	.B2(n2387), 
	.B1(n16645), 
	.A2(n2895), 
	.A1(n417));
   INV_X1 U2888 (.ZN(n417), 
	.A(n412));
   OAI21_X1 U2889 (.ZN(n412), 
	.B2(n3066), 
	.B1(n3065), 
	.A(n4965));
   AOI211_X1 U2890 (.ZN(n3065), 
	.C2(n2903), 
	.C1(n1370), 
	.B(n3067), 
	.A(n1067));
   AOI211_X1 U2891 (.ZN(n3067), 
	.C2(n2911), 
	.C1(n3068), 
	.B(n1370), 
	.A(n3069));
   OAI21_X1 U2892 (.ZN(n3069), 
	.B2(n2911), 
	.B1(n3070), 
	.A(n2907));
   AOI221_X1 U2893 (.ZN(n3070), 
	.C2(n3074), 
	.C1(n3073), 
	.B2(n3072), 
	.B1(n3071), 
	.A(n3075));
   NOR3_X1 U2894 (.ZN(n3075), 
	.A3(n3077), 
	.A2(n3073), 
	.A1(n3076));
   OAI21_X1 U2895 (.ZN(n3074), 
	.B2(n3079), 
	.B1(n3078), 
	.A(n3080));
   INV_X1 U2896 (.ZN(n3071), 
	.A(n2997));
   OAI22_X1 U2897 (.ZN(n3068), 
	.B2(n2909), 
	.B1(n3082), 
	.A2(n3081), 
	.A1(n2993));
   INV_X1 U2898 (.ZN(n3082), 
	.A(n3083));
   OAI21_X1 U2899 (.ZN(n3083), 
	.B2(n3084), 
	.B1(n2994), 
	.A(n3085));
   AOI22_X1 U2900 (.ZN(n3081), 
	.B2(n3088), 
	.B1(n2995), 
	.A2(n3087), 
	.A1(n3086));
   AOI22_X1 U2901 (.ZN(n3061), 
	.B2(n3089), 
	.B1(n2913), 
	.A2(n2385), 
	.A1(n2912));
   AOI221_X1 U2902 (.ZN(n2596), 
	.C2(n2922), 
	.C1(n2364), 
	.B2(n2895), 
	.B1(n209), 
	.A(n3090));
   OAI21_X1 U2903 (.ZN(n3090), 
	.B2(n2918), 
	.B1(FE_PHN806_n1143), 
	.A(n3003));
   INV_X1 U2904 (.ZN(n1143), 
	.A(hrdata_i[28]));
   OAI22_X1 U2905 (.ZN(n2364), 
	.B2(n3093), 
	.B1(n2940), 
	.A2(n3092), 
	.A1(n3091));
   AOI22_X1 U2906 (.ZN(n3093), 
	.B2(n3095), 
	.B1(n2337), 
	.A2(n3094), 
	.A1(n16788));
   INV_X1 U2907 (.ZN(n2757), 
	.A(n2066));
   OAI221_X1 U2908 (.ZN(n2066), 
	.C2(n272), 
	.C1(n2981), 
	.B2(n16685), 
	.B1(FE_PHN2378_n5618), 
	.A(FE_PHN743_n3096));
   AOI222_X1 U2909 (.ZN(n3096), 
	.C2(FE_OFN530_n2350), 
	.C1(n2912), 
	.B2(n2355), 
	.B1(n16645), 
	.A2(n2879), 
	.A1(hrdata_i[20]));
   OAI22_X1 U2911 (.ZN(U349_Z_0), 
	.B2(n17005), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17001), 
	.A1(FE_PHN2452_n5569));
   OAI22_X1 U2912 (.ZN(U348_Z_0), 
	.B2(n17000), 
	.B1(FE_PSN5238_n3097), 
	.A2(n16996), 
	.A1(FE_PHN2784_n5568));
   OAI22_X1 U2913 (.ZN(U347_Z_0), 
	.B2(n17042), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17038), 
	.A1(FE_PHN2660_n5567));
   OAI22_X1 U2914 (.ZN(U346_Z_0), 
	.B2(n17037), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17033), 
	.A1(FE_PHN2531_n5566));
   OAI22_X1 U2915 (.ZN(U345_Z_0), 
	.B2(n17031), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17028), 
	.A1(FE_PHN4750_n5565));
   OAI22_X1 U2916 (.ZN(U344_Z_0), 
	.B2(FE_OFN651_n17027), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17023), 
	.A1(FE_PHN2709_n5564));
   OAI22_X1 U2917 (.ZN(U343_Z_0), 
	.B2(n17022), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17018), 
	.A1(FE_PHN2523_n5563));
   OAI22_X1 U2918 (.ZN(U342_Z_0), 
	.B2(FE_OFN648_n17017), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17013), 
	.A1(FE_PHN2552_n5562));
   OAI22_X1 U2919 (.ZN(U341_Z_0), 
	.B2(n17046), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17043), 
	.A1(FE_PHN4732_n5561));
   OAI22_X1 U2920 (.ZN(U340_Z_0), 
	.B2(n17052), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17048), 
	.A1(FE_PHN2560_n5560));
   OAI22_X1 U2921 (.ZN(U339_Z_0), 
	.B2(n17057), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17053), 
	.A1(FE_PHN2465_n5559));
   OAI22_X1 U2922 (.ZN(U338_Z_0), 
	.B2(n17062), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17058), 
	.A1(FE_PHN2644_n5558));
   OAI22_X1 U2923 (.ZN(U337_Z_0), 
	.B2(n17067), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17063), 
	.A1(FE_PHN2777_n5557));
   OAI22_X1 U2924 (.ZN(U336_Z_0), 
	.B2(n17071), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17068), 
	.A1(FE_PHN3568_n5556));
   OAI22_X1 U2925 (.ZN(U335_Z_0), 
	.B2(n17077), 
	.B1(FE_PSN5238_n3097), 
	.A2(FE_OFN665_n17074), 
	.A1(FE_PHN4734_n5555));
   OAI22_X1 U2926 (.ZN(U334_Z_0), 
	.B2(n17082), 
	.B1(FE_PSN5238_n3097), 
	.A2(n17078), 
	.A1(FE_PHN2590_n5554));
   INV_X2 U2928 (.ZN(n3098), 
	.A(n3099));
   AOI221_X1 U2929 (.ZN(n3099), 
	.C2(n2246), 
	.C1(n17008), 
	.B2(FE_OFN208_n2015), 
	.B1(n16719), 
	.A(n126));
   OAI221_X1 U2930 (.ZN(n126), 
	.C2(n2419), 
	.C1(n2869), 
	.B2(n2418), 
	.B1(n3051), 
	.A(n3100));
   AOI221_X1 U2931 (.ZN(n3100), 
	.C2(n2954), 
	.C1(n2422), 
	.B2(n2871), 
	.B1(FE_PHN728_n2421), 
	.A(n2873));
   NAND3_X1 U2932 (.ZN(n2422), 
	.A3(n3103), 
	.A2(n3102), 
	.A1(n3101));
   AOI221_X1 U2933 (.ZN(n3103), 
	.C2(n2878), 
	.C1(sub_2068_A_3_), 
	.B2(n3104), 
	.B1(n16787), 
	.A(n3105));
   OAI22_X1 U2934 (.ZN(n3105), 
	.B2(n2948), 
	.B1(n5536), 
	.A2(FE_PHN875_n423), 
	.A1(n2918));
   INV_X1 U2935 (.ZN(n423), 
	.A(hrdata_i[3]));
   AOI21_X1 U2937 (.ZN(n3102), 
	.B2(n2334), 
	.B1(n16645), 
	.A(n3106));
   AOI22_X1 U2938 (.ZN(n3101), 
	.B2(n3107), 
	.B1(n2913), 
	.A2(n2338), 
	.A1(n2912));
   NAND3_X1 U2939 (.ZN(n2421), 
	.A3(n3110), 
	.A2(n3109), 
	.A1(n3108));
   AOI222_X1 U2940 (.ZN(n3110), 
	.C2(n3111), 
	.C1(n16787), 
	.B2(n2879), 
	.B1(hrdata_i[11]), 
	.A2(n2878), 
	.A1(sub_2068_A_11_));
   AOI22_X1 U2942 (.ZN(n3109), 
	.B2(n2384), 
	.B1(n2912), 
	.A2(n2386), 
	.A1(n16645));
   INV_X1 U2943 (.ZN(n3108), 
	.A(n3112));
   OAI22_X1 U2944 (.ZN(n3112), 
	.B2(n5570), 
	.B1(n2948), 
	.A2(n5572), 
	.A1(n3011));
   INV_X1 U2945 (.ZN(n2419), 
	.A(n2623));
   OAI211_X1 U2946 (.ZN(n2623), 
	.C2(n2368), 
	.C1(n3113), 
	.B(n3114), 
	.A(n3003));
   INV_X1 U2947 (.ZN(n3114), 
	.A(n3115));
   OAI22_X1 U2948 (.ZN(n3115), 
	.B2(n2918), 
	.B1(FE_PHN755_n1142), 
	.A2(n3001), 
	.A1(n3116));
   INV_X1 U2949 (.ZN(n1142), 
	.A(hrdata_i[27]));
   OAI21_X1 U2950 (.ZN(n2368), 
	.B2(n3117), 
	.B1(n16788), 
	.A(n3116));
   OAI221_X1 U2951 (.ZN(n3116), 
	.C2(n16951), 
	.C1(n3120), 
	.B2(n3119), 
	.B1(n3118), 
	.A(n3122));
   AOI21_X1 U2952 (.ZN(n3113), 
	.B2(n2369), 
	.B1(n2922), 
	.A(n16645));
   INV_X1 U2953 (.ZN(n2418), 
	.A(FE_PHN859_n2624));
   OAI211_X1 U2954 (.ZN(n2624), 
	.C2(n2875), 
	.C1(n3123), 
	.B(n3125), 
	.A(n3124));
   AOI222_X1 U2955 (.ZN(n3125), 
	.C2(n3126), 
	.C1(n16787), 
	.B2(n2879), 
	.B1(hrdata_i[19]), 
	.A2(n2878), 
	.A1(sub_2068_A_19_));
   AOI21_X1 U2957 (.ZN(n3124), 
	.B2(n2354), 
	.B1(n16645), 
	.A(n2897));
   INV_X1 U2958 (.ZN(n3123), 
	.A(n2356));
   AOI221_X1 U2959 (.ZN(n2310), 
	.C2(n16992), 
	.C1(n3127), 
	.B2(n2131), 
	.B1(n5820), 
	.A(n1695));
   INV_X1 U2960 (.ZN(n1695), 
	.A(n3128));
   NOR3_X1 U2961 (.ZN(n2309), 
	.A3(n3128), 
	.A2(n2501), 
	.A1(n3127));
   NAND4_X1 U2962 (.ZN(n3128), 
	.A4(n3132), 
	.A3(n3131), 
	.A2(n3130), 
	.A1(n3129));
   AOI222_X1 U2963 (.ZN(n3132), 
	.C2(vis_psp_o[9]), 
	.C1(n16968), 
	.B2(n3134), 
	.B1(n16970), 
	.A2(vis_msp_o[9]), 
	.A1(n16974));
   AOI222_X1 U2965 (.ZN(n3131), 
	.C2(vis_r11_o[11]), 
	.C1(n16987), 
	.B2(vis_r12_o[11]), 
	.B1(n16966), 
	.A2(vis_r14_o[11]), 
	.A1(n16983));
   AOI222_X1 U2968 (.ZN(n3130), 
	.C2(vis_r8_o[11]), 
	.C1(FE_PSN5236_n16960), 
	.B2(vis_r10_o[11]), 
	.B1(n16963), 
	.A2(vis_r9_o[11]), 
	.A1(n16980));
   AOI22_X1 U2970 (.ZN(n3129), 
	.B2(n3142), 
	.B1(n16956), 
	.A2(n3049), 
	.A1(n16976));
   INV_X1 U2972 (.ZN(n3127), 
	.A(n5820));
   XOR2_X1 U2973 (.Z(n5820), 
	.B(n3143), 
	.A(n2169));
   AOI221_X1 U2974 (.ZN(n3143), 
	.C2(n16817), 
	.C1(n2198), 
	.B2(n2246), 
	.B1(n16989), 
	.A(n2732));
   OAI22_X1 U2975 (.ZN(U333_Z_0), 
	.B2(n17005), 
	.B1(n3144), 
	.A2(n17001), 
	.A1(FE_PHN3580_n5148));
   OAI22_X1 U2976 (.ZN(U332_Z_0), 
	.B2(n17000), 
	.B1(n3144), 
	.A2(n16996), 
	.A1(FE_PHN3627_n5147));
   OAI22_X1 U2977 (.ZN(U331_Z_0), 
	.B2(n17042), 
	.B1(n3144), 
	.A2(n17038), 
	.A1(FE_PHN3681_n5302));
   OAI22_X1 U2978 (.ZN(U330_Z_0), 
	.B2(n17037), 
	.B1(n3144), 
	.A2(n17033), 
	.A1(FE_PHN3555_n5281));
   OAI22_X1 U2979 (.ZN(U329_Z_0), 
	.B2(n17031), 
	.B1(n3144), 
	.A2(n17028), 
	.A1(n5146));
   OAI22_X1 U2980 (.ZN(U328_Z_0), 
	.B2(FE_OFN651_n17027), 
	.B1(n3144), 
	.A2(n17023), 
	.A1(FE_PHN3726_n5193));
   OAI22_X1 U2981 (.ZN(U327_Z_0), 
	.B2(n17022), 
	.B1(n3144), 
	.A2(n17018), 
	.A1(FE_PHN3596_n5145));
   OAI22_X1 U2982 (.ZN(U326_Z_0), 
	.B2(n17017), 
	.B1(n3144), 
	.A2(n17013), 
	.A1(FE_PHN3570_n5222));
   OAI22_X1 U2983 (.ZN(U325_Z_0), 
	.B2(n17046), 
	.B1(n3144), 
	.A2(n17043), 
	.A1(n5329));
   OAI22_X1 U2984 (.ZN(U324_Z_0), 
	.B2(n17052), 
	.B1(n3144), 
	.A2(n17048), 
	.A1(n5358));
   OAI22_X1 U2985 (.ZN(U323_Z_0), 
	.B2(n17057), 
	.B1(n3144), 
	.A2(n17053), 
	.A1(n5387));
   OAI22_X1 U2986 (.ZN(U322_Z_0), 
	.B2(n17062), 
	.B1(n3144), 
	.A2(n17058), 
	.A1(FE_PHN3622_n5416));
   OAI22_X1 U2987 (.ZN(U321_Z_0), 
	.B2(n17067), 
	.B1(n3144), 
	.A2(n17063), 
	.A1(n5445));
   OAI22_X1 U2988 (.ZN(U320_Z_0), 
	.B2(n17071), 
	.B1(n3144), 
	.A2(n17068), 
	.A1(n5474));
   OAI22_X1 U2989 (.ZN(U319_Z_0), 
	.B2(n17077), 
	.B1(n3144), 
	.A2(n17074), 
	.A1(n5144));
   OAI22_X2 U2990 (.ZN(U318_Z_0), 
	.B2(n17082), 
	.B1(n3144), 
	.A2(n17078), 
	.A1(n5498));
   AOI221_X1 U2992 (.ZN(n2114), 
	.C2(n17008), 
	.C1(n3145), 
	.B2(n16723), 
	.B1(n2495), 
	.A(n3146));
   INV_X1 U2993 (.ZN(n3146), 
	.A(n3147));
   AOI211_X1 U2994 (.ZN(n3147), 
	.C2(n3148), 
	.C1(n5804), 
	.B(n3149), 
	.A(n2055));
   NOR3_X1 U2995 (.ZN(n3149), 
	.A3(n1696), 
	.A2(n16992), 
	.A1(n5804));
   OAI22_X1 U2996 (.ZN(n3148), 
	.B2(n1667), 
	.B1(n2501), 
	.A2(n1696), 
	.A1(n2131));
   INV_X1 U2997 (.ZN(n1696), 
	.A(n1667));
   NAND4_X1 U2998 (.ZN(n1667), 
	.A4(n3153), 
	.A3(n3152), 
	.A2(n3151), 
	.A1(n3150));
   AOI222_X1 U2999 (.ZN(n3153), 
	.C2(vis_psp_o[8]), 
	.C1(n16969), 
	.B2(n3155), 
	.B1(n16970), 
	.A2(vis_msp_o[8]), 
	.A1(n16974));
   AOI222_X1 U3001 (.ZN(n3152), 
	.C2(vis_r11_o[10]), 
	.C1(n16987), 
	.B2(vis_r12_o[10]), 
	.B1(n16966), 
	.A2(vis_r14_o[10]), 
	.A1(n16983));
   AOI222_X1 U3004 (.ZN(n3151), 
	.C2(vis_r8_o[10]), 
	.C1(FE_PSN5236_n16960), 
	.B2(vis_r10_o[10]), 
	.B1(n16963), 
	.A2(vis_r9_o[10]), 
	.A1(n16980));
   AOI22_X1 U3006 (.ZN(n3150), 
	.B2(n869), 
	.B1(n16956), 
	.A2(n3142), 
	.A1(n16976));
   XOR2_X1 U3008 (.Z(n5804), 
	.B(n3163), 
	.A(n2169));
   AOI222_X1 U3009 (.ZN(n3163), 
	.C2(n2731), 
	.C1(n3164), 
	.B2(n16657), 
	.B1(n2198), 
	.A2(n3145), 
	.A1(n16988));
   AOI221_X1 U3010 (.ZN(n140), 
	.C2(n2871), 
	.C1(FE_PHN679_n2465), 
	.B2(n2954), 
	.B1(n2464), 
	.A(n3165));
   INV_X2 U3011 (.ZN(n3165), 
	.A(n3166));
   AOI221_X1 U3012 (.ZN(n3166), 
	.C2(n2872), 
	.C1(n2469), 
	.B2(n2977), 
	.B1(n2468), 
	.A(n2873));
   OAI22_X1 U3013 (.ZN(U317_Z_0), 
	.B2(n3169), 
	.B1(n3168), 
	.A2(n3167), 
	.A1(n5546));
   AOI22_X1 U3014 (.ZN(n3168), 
	.B2(n1058), 
	.B1(n3170), 
	.A2(n1640), 
	.A1(n1040));
   INV_X1 U3015 (.ZN(n3167), 
	.A(n3169));
   OAI211_X1 U3016 (.ZN(n3169), 
	.C2(n1880), 
	.C1(n1173), 
	.B(n195), 
	.A(n17122));
   INV_X1 U3017 (.ZN(n1880), 
	.A(FE_OFN461_n890));
   OAI22_X1 U3018 (.ZN(U315_Z_0), 
	.B2(n17005), 
	.B1(n3171), 
	.A2(n17001), 
	.A1(FE_PHN3554_n5060));
   OAI22_X1 U3019 (.ZN(U314_Z_0), 
	.B2(n17000), 
	.B1(n3171), 
	.A2(n16996), 
	.A1(FE_PHN3589_n5059));
   OAI22_X1 U3020 (.ZN(U313_Z_0), 
	.B2(n17042), 
	.B1(n3171), 
	.A2(n17038), 
	.A1(FE_PHN3560_n5303));
   OAI22_X1 U3021 (.ZN(U312_Z_0), 
	.B2(n17037), 
	.B1(n3171), 
	.A2(n17033), 
	.A1(FE_PHN3569_n5282));
   OAI22_X1 U3022 (.ZN(U311_Z_0), 
	.B2(n17031), 
	.B1(n3171), 
	.A2(n17028), 
	.A1(FE_PHN3623_n5058));
   OAI22_X1 U3023 (.ZN(U310_Z_0), 
	.B2(n17027), 
	.B1(n3171), 
	.A2(n17023), 
	.A1(FE_PHN3630_n5194));
   OAI22_X1 U3024 (.ZN(U309_Z_0), 
	.B2(n17022), 
	.B1(n3171), 
	.A2(n17018), 
	.A1(n5057));
   OAI22_X1 U3025 (.ZN(U308_Z_0), 
	.B2(n17017), 
	.B1(n3171), 
	.A2(n17013), 
	.A1(FE_PHN5065_n5223));
   OAI22_X1 U3026 (.ZN(U307_Z_0), 
	.B2(n17046), 
	.B1(n3171), 
	.A2(n17043), 
	.A1(FE_PHN3594_n5330));
   OAI22_X1 U3027 (.ZN(U306_Z_0), 
	.B2(n17052), 
	.B1(n3171), 
	.A2(n17048), 
	.A1(FE_PHN3587_n5359));
   OAI22_X1 U3028 (.ZN(U305_Z_0), 
	.B2(n17057), 
	.B1(n3171), 
	.A2(n17053), 
	.A1(n5388));
   OAI22_X1 U3029 (.ZN(U304_Z_0), 
	.B2(n17062), 
	.B1(n3171), 
	.A2(n17058), 
	.A1(FE_PHN3550_n5417));
   OAI22_X1 U3030 (.ZN(U303_Z_0), 
	.B2(n17067), 
	.B1(n3171), 
	.A2(n17063), 
	.A1(FE_PHN3626_n5446));
   OAI22_X1 U3031 (.ZN(U302_Z_0), 
	.B2(n17071), 
	.B1(n3171), 
	.A2(n17068), 
	.A1(FE_PHN3634_n5475));
   OAI22_X1 U3032 (.ZN(U301_Z_0), 
	.B2(n17077), 
	.B1(n3171), 
	.A2(n17074), 
	.A1(FE_PHN4756_n5056));
   OAI22_X1 U3033 (.ZN(U300_Z_0), 
	.B2(n17082), 
	.B1(n3171), 
	.A2(n17078), 
	.A1(FE_PHN3621_n5499));
   AND4_X1 U3035 (.ZN(n2115), 
	.A4(n3175), 
	.A3(n3174), 
	.A2(n3173), 
	.A1(n3172));
   AOI222_X1 U3036 (.ZN(n3175), 
	.C2(n3177), 
	.C1(n17008), 
	.B2(vis_control_o), 
	.B1(n2055), 
	.A2(FE_OFN2_n2015), 
	.A1(n16729));
   AOI22_X1 U3038 (.ZN(n3174), 
	.B2(vis_ipsr_o[2]), 
	.B1(n2227), 
	.A2(n3178), 
	.A1(n5806));
   NOR3_X1 U3039 (.ZN(n2227), 
	.A3(n2168), 
	.A2(n5120), 
	.A1(FE_OFN15_n16671));
   OAI22_X2 U3040 (.ZN(n3178), 
	.B2(n1640), 
	.B1(n2501), 
	.A2(n1676), 
	.A1(n2131));
   OR4_X1 U3041 (.ZN(n3173), 
	.A4(n4950), 
	.A3(n16854), 
	.A2(n5546), 
	.A1(n1308));
   NAND2_X1 U3042 (.ZN(n1308), 
	.A2(n16728), 
	.A1(n17096));
   OR3_X1 U3043 (.ZN(n3172), 
	.A3(n5806), 
	.A2(n16992), 
	.A1(n1676));
   XNOR2_X1 U3044 (.ZN(n5806), 
	.B(n3179), 
	.A(n16990));
   OAI221_X1 U3045 (.ZN(n3179), 
	.C2(n3181), 
	.C1(n3180), 
	.B2(n2554), 
	.B1(n5120), 
	.A(n3182));
   AOI22_X1 U3046 (.ZN(n3182), 
	.B2(n2173), 
	.B1(n16656), 
	.A2(n2198), 
	.A1(n461));
   NAND2_X1 U3047 (.ZN(n2173), 
	.A2(n3183), 
	.A1(n2201));
   NAND4_X1 U3048 (.ZN(n3183), 
	.A4(FE_OFN10_n1697), 
	.A3(n16843), 
	.A2(n2661), 
	.A1(n1097));
   INV_X1 U3049 (.ZN(n2201), 
	.A(n3184));
   OAI21_X1 U3050 (.ZN(n3184), 
	.B2(n3185), 
	.B1(n4950), 
	.A(n3186));
   AOI221_X1 U3051 (.ZN(n3185), 
	.C2(n16871), 
	.C1(n3188), 
	.B2(n3187), 
	.B1(n16862), 
	.A(n3189));
   OAI22_X1 U3052 (.ZN(n3189), 
	.B2(n655), 
	.B1(n919), 
	.A2(n1517), 
	.A1(n1104));
   NAND2_X1 U3053 (.ZN(n655), 
	.A2(n16838), 
	.A1(n17097));
   OAI21_X1 U3054 (.ZN(n3188), 
	.B2(n1211), 
	.B1(n16837), 
	.A(n919));
   NAND2_X1 U3055 (.ZN(n919), 
	.A2(FE_OFN81_n16856), 
	.A1(n16828));
   OAI22_X1 U3056 (.ZN(n3187), 
	.B2(n648), 
	.B1(FE_OFN17_n16805), 
	.A2(n1104), 
	.A1(n16851));
   INV_X1 U3057 (.ZN(n3181), 
	.A(n3177));
   INV_X1 U3058 (.ZN(n2554), 
	.A(n2577));
   OAI21_X1 U3059 (.ZN(n2577), 
	.B2(n3190), 
	.B1(n4950), 
	.A(n2200));
   AOI221_X1 U3060 (.ZN(n3190), 
	.C2(FE_OFN84_n16839), 
	.C1(n507), 
	.B2(FE_OFN633_n16868), 
	.B1(n3191), 
	.A(n3192));
   OAI22_X1 U3061 (.ZN(n3192), 
	.B2(n1211), 
	.B1(FE_OFN107_n585), 
	.A2(n673), 
	.A1(FE_OFN73_n16806));
   NAND2_X1 U3062 (.ZN(n507), 
	.A2(n994), 
	.A1(n499));
   AOI21_X1 U3063 (.ZN(n3191), 
	.B2(n3193), 
	.B1(n1603), 
	.A(FE_OFN70_n16867));
   NAND2_X1 U3064 (.ZN(n3193), 
	.A2(FE_OFN632_n16859), 
	.A1(n1564));
   INV_X4 U3065 (.ZN(n1676), 
	.A(n1640));
   NAND4_X2 U3066 (.ZN(n1640), 
	.A4(n3197), 
	.A3(n3196), 
	.A2(n3195), 
	.A1(n3194));
   AOI222_X1 U3067 (.ZN(n3197), 
	.C2(vis_psp_o[0]), 
	.C1(n16969), 
	.B2(n3199), 
	.B1(n16970), 
	.A2(vis_msp_o[0]), 
	.A1(n16975));
   AOI222_X1 U3068 (.ZN(n3196), 
	.C2(vis_r11_o[2]), 
	.C1(n16987), 
	.B2(vis_r12_o[2]), 
	.B1(n16966), 
	.A2(vis_r14_o[2]), 
	.A1(n16984));
   AOI222_X1 U3069 (.ZN(n3195), 
	.C2(vis_r8_o[2]), 
	.C1(n16960), 
	.B2(vis_r10_o[2]), 
	.B1(n16963), 
	.A2(vis_r9_o[2]), 
	.A1(n16979));
   AOI22_X1 U3070 (.ZN(n3194), 
	.B2(n2635), 
	.B1(n16955), 
	.A2(n2620), 
	.A1(n16976));
   AOI221_X1 U3072 (.ZN(n171), 
	.C2(FE_PHN679_n2465), 
	.C1(n2002), 
	.B2(n2468), 
	.B1(n2008), 
	.A(n3207));
   INV_X2 U3073 (.ZN(n3207), 
	.A(n3208));
   AOI221_X1 U3074 (.ZN(n3208), 
	.C2(n2004), 
	.C1(n2464), 
	.B2(n2011), 
	.B1(n2469), 
	.A(n2012));
   AND4_X1 U3075 (.ZN(n2012), 
	.A4(n3212), 
	.A3(n3211), 
	.A2(n3210), 
	.A1(n3209));
   AOI222_X1 U3076 (.ZN(n3212), 
	.C2(1'b1), 
	.C1(n3215), 
	.B2(n2341), 
	.B1(n3214), 
	.A2(n3213), 
	.A1(n2360));
   INV_X1 U3077 (.ZN(n2360), 
	.A(n3217));
   AOI211_X1 U3079 (.ZN(n3218), 
	.C2(n606), 
	.C1(n3219), 
	.B(n3220), 
	.A(n1712));
   AOI211_X1 U3080 (.ZN(n3220), 
	.C2(n3221), 
	.C1(n16843), 
	.B(n3223), 
	.A(n3222));
   NAND2_X1 U3081 (.ZN(n3219), 
	.A2(FE_OFN81_n16856), 
	.A1(n16838));
   NAND3_X1 U3082 (.ZN(n2464), 
	.A3(n3226), 
	.A2(n3225), 
	.A1(n3224));
   AOI221_X1 U3083 (.ZN(n3226), 
	.C2(n2878), 
	.C1(sub_2068_A_2_), 
	.B2(n3227), 
	.B1(n16787), 
	.A(n3228));
   OAI22_X1 U3084 (.ZN(n3228), 
	.B2(n2948), 
	.B1(n4801), 
	.A2(FE_PHN844_n425), 
	.A1(n2918));
   INV_X1 U3085 (.ZN(n425), 
	.A(hrdata_i[2]));
   AOI221_X1 U3087 (.ZN(n3225), 
	.C2(n3229), 
	.C1(n3058), 
	.B2(n2325), 
	.B1(n2912), 
	.A(n3230));
   OAI221_X1 U3089 (.ZN(n2325), 
	.C2(n16951), 
	.C1(n3233), 
	.B2(n16948), 
	.B1(n3231), 
	.A(n3234));
   AOI22_X1 U3090 (.ZN(n3234), 
	.B2(n3237), 
	.B1(n16942), 
	.A2(n2209), 
	.A1(n16945));
   AOI22_X1 U3091 (.ZN(n3224), 
	.B2(n3238), 
	.B1(n2913), 
	.A2(n2332), 
	.A1(n16645));
   OAI221_X1 U3092 (.ZN(n2332), 
	.C2(n16951), 
	.C1(n3240), 
	.B2(n16948), 
	.B1(n3239), 
	.A(n3241));
   AOI22_X1 U3093 (.ZN(n3241), 
	.B2(FE_OFN542_n2562), 
	.B1(n16942), 
	.A2(FE_OFN544_n2612), 
	.A1(n16945));
   NAND3_X1 U3095 (.ZN(n3244), 
	.A3(n3246), 
	.A2(n3223), 
	.A1(n5227));
   NAND4_X1 U3096 (.ZN(n2469), 
	.A4(n3249), 
	.A3(n3248), 
	.A2(n3003), 
	.A1(n3247));
   AOI222_X1 U3097 (.ZN(n3249), 
	.C2(n3250), 
	.C1(n16787), 
	.B2(n2879), 
	.B1(hrdata_i[18]), 
	.A2(n2878), 
	.A1(sub_2068_A_18_));
   AOI22_X1 U3099 (.ZN(n3248), 
	.B2(n2344), 
	.B1(n2912), 
	.A2(n2352), 
	.A1(n16645));
   OAI221_X1 U3100 (.ZN(n2344), 
	.C2(n16951), 
	.C1(n3252), 
	.B2(n16948), 
	.B1(n3251), 
	.A(n3253));
   AOI22_X1 U3101 (.ZN(n3253), 
	.B2(n2484), 
	.B1(n16942), 
	.A2(n3254), 
	.A1(n16945));
   OAI221_X1 U3102 (.ZN(n2352), 
	.C2(n16951), 
	.C1(n3256), 
	.B2(n16948), 
	.B1(n3255), 
	.A(n3257));
   AOI22_X1 U3103 (.ZN(n3257), 
	.B2(n2738), 
	.B1(n16942), 
	.A2(n2787), 
	.A1(n16945));
   NAND2_X1 U3104 (.ZN(n2465), 
	.A2(n3259), 
	.A1(n3258));
   AOI221_X1 U3105 (.ZN(n3259), 
	.C2(n2329), 
	.C1(n16645), 
	.B2(n2388), 
	.B1(n2912), 
	.A(n3260));
   OAI22_X1 U3106 (.ZN(n3260), 
	.B2(n3011), 
	.B1(n4748), 
	.A2(n2948), 
	.A1(n5537));
   OAI221_X1 U3107 (.ZN(n2329), 
	.C2(n16951), 
	.C1(n3262), 
	.B2(n16948), 
	.B1(n3261), 
	.A(n3263));
   AOI22_X1 U3108 (.ZN(n3263), 
	.B2(n3022), 
	.B1(n16942), 
	.A2(n3134), 
	.A1(n16945));
   OAI221_X1 U3109 (.ZN(n2388), 
	.C2(n16951), 
	.C1(n3265), 
	.B2(n16948), 
	.B1(n3264), 
	.A(n3266));
   AOI22_X1 U3110 (.ZN(n3266), 
	.B2(n2833), 
	.B1(n16942), 
	.A2(n3267), 
	.A1(n16945));
   AOI222_X1 U3111 (.ZN(n3258), 
	.C2(n3268), 
	.C1(n16787), 
	.B2(n2879), 
	.B1(hrdata_i[10]), 
	.A2(n2878), 
	.A1(sub_2068_A_10_));
   NAND3_X1 U3113 (.ZN(n2002), 
	.A3(n3270), 
	.A2(n3210), 
	.A1(n3269));
   AOI22_X1 U3114 (.ZN(n3270), 
	.B2(n3215), 
	.B1(n1207), 
	.A2(n3246), 
	.A1(n3271));
   NOR2_X1 U3115 (.ZN(n3271), 
	.A2(n3223), 
	.A1(n5227));
   OAI211_X1 U3116 (.ZN(n2468), 
	.C2(n2371), 
	.C1(n3001), 
	.B(FE_PHN4653_n3273), 
	.A(n3272));
   AOI22_X1 U3117 (.ZN(n3273), 
	.B2(n2879), 
	.B1(hrdata_i[26]), 
	.A2(n203), 
	.A1(n2895));
   NAND3_X1 U3118 (.ZN(n3272), 
	.A3(n2922), 
	.A2(n2371), 
	.A1(n2370));
   OAI22_X1 U3119 (.ZN(n2370), 
	.B2(n2337), 
	.B1(n2937), 
	.A2(n16788), 
	.A1(n2874));
   AOI221_X1 U3120 (.ZN(n2937), 
	.C2(n3118), 
	.C1(n2297), 
	.B2(n3275), 
	.B1(n3274), 
	.A(n3276));
   OAI22_X1 U3121 (.ZN(n3276), 
	.B2(n3280), 
	.B1(n3279), 
	.A2(n3278), 
	.A1(n3277));
   INV_X1 U3122 (.ZN(n2874), 
	.A(n2349));
   OAI221_X1 U3123 (.ZN(n2349), 
	.C2(n16951), 
	.C1(n3282), 
	.B2(n16948), 
	.B1(n3281), 
	.A(n3283));
   AOI22_X1 U3124 (.ZN(n3283), 
	.B2(n2402), 
	.B1(n16942), 
	.A2(n2433), 
	.A1(n16945));
   OAI221_X1 U3125 (.ZN(n2371), 
	.C2(n2942), 
	.C1(n3120), 
	.B2(n3119), 
	.B1(n2939), 
	.A(n3122));
   INV_X1 U3126 (.ZN(n2939), 
	.A(n2942));
   NAND3_X1 U3128 (.ZN(n3284), 
	.A3(n3246), 
	.A2(n3223), 
	.A1(n3222));
   NOR3_X1 U3129 (.ZN(n3246), 
	.A3(n3213), 
	.A2(n16843), 
	.A1(n17096));
   OAI22_X1 U3131 (.ZN(U299_Z_0), 
	.B2(n17005), 
	.B1(n3286), 
	.A2(n17001), 
	.A1(FE_PHN2436_n5577));
   OAI22_X1 U3132 (.ZN(U298_Z_0), 
	.B2(n17000), 
	.B1(n3286), 
	.A2(n16996), 
	.A1(FE_PHN2686_n5576));
   OAI22_X1 U3133 (.ZN(U297_Z_0), 
	.B2(n17042), 
	.B1(n3286), 
	.A2(n17038), 
	.A1(FE_PHN2706_n5575));
   OAI22_X1 U3134 (.ZN(U296_Z_0), 
	.B2(n17037), 
	.B1(n3286), 
	.A2(n17033), 
	.A1(FE_PHN2484_n5574));
   OAI22_X1 U3135 (.ZN(U295_Z_0), 
	.B2(n17031), 
	.B1(n3286), 
	.A2(n17028), 
	.A1(n5143));
   OAI22_X1 U3136 (.ZN(U294_Z_0), 
	.B2(FE_OFN651_n17027), 
	.B1(n3286), 
	.A2(n17023), 
	.A1(FE_PHN2663_n5195));
   OAI22_X1 U3137 (.ZN(U293_Z_0), 
	.B2(n17022), 
	.B1(n3286), 
	.A2(n17018), 
	.A1(FE_PHN2499_n5142));
   OAI22_X1 U3138 (.ZN(U292_Z_0), 
	.B2(n17017), 
	.B1(n3286), 
	.A2(n17013), 
	.A1(FE_PHN2598_n5224));
   OAI22_X2 U3139 (.ZN(U291_Z_0), 
	.B2(n17046), 
	.B1(n3286), 
	.A2(n17043), 
	.A1(n5331));
   OAI22_X1 U3140 (.ZN(U290_Z_0), 
	.B2(n17052), 
	.B1(n3286), 
	.A2(n17048), 
	.A1(FE_PHN2626_n5360));
   OAI22_X1 U3142 (.ZN(U289_Z_0), 
	.B2(n17057), 
	.B1(n3286), 
	.A2(n17053), 
	.A1(FE_PHN2443_n5389));
   OAI22_X1 U3143 (.ZN(U288_Z_0), 
	.B2(n17062), 
	.B1(n3286), 
	.A2(n17058), 
	.A1(FE_PHN2640_n5418));
   OAI22_X1 U3144 (.ZN(U287_Z_0), 
	.B2(n17067), 
	.B1(n3286), 
	.A2(n17063), 
	.A1(FE_PHN2682_n5447));
   OAI22_X1 U3145 (.ZN(U286_Z_0), 
	.B2(n17071), 
	.B1(n3286), 
	.A2(n17068), 
	.A1(FE_PHN2674_n5476));
   OAI22_X1 U3146 (.ZN(U285_Z_0), 
	.B2(n17077), 
	.B1(n3286), 
	.A2(n17074), 
	.A1(FE_PHN2776_n5141));
   OAI22_X1 U3147 (.ZN(U284_Z_0), 
	.B2(n17082), 
	.B1(n3286), 
	.A2(n17078), 
	.A1(FE_PHN2453_n5541));
   AOI221_X1 U3149 (.ZN(n2113), 
	.C2(n17008), 
	.C1(n3287), 
	.B2(n16727), 
	.B1(n2495), 
	.A(n3288));
   INV_X1 U3150 (.ZN(n3288), 
	.A(n3289));
   AOI211_X1 U3151 (.ZN(n3289), 
	.C2(n3290), 
	.C1(FE_OFN598_n5805), 
	.B(n3291), 
	.A(n2055));
   NOR3_X1 U3152 (.ZN(n3291), 
	.A3(n1621), 
	.A2(n16992), 
	.A1(FE_OFN598_n5805));
   OAI22_X1 U3153 (.ZN(n3290), 
	.B2(n3292), 
	.B1(n2501), 
	.A2(n1621), 
	.A1(n2131));
   INV_X1 U3154 (.ZN(n1621), 
	.A(n3292));
   NAND4_X1 U3155 (.ZN(n3292), 
	.A4(n3296), 
	.A3(n3295), 
	.A2(n3294), 
	.A1(n3293));
   AOI222_X1 U3156 (.ZN(n3296), 
	.C2(vis_psp_o[7]), 
	.C1(n16969), 
	.B2(n3237), 
	.B1(n16970), 
	.A2(vis_msp_o[7]), 
	.A1(n16975));
   AOI222_X1 U3158 (.ZN(n3295), 
	.C2(vis_r11_o[9]), 
	.C1(n16987), 
	.B2(vis_r12_o[9]), 
	.B1(n16966), 
	.A2(vis_r14_o[9]), 
	.A1(n16984));
   AOI222_X1 U3161 (.ZN(n3294), 
	.C2(vis_r8_o[9]), 
	.C1(FE_PSN5236_n16960), 
	.B2(vis_r10_o[9]), 
	.B1(n16963), 
	.A2(vis_r9_o[9]), 
	.A1(n16979));
   AOI22_X1 U3163 (.ZN(n3293), 
	.B2(n1161), 
	.B1(n16956), 
	.A2(n869), 
	.A1(n16976));
   XOR2_X1 U3165 (.Z(n5805), 
	.B(n3305), 
	.A(n2169));
   AOI221_X1 U3166 (.ZN(n3305), 
	.C2(n3287), 
	.C1(n16988), 
	.B2(n17098), 
	.B1(n2198), 
	.A(n3306));
   OAI22_X1 U3167 (.ZN(n3306), 
	.B2(n2200), 
	.B1(n5258), 
	.A2(n3186), 
	.A1(n5003));
   INV_X1 U3168 (.ZN(n127), 
	.A(n3170));
   OAI221_X1 U3169 (.ZN(n3170), 
	.C2(n2869), 
	.C1(n2473), 
	.B2(n2472), 
	.B1(n3051), 
	.A(n3307));
   AOI221_X1 U3170 (.ZN(n3307), 
	.C2(n2954), 
	.C1(n2005), 
	.B2(n2871), 
	.B1(n2003), 
	.A(n2873));
   NAND3_X1 U3171 (.ZN(n2005), 
	.A3(n3310), 
	.A2(n3309), 
	.A1(n3308));
   AOI221_X1 U3172 (.ZN(n3310), 
	.C2(n2878), 
	.C1(sub_2068_A_1_), 
	.B2(n3311), 
	.B1(n16787), 
	.A(n3312));
   OAI22_X1 U3173 (.ZN(n3312), 
	.B2(n2948), 
	.B1(n5535), 
	.A2(FE_PHN869_n427), 
	.A1(n2918));
   INV_X1 U3174 (.ZN(n427), 
	.A(hrdata_i[1]));
   AOI222_X1 U3176 (.ZN(n3309), 
	.C2(n2326), 
	.C1(n2912), 
	.B2(n3313), 
	.B1(n3058), 
	.A2(n2336), 
	.A1(n16645));
   OAI221_X1 U3177 (.ZN(n2326), 
	.C2(n16951), 
	.C1(n3315), 
	.B2(n16948), 
	.B1(n3314), 
	.A(n3316));
   AOI22_X1 U3178 (.ZN(n3316), 
	.B2(n3317), 
	.B1(n16942), 
	.A2(n2531), 
	.A1(n16945));
   AND2_X1 U3179 (.ZN(n3058), 
	.A2(n1111), 
	.A1(n3318));
   OAI221_X1 U3180 (.ZN(n2336), 
	.C2(n16951), 
	.C1(n3280), 
	.B2(n16948), 
	.B1(n3319), 
	.A(n3320));
   AOI22_X1 U3181 (.ZN(n3320), 
	.B2(FE_OFN543_n2585), 
	.B1(n16942), 
	.A2(FE_OFN560_n3199), 
	.A1(n16945));
   INV_X1 U3182 (.ZN(n3308), 
	.A(n3321));
   OAI22_X1 U3183 (.ZN(n3321), 
	.B2(n5534), 
	.B1(n3011), 
	.A2(n4833), 
	.A1(n3322));
   NAND3_X1 U3184 (.ZN(n2003), 
	.A3(n3325), 
	.A2(n3324), 
	.A1(n3323));
   AOI221_X1 U3185 (.ZN(n3325), 
	.C2(n2878), 
	.C1(sub_2068_A_9_), 
	.B2(n3326), 
	.B1(n16787), 
	.A(n3327));
   OAI22_X1 U3186 (.ZN(n3327), 
	.B2(n2948), 
	.B1(n5578), 
	.A2(n391), 
	.A1(n2918));
   INV_X1 U3187 (.ZN(n391), 
	.A(hrdata_i[9]));
   AOI211_X1 U3189 (.ZN(n3324), 
	.C2(n2330), 
	.C1(n16645), 
	.B(n2897), 
	.A(n3106));
   AND4_X1 U3190 (.ZN(n3106), 
	.A4(n251), 
	.A3(n5096), 
	.A2(n1189), 
	.A1(n3318));
   OAI221_X1 U3191 (.ZN(n2330), 
	.C2(n16951), 
	.C1(n3329), 
	.B2(n16948), 
	.B1(n3328), 
	.A(n3330));
   AOI22_X1 U3192 (.ZN(n3330), 
	.B2(n3041), 
	.B1(n16942), 
	.A2(n3155), 
	.A1(n16945));
   INV_X1 U3193 (.ZN(n3323), 
	.A(n3331));
   OAI22_X1 U3194 (.ZN(n3331), 
	.B2(n5011), 
	.B1(n3011), 
	.A2(n2378), 
	.A1(n2875));
   INV_X1 U3195 (.ZN(n2378), 
	.A(n2988));
   OAI221_X1 U3196 (.ZN(n2988), 
	.C2(n16951), 
	.C1(n3333), 
	.B2(n16948), 
	.B1(n3332), 
	.A(n3334));
   AOI22_X1 U3197 (.ZN(n3334), 
	.B2(n2856), 
	.B1(n16942), 
	.A2(n2964), 
	.A1(n16945));
   INV_X1 U3198 (.ZN(n2869), 
	.A(n2977));
   INV_X1 U3199 (.ZN(n2473), 
	.A(n2009));
   OAI211_X1 U3200 (.ZN(n2009), 
	.C2(n3335), 
	.C1(n3001), 
	.B(n3336), 
	.A(n3003));
   INV_X1 U3201 (.ZN(n3336), 
	.A(n3337));
   OAI22_X1 U3202 (.ZN(n3337), 
	.B2(n2918), 
	.B1(FE_PHN763_n1140), 
	.A2(n2998), 
	.A1(n2372));
   INV_X1 U3203 (.ZN(n1140), 
	.A(hrdata_i[25]));
   OAI221_X1 U3204 (.ZN(n2372), 
	.C2(FE_OFN533_n2357), 
	.C1(n16788), 
	.B2(n3004), 
	.B1(n2337), 
	.A(n3335));
   OAI221_X1 U3205 (.ZN(n2357), 
	.C2(n16951), 
	.C1(n3339), 
	.B2(n16948), 
	.B1(n3338), 
	.A(n3340));
   AOI22_X1 U3206 (.ZN(n3340), 
	.B2(n2271), 
	.B1(n16942), 
	.A2(n2452), 
	.A1(n16945));
   OAI221_X1 U3207 (.ZN(n3004), 
	.C2(n16951), 
	.C1(n3341), 
	.B2(n16948), 
	.B1(n3278), 
	.A(n3342));
   AOI22_X1 U3208 (.ZN(n3342), 
	.B2(n3274), 
	.B1(n16942), 
	.A2(n2297), 
	.A1(n16945));
   OAI221_X1 U3209 (.ZN(n3335), 
	.C2(n3006), 
	.C1(n3120), 
	.B2(n3119), 
	.B1(n3005), 
	.A(n3122));
   AOI21_X1 U3210 (.ZN(n3122), 
	.B2(n2337), 
	.B1(n3343), 
	.A(FE_OFN631_n16851));
   INV_X1 U3211 (.ZN(n3006), 
	.A(n3005));
   NAND2_X1 U3212 (.ZN(n3005), 
	.A2(n16948), 
	.A1(n2942));
   NOR2_X1 U3213 (.ZN(n2942), 
	.A2(n16945), 
	.A1(n3118));
   NAND2_X1 U3214 (.ZN(n3001), 
	.A2(n2922), 
	.A1(n2313));
   INV_X1 U3215 (.ZN(n2472), 
	.A(n2010));
   OAI221_X1 U3216 (.ZN(n2010), 
	.C2(n278), 
	.C1(n2981), 
	.B2(n16685), 
	.B1(FE_PHN2364_n5639), 
	.A(FE_PHN727_n3344));
   AOI222_X1 U3217 (.ZN(n3344), 
	.C2(n2345), 
	.C1(n2912), 
	.B2(n2353), 
	.B1(n16645), 
	.A2(n2879), 
	.A1(hrdata_i[17]));
   OAI221_X1 U3218 (.ZN(n2345), 
	.C2(n16951), 
	.C1(n3346), 
	.B2(n16948), 
	.B1(n3345), 
	.A(n3347));
   AOI22_X1 U3219 (.ZN(n3347), 
	.B2(n2507), 
	.B1(n16942), 
	.A2(n2705), 
	.A1(n16945));
   NAND2_X1 U3221 (.ZN(n2875), 
	.A2(n16788), 
	.A1(n2922));
   OAI221_X1 U3222 (.ZN(n2353), 
	.C2(n16951), 
	.C1(n3349), 
	.B2(n16948), 
	.B1(n3348), 
	.A(n3350));
   AOI22_X1 U3223 (.ZN(n3350), 
	.B2(n2764), 
	.B1(n16942), 
	.A2(n2809), 
	.A1(n16945));
   INV_X1 U3226 (.ZN(n3051), 
	.A(n2872));
   OAI22_X1 U3227 (.ZN(U283_Z_0), 
	.B2(n17005), 
	.B1(n3351), 
	.A2(n17001), 
	.A1(FE_PHN2561_n5139));
   OAI22_X1 U3228 (.ZN(U282_Z_0), 
	.B2(n17000), 
	.B1(n3351), 
	.A2(n16996), 
	.A1(FE_PHN2731_n5138));
   OAI22_X1 U3229 (.ZN(U281_Z_0), 
	.B2(n17042), 
	.B1(n3351), 
	.A2(FE_OFN654_n17038), 
	.A1(FE_PHN2661_n5304));
   OAI22_X1 U3230 (.ZN(U280_Z_0), 
	.B2(n17037), 
	.B1(n3351), 
	.A2(FE_OFN652_n17033), 
	.A1(FE_PHN2528_n5283));
   OAI22_X1 U3231 (.ZN(U279_Z_0), 
	.B2(n17031), 
	.B1(n3351), 
	.A2(n17028), 
	.A1(n5137));
   OAI22_X1 U3232 (.ZN(U278_Z_0), 
	.B2(n17027), 
	.B1(n3351), 
	.A2(n17023), 
	.A1(FE_PHN2763_n5196));
   OAI22_X1 U3233 (.ZN(U277_Z_0), 
	.B2(n17022), 
	.B1(n3351), 
	.A2(n17018), 
	.A1(FE_PHN2569_n5136));
   OAI22_X1 U3234 (.ZN(U276_Z_0), 
	.B2(FE_OFN648_n17017), 
	.B1(n3351), 
	.A2(n17013), 
	.A1(FE_PHN2588_n5225));
   OAI22_X2 U3235 (.ZN(U275_Z_0), 
	.B2(n17046), 
	.B1(n3351), 
	.A2(n17043), 
	.A1(n5332));
   OAI22_X1 U3236 (.ZN(U274_Z_0), 
	.B2(n17052), 
	.B1(n3351), 
	.A2(n17048), 
	.A1(FE_PHN2599_n5361));
   OAI22_X1 U3237 (.ZN(U273_Z_0), 
	.B2(n17057), 
	.B1(n3351), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2444_n5390));
   OAI22_X1 U3238 (.ZN(U272_Z_0), 
	.B2(n17062), 
	.B1(n3351), 
	.A2(FE_OFN663_n17058), 
	.A1(FE_PHN2632_n5419));
   OAI22_X1 U3239 (.ZN(U271_Z_0), 
	.B2(n17067), 
	.B1(n3351), 
	.A2(n17063), 
	.A1(FE_PHN2658_n5448));
   OAI22_X1 U3240 (.ZN(U270_Z_0), 
	.B2(n17071), 
	.B1(n3351), 
	.A2(n17068), 
	.A1(FE_PHN2724_n5477));
   OAI22_X1 U3242 (.ZN(U269_Z_0), 
	.B2(FE_OFN666_n17077), 
	.B1(n3351), 
	.A2(n17074), 
	.A1(FE_PHN2737_n5135));
   OAI22_X1 U3243 (.ZN(U268_Z_0), 
	.B2(n17082), 
	.B1(n3351), 
	.A2(n17078), 
	.A1(FE_PHN2516_n5542));
   AOI221_X1 U3245 (.ZN(n3353), 
	.C2(FE_OFN208_n2015), 
	.C1(n16722), 
	.B2(n2261), 
	.B1(n17008), 
	.A(n2055));
   OAI221_X1 U3246 (.ZN(n3352), 
	.C2(n2148), 
	.C1(n16994), 
	.B2(n5819), 
	.B1(n3354), 
	.A(n3355));
   NAND3_X1 U3247 (.ZN(n3355), 
	.A3(n5819), 
	.A2(n2148), 
	.A1(n2131));
   AOI221_X1 U3249 (.ZN(n3356), 
	.C2(n2261), 
	.C1(n16988), 
	.B2(n16798), 
	.B1(n2198), 
	.A(n3357));
   OAI22_X1 U3250 (.ZN(n3357), 
	.B2(n2200), 
	.B1(n5257), 
	.A2(n3186), 
	.A1(FE_OFN587_n5162));
   OAI21_X1 U3251 (.ZN(n2200), 
	.B2(n3359), 
	.B1(n3358), 
	.A(FE_OFN10_n1697));
   OAI22_X1 U3252 (.ZN(n3359), 
	.B2(n3361), 
	.B1(n758), 
	.A2(n745), 
	.A1(n3360));
   NAND2_X1 U3253 (.ZN(n3361), 
	.A2(n991), 
	.A1(n16851));
   NOR3_X1 U3254 (.ZN(n3360), 
	.A3(n798), 
	.A2(n760), 
	.A1(n16847));
   INV_X1 U3255 (.ZN(n798), 
	.A(n3362));
   OAI33_X1 U3256 (.ZN(n3358), 
	.B3(n3362), 
	.B2(n16851), 
	.B1(n863), 
	.A3(n653), 
	.A2(FE_OFN100_n1086), 
	.A1(n3363));
   NAND2_X1 U3257 (.ZN(n863), 
	.A2(n16860), 
	.A1(n991));
   NOR2_X1 U3258 (.ZN(n3354), 
	.A2(n16992), 
	.A1(n1625));
   INV_X1 U3259 (.ZN(n1625), 
	.A(n2148));
   NAND4_X1 U3260 (.ZN(n2148), 
	.A4(n3367), 
	.A3(n3366), 
	.A2(n3365), 
	.A1(n3364));
   AOI222_X1 U3261 (.ZN(n3367), 
	.C2(vis_psp_o[6]), 
	.C1(n16969), 
	.B2(n3317), 
	.B1(n16970), 
	.A2(vis_msp_o[6]), 
	.A1(n16975));
   AOI222_X1 U3263 (.ZN(n3366), 
	.C2(vis_r11_o[8]), 
	.C1(n16987), 
	.B2(vis_r12_o[8]), 
	.B1(n16966), 
	.A2(vis_r14_o[8]), 
	.A1(n16983));
   AOI222_X1 U3266 (.ZN(n3365), 
	.C2(vis_r8_o[8]), 
	.C1(FE_PSN5236_n16960), 
	.B2(vis_r10_o[8]), 
	.B1(n16963), 
	.A2(vis_r9_o[8]), 
	.A1(n16979));
   AOI22_X1 U3268 (.ZN(n3364), 
	.B2(n2221), 
	.B1(n16956), 
	.A2(n1161), 
	.A1(n16976));
   AOI221_X1 U3270 (.ZN(n144), 
	.C2(n2954), 
	.C1(n2018), 
	.B2(n2977), 
	.B1(n2022), 
	.A(n3376));
   INV_X2 U3271 (.ZN(n3376), 
	.A(n3377));
   AOI221_X1 U3272 (.ZN(n3377), 
	.C2(n2872), 
	.C1(n2023), 
	.B2(n2019), 
	.B1(n2871), 
	.A(n2873));
   NAND4_X1 U3273 (.ZN(n2023), 
	.A4(n3380), 
	.A3(n3379), 
	.A2(n3003), 
	.A1(n3378));
   AOI222_X1 U3274 (.ZN(n3380), 
	.C2(n3381), 
	.C1(n16787), 
	.B2(n2879), 
	.B1(hrdata_i[16]), 
	.A2(n2878), 
	.A1(sub_2068_A_16_));
   INV_X1 U3276 (.ZN(n3379), 
	.A(n3382));
   OAI22_X1 U3277 (.ZN(n3382), 
	.B2(n5068), 
	.B1(n3322), 
	.A2(n2998), 
	.A1(n1779));
   OAI22_X1 U3278 (.ZN(n1779), 
	.B2(n2385), 
	.B1(n16788), 
	.A2(n2355), 
	.A1(n2337));
   OAI221_X1 U3279 (.ZN(n2385), 
	.C2(n16951), 
	.C1(n3264), 
	.B2(n16948), 
	.B1(n3256), 
	.A(n3383));
   AOI22_X1 U3280 (.ZN(n3383), 
	.B2(n2787), 
	.B1(n16942), 
	.A2(n2833), 
	.A1(n16945));
   OAI221_X1 U3281 (.ZN(n2355), 
	.C2(n16951), 
	.C1(n3255), 
	.B2(n16948), 
	.B1(n3252), 
	.A(n3384));
   AOI22_X1 U3282 (.ZN(n3384), 
	.B2(n3254), 
	.B1(n16942), 
	.A2(n2738), 
	.A1(n16945));
   NAND2_X1 U3283 (.ZN(n3378), 
	.A2(n2895), 
	.A1(n405));
   INV_X1 U3284 (.ZN(n405), 
	.A(n421));
   NAND3_X1 U3285 (.ZN(n421), 
	.A3(n2905), 
	.A2(n1372), 
	.A1(n2907));
   INV_X1 U3286 (.ZN(n2019), 
	.A(n3385));
   AOI211_X1 U3287 (.ZN(n3385), 
	.C2(sub_2068_A_8_), 
	.C1(n2878), 
	.B(n3387), 
	.A(n3386));
   OAI222_X1 U3288 (.ZN(n3387), 
	.C2(n2918), 
	.C1(FE_PHN904_n393), 
	.B2(n4796), 
	.B1(n2948), 
	.A2(n4747), 
	.A1(n3011));
   INV_X1 U3289 (.ZN(n393), 
	.A(hrdata_i[8]));
   OAI22_X1 U3290 (.ZN(n3386), 
	.B2(FE_PHN2426_n5581), 
	.B1(n16685), 
	.A2(n2998), 
	.A1(n1772));
   OAI22_X1 U3291 (.ZN(n1772), 
	.B2(n2339), 
	.B1(n16788), 
	.A2(n2387), 
	.A1(n2337));
   OAI221_X1 U3292 (.ZN(n2339), 
	.C2(n16951), 
	.C1(n3231), 
	.B2(n16948), 
	.B1(n3262), 
	.A(n3388));
   AOI22_X1 U3293 (.ZN(n3388), 
	.B2(n3134), 
	.B1(n16942), 
	.A2(n3237), 
	.A1(n16945));
   OAI221_X1 U3294 (.ZN(n2387), 
	.C2(n16951), 
	.C1(n3261), 
	.B2(n16948), 
	.B1(n3265), 
	.A(n3389));
   AOI22_X1 U3295 (.ZN(n3389), 
	.B2(n3267), 
	.B1(n16942), 
	.A2(n3022), 
	.A1(n16945));
   INV_X1 U3297 (.ZN(n2018), 
	.A(n2517));
   NOR2_X1 U3298 (.ZN(n2517), 
	.A2(n3391), 
	.A1(n3390));
   OAI221_X1 U3299 (.ZN(n3391), 
	.C2(n2998), 
	.C1(n1781), 
	.B2(FE_PHN3501_n5516), 
	.B1(n3322), 
	.A(n3392));
   INV_X1 U3300 (.ZN(n3392), 
	.A(n3393));
   OAI22_X1 U3301 (.ZN(n3393), 
	.B2(n3011), 
	.B1(n5005), 
	.A2(n2948), 
	.A1(n5540));
   OAI22_X1 U3302 (.ZN(n1781), 
	.B2(n3094), 
	.B1(n16788), 
	.A2(n2333), 
	.A1(n2337));
   OAI221_X1 U3303 (.ZN(n3094), 
	.C2(n16951), 
	.C1(n2183), 
	.B2(n16948), 
	.B1(n3240), 
	.A(n3394));
   AOI22_X1 U3304 (.ZN(n3394), 
	.B2(FE_OFN544_n2612), 
	.B1(n16942), 
	.A2(n2639), 
	.A1(n16945));
   OAI221_X1 U3305 (.ZN(n2333), 
	.C2(n16951), 
	.C1(n3239), 
	.B2(n3279), 
	.B1(n3314), 
	.A(n3395));
   AOI22_X1 U3306 (.ZN(n3395), 
	.B2(n2531), 
	.B1(n3275), 
	.A2(FE_OFN542_n2562), 
	.A1(n16945));
   INV_X1 U3307 (.ZN(n3322), 
	.A(n3230));
   NOR3_X1 U3308 (.ZN(n3230), 
	.A3(n261), 
	.A2(n2926), 
	.A1(n251));
   OAI222_X1 U3309 (.ZN(n3390), 
	.C2(FE_PHN3512_n5510), 
	.C1(n16685), 
	.B2(n2918), 
	.B1(FE_PHN804_n429), 
	.A2(n2981), 
	.A1(n260));
   INV_X1 U3310 (.ZN(n429), 
	.A(hrdata_i[0]));
   INV_X1 U3311 (.ZN(n2022), 
	.A(FE_PHN685_n2516));
   AOI221_X1 U3312 (.ZN(n2516), 
	.C2(n2922), 
	.C1(n2363), 
	.B2(hrdata_i[24]), 
	.B1(n2879), 
	.A(n2897));
   OAI22_X1 U3313 (.ZN(n2363), 
	.B2(n3397), 
	.B1(n3092), 
	.A2(n3396), 
	.A1(n1782));
   INV_X1 U3314 (.ZN(n3396), 
	.A(n3397));
   NAND2_X1 U3315 (.ZN(n3397), 
	.A2(FE_OFN90_n16849), 
	.A1(n3120));
   AOI22_X1 U3316 (.ZN(n1782), 
	.B2(n16788), 
	.B1(n3095), 
	.A2(n2337), 
	.A1(n2350));
   OAI221_X1 U3317 (.ZN(n3095), 
	.C2(n16951), 
	.C1(n3281), 
	.B2(n16948), 
	.B1(n3398), 
	.A(n3399));
   AOI22_X1 U3318 (.ZN(n3399), 
	.B2(n3400), 
	.B1(n16942), 
	.A2(n2402), 
	.A1(n16945));
   OAI221_X1 U3319 (.ZN(n2350), 
	.C2(n16951), 
	.C1(n3251), 
	.B2(n16948), 
	.B1(n3282), 
	.A(n3401));
   AOI22_X1 U3320 (.ZN(n3401), 
	.B2(n2433), 
	.B1(n16942), 
	.A2(n2484), 
	.A1(n16945));
   OAI22_X1 U3321 (.ZN(U265_Z_0), 
	.B2(n17005), 
	.B1(n3402), 
	.A2(n17001), 
	.A1(FE_PHN2529_n5634));
   OAI22_X1 U3322 (.ZN(U264_Z_0), 
	.B2(n17000), 
	.B1(n3402), 
	.A2(n16996), 
	.A1(FE_PHN2754_n5633));
   OAI22_X1 U3323 (.ZN(U263_Z_0), 
	.B2(n17042), 
	.B1(n3402), 
	.A2(n17038), 
	.A1(n5632));
   OAI22_X1 U3324 (.ZN(U262_Z_0), 
	.B2(n17037), 
	.B1(n3402), 
	.A2(FE_OFN652_n17033), 
	.A1(FE_PHN2478_n5631));
   OAI22_X1 U3325 (.ZN(U261_Z_0), 
	.B2(n17031), 
	.B1(n3402), 
	.A2(n17028), 
	.A1(n5110));
   OAI22_X1 U3326 (.ZN(U260_Z_0), 
	.B2(n17027), 
	.B1(n3402), 
	.A2(n17023), 
	.A1(FE_PHN2703_n5197));
   OAI22_X1 U3328 (.ZN(U259_Z_0), 
	.B2(n17022), 
	.B1(n3402), 
	.A2(n17018), 
	.A1(FE_PHN2538_n5109));
   OAI22_X1 U3329 (.ZN(U258_Z_0), 
	.B2(FE_OFN648_n17017), 
	.B1(n3402), 
	.A2(n17013), 
	.A1(FE_PHN2483_n5226));
   OAI22_X1 U3330 (.ZN(U257_Z_0), 
	.B2(n17046), 
	.B1(n3402), 
	.A2(n17043), 
	.A1(n5333));
   OAI22_X1 U3331 (.ZN(U256_Z_0), 
	.B2(n17052), 
	.B1(n3402), 
	.A2(FE_OFN656_n17048), 
	.A1(FE_PHN2600_n5362));
   OAI22_X1 U3332 (.ZN(U255_Z_0), 
	.B2(n17057), 
	.B1(n3402), 
	.A2(FE_OFN659_n17053), 
	.A1(FE_PHN2512_n5391));
   OAI22_X1 U3333 (.ZN(U254_Z_0), 
	.B2(n17062), 
	.B1(n3402), 
	.A2(FE_OFN663_n17058), 
	.A1(FE_PHN2740_n5420));
   OAI22_X1 U3334 (.ZN(U253_Z_0), 
	.B2(n17067), 
	.B1(n3402), 
	.A2(n17063), 
	.A1(FE_PHN2702_n5449));
   OAI22_X1 U3335 (.ZN(U252_Z_0), 
	.B2(n17071), 
	.B1(n3402), 
	.A2(n17068), 
	.A1(FE_PHN2768_n5478));
   OAI22_X1 U3336 (.ZN(U251_Z_0), 
	.B2(FE_OFN666_n17077), 
	.B1(n3402), 
	.A2(n17074), 
	.A1(FE_PHN2681_n5108));
   OAI22_X1 U3337 (.ZN(U250_Z_0), 
	.B2(n17082), 
	.B1(n3402), 
	.A2(n17078), 
	.A1(FE_PHN2518_n5543));
   AOI221_X1 U3339 (.ZN(n3404), 
	.C2(FE_OFN208_n2015), 
	.C1(n16715), 
	.B2(n2254), 
	.B1(n17008), 
	.A(n2055));
   OAI221_X1 U3340 (.ZN(n3403), 
	.C2(n2144), 
	.C1(n16994), 
	.B2(n5818), 
	.B1(n3405), 
	.A(n3406));
   NAND3_X1 U3341 (.ZN(n3406), 
	.A3(n5818), 
	.A2(n2144), 
	.A1(n2131));
   AOI221_X1 U3343 (.ZN(n3407), 
	.C2(FE_OFN15_n16671), 
	.C1(n2198), 
	.B2(n2254), 
	.B1(n16989), 
	.A(n2732));
   NOR2_X1 U3344 (.ZN(n3405), 
	.A2(n16992), 
	.A1(n1661));
   INV_X1 U3345 (.ZN(n1661), 
	.A(n2144));
   NAND4_X1 U3346 (.ZN(n2144), 
	.A4(n3411), 
	.A3(n3410), 
	.A2(n3409), 
	.A1(n3408));
   AOI222_X1 U3347 (.ZN(n3411), 
	.C2(vis_psp_o[13]), 
	.C1(n16969), 
	.B2(n3267), 
	.B1(n16970), 
	.A2(vis_msp_o[13]), 
	.A1(n16975));
   AOI222_X1 U3349 (.ZN(n3410), 
	.C2(vis_r11_o[15]), 
	.C1(n16987), 
	.B2(vis_r12_o[15]), 
	.B1(n16966), 
	.A2(vis_r14_o[15]), 
	.A1(n16984));
   AOI222_X1 U3352 (.ZN(n3409), 
	.C2(vis_r8_o[15]), 
	.C1(FE_PSN5236_n16960), 
	.B2(vis_r10_o[15]), 
	.B1(n16963), 
	.A2(vis_r9_o[15]), 
	.A1(n16979));
   AOI22_X1 U3354 (.ZN(n3408), 
	.B2(n2961), 
	.B1(n16956), 
	.A2(n1163), 
	.A1(n16976));
   AOI221_X1 U3357 (.ZN(n48), 
	.C2(FE_PSN5239_n2057), 
	.C1(n2977), 
	.B2(n2061), 
	.B1(n2872), 
	.A(n3420));
   INV_X2 U3358 (.ZN(n3420), 
	.A(n3421));
   AOI221_X1 U3359 (.ZN(n3421), 
	.C2(n2058), 
	.C1(n2871), 
	.B2(n2062), 
	.B1(n2954), 
	.A(n2873));
   INV_X4 U3360 (.ZN(n2873), 
	.A(n3422));
   OAI211_X1 U3361 (.ZN(n3422), 
	.C2(n3215), 
	.C1(n2377), 
	.B(n3424), 
	.A(n3423));
   NOR2_X2 U3362 (.ZN(n3424), 
	.A2(n3425), 
	.A1(n3214));
   NAND4_X1 U3363 (.ZN(n3423), 
	.A4(n3426), 
	.A3(1'b1), 
	.A2(n1518), 
	.A1(n3215));
   NAND3_X1 U3364 (.ZN(n3426), 
	.A3(n195), 
	.A2(n16871), 
	.A1(n16837));
   AOI211_X1 U3365 (.ZN(n2377), 
	.C2(n2358), 
	.C1(n2341), 
	.B(n2322), 
	.A(n2321));
   INV_X1 U3367 (.ZN(n2756), 
	.A(n2720));
   AOI211_X1 U3368 (.ZN(n3427), 
	.C2(n3428), 
	.C1(n5102), 
	.B(n728), 
	.A(n1712));
   INV_X4 U3369 (.ZN(n728), 
	.A(n605));
   NOR2_X1 U3370 (.ZN(n1712), 
	.A2(n16851), 
	.A1(n1210));
   NAND2_X1 U3371 (.ZN(n1210), 
	.A2(n16860), 
	.A1(n16842));
   OAI21_X1 U3372 (.ZN(n3428), 
	.B2(n1580), 
	.B1(FE_OFN84_n16839), 
	.A(n3429));
   NAND2_X1 U3373 (.ZN(n2954), 
	.A2(n3269), 
	.A1(n2417));
   NAND3_X1 U3374 (.ZN(n3269), 
	.A3(n3215), 
	.A2(n3430), 
	.A1(n827));
   INV_X1 U3375 (.ZN(n2417), 
	.A(n2067));
   NAND3_X1 U3376 (.ZN(n2977), 
	.A3(n3431), 
	.A2(n3245), 
	.A1(n3243));
   NAND3_X1 U3377 (.ZN(n3431), 
	.A3(n3432), 
	.A2(n3223), 
	.A1(n3215));
   NAND4_X1 U3378 (.ZN(n3245), 
	.A4(n16843), 
	.A3(n3223), 
	.A2(n990), 
	.A1(n3215));
   INV_X1 U3379 (.ZN(n990), 
	.A(n1964));
   NAND2_X1 U3380 (.ZN(n2872), 
	.A2(n3210), 
	.A1(n3285));
   NAND2_X1 U3381 (.ZN(n3210), 
	.A2(n2341), 
	.A1(n3433));
   OAI22_X1 U3382 (.ZN(U247_Z_0), 
	.B2(n17005), 
	.B1(n3434), 
	.A2(n17001), 
	.A1(n5595));
   OAI22_X1 U3385 (.ZN(U246_Z_0), 
	.B2(n17000), 
	.B1(n3434), 
	.A2(n16996), 
	.A1(n4970));
   OAI22_X1 U3388 (.ZN(U245_Z_0), 
	.B2(n17042), 
	.B1(n3434), 
	.A2(n17038), 
	.A1(FE_PHN3648_n5594));
   OAI22_X1 U3391 (.ZN(U244_Z_0), 
	.B2(n17037), 
	.B1(n3434), 
	.A2(n17033), 
	.A1(FE_PHN3551_n5593));
   AND2_X1 U3394 (.ZN(n3437), 
	.A2(n3441), 
	.A1(n3440));
   OAI22_X1 U3395 (.ZN(U243_Z_0), 
	.B2(n17031), 
	.B1(n3434), 
	.A2(n17028), 
	.A1(n4960));
   OAI22_X1 U3398 (.ZN(U242_Z_0), 
	.B2(n17027), 
	.B1(n3434), 
	.A2(n17023), 
	.A1(n5592));
   OAI22_X1 U3401 (.ZN(U241_Z_0), 
	.B2(n17022), 
	.B1(n3434), 
	.A2(n17018), 
	.A1(FE_PHN3558_n5591));
   OAI22_X1 U3404 (.ZN(U240_Z_0), 
	.B2(n17017), 
	.B1(n3434), 
	.A2(n17013), 
	.A1(FE_PHN3572_n5590));
   AND2_X1 U3407 (.ZN(n3442), 
	.A2(n3441), 
	.A1(n3444));
   OAI22_X1 U3408 (.ZN(U239_Z_0), 
	.B2(n17046), 
	.B1(n3434), 
	.A2(n17043), 
	.A1(n5589));
   OAI22_X1 U3411 (.ZN(U238_Z_0), 
	.B2(n17052), 
	.B1(n3434), 
	.A2(n17048), 
	.A1(FE_PHN3590_n5588));
   OAI22_X1 U3414 (.ZN(U237_Z_0), 
	.B2(n17057), 
	.B1(n3434), 
	.A2(n17053), 
	.A1(FE_PHN3574_n5587));
   OAI22_X1 U3417 (.ZN(U236_Z_0), 
	.B2(n17062), 
	.B1(n3434), 
	.A2(n17058), 
	.A1(FE_PHN4739_n5586));
   NOR2_X1 U3420 (.ZN(n3445), 
	.A2(n3444), 
	.A1(n3441));
   INV_X1 U3421 (.ZN(n3444), 
	.A(n3440));
   OAI22_X1 U3422 (.ZN(U235_Z_0), 
	.B2(n17067), 
	.B1(n3434), 
	.A2(n17063), 
	.A1(n5585));
   AND2_X1 U3425 (.ZN(n3443), 
	.A2(n3448), 
	.A1(n3447));
   OAI22_X1 U3426 (.ZN(U234_Z_0), 
	.B2(n17071), 
	.B1(n3434), 
	.A2(n17068), 
	.A1(n5584));
   AND2_X1 U3429 (.ZN(n3438), 
	.A2(n3448), 
	.A1(n3449));
   OAI22_X1 U3430 (.ZN(U233_Z_0), 
	.B2(n17077), 
	.B1(n3434), 
	.A2(n17074), 
	.A1(n4983));
   NOR2_X1 U3433 (.ZN(n3435), 
	.A2(n3449), 
	.A1(n3448));
   INV_X1 U3434 (.ZN(n3449), 
	.A(n3447));
   OAI22_X1 U3435 (.ZN(U232_Z_0), 
	.B2(n17082), 
	.B1(n3434), 
	.A2(n17078), 
	.A1(FE_PHN3603_n5583));
   AOI221_X1 U3437 (.ZN(n2103), 
	.C2(n17008), 
	.C1(n3450), 
	.B2(n16705), 
	.B1(n2495), 
	.A(n3451));
   INV_X1 U3438 (.ZN(n3451), 
	.A(n3452));
   AOI211_X1 U3439 (.ZN(n3452), 
	.C2(n3453), 
	.C1(n5803), 
	.B(n3454), 
	.A(n2055));
   NOR3_X1 U3440 (.ZN(n3454), 
	.A3(n1685), 
	.A2(n16992), 
	.A1(n5803));
   OAI22_X1 U3441 (.ZN(n3453), 
	.B2(n1649), 
	.B1(FE_OFN538_n2501), 
	.A2(n1685), 
	.A1(n2131));
   INV_X1 U3442 (.ZN(n1685), 
	.A(n1649));
   NAND4_X1 U3443 (.ZN(n1649), 
	.A4(n3458), 
	.A3(n3457), 
	.A2(n3456), 
	.A1(n3455));
   AOI222_X1 U3444 (.ZN(n3458), 
	.C2(vis_psp_o[21]), 
	.C1(n16969), 
	.B2(n3254), 
	.B1(n16970), 
	.A2(vis_msp_o[21]), 
	.A1(n16975));
   AOI222_X1 U3446 (.ZN(n3457), 
	.C2(vis_r11_o[23]), 
	.C1(n16987), 
	.B2(vis_r12_o[23]), 
	.B1(FE_OFN109_n16964), 
	.A2(vis_r14_o[23]), 
	.A1(n16984));
   AOI222_X1 U3449 (.ZN(n3456), 
	.C2(vis_r8_o[23]), 
	.C1(FE_PSN5236_n16960), 
	.B2(vis_r10_o[23]), 
	.B1(n16961), 
	.A2(vis_r9_o[23]), 
	.A1(n16979));
   AOI22_X1 U3451 (.ZN(n3455), 
	.B2(n2713), 
	.B1(n16956), 
	.A2(n2515), 
	.A1(n16976));
   XOR2_X1 U3455 (.Z(n5803), 
	.B(n3467), 
	.A(n16990));
   AOI221_X1 U3456 (.ZN(n3467), 
	.C2(n3450), 
	.C1(n16988), 
	.B2(n16683), 
	.B1(n2716), 
	.A(n3468));
   NAND2_X1 U3457 (.ZN(n3468), 
	.A2(n2719), 
	.A1(n3469));
   NAND3_X1 U3458 (.ZN(n3469), 
	.A3(n16807), 
	.A2(n2198), 
	.A1(n5254));
   INV_X1 U3460 (.ZN(n2495), 
	.A(n2544));
   NOR2_X1 U3461 (.ZN(n2544), 
	.A2(n2055), 
	.A1(FE_OFN2_n2015));
   AOI221_X1 U3462 (.ZN(n44), 
	.C2(n2074), 
	.C1(n2062), 
	.B2(FE_PSN5239_n2057), 
	.B1(n2749), 
	.A(n3470));
   INV_X1 U3463 (.ZN(n3470), 
	.A(n3471));
   AOI221_X1 U3464 (.ZN(n3471), 
	.C2(n2061), 
	.C1(n2720), 
	.B2(n2721), 
	.B1(n2058), 
	.A(n71));
   AND4_X4 U3465 (.ZN(n71), 
	.A4(n3474), 
	.A3(n3211), 
	.A2(n3473), 
	.A1(n3472));
   NOR3_X1 U3466 (.ZN(n3474), 
	.A3(n2074), 
	.A2(n3433), 
	.A1(n3425));
   INV_X1 U3467 (.ZN(n3433), 
	.A(n3475));
   NAND2_X1 U3468 (.ZN(n2720), 
	.A2(n3211), 
	.A1(n3476));
   NAND2_X1 U3469 (.ZN(n3211), 
	.A2(n3213), 
	.A1(n2321));
   NOR2_X1 U3470 (.ZN(n2321), 
	.A2(n3242), 
	.A1(n3477));
   INV_X1 U3471 (.ZN(n3242), 
	.A(n2341));
   NAND2_X1 U3472 (.ZN(n2341), 
	.A2(n3478), 
	.A1(n16828));
   NAND2_X1 U3473 (.ZN(n2721), 
	.A2(n3285), 
	.A1(n3472));
   OAI21_X1 U3474 (.ZN(n2749), 
	.B2(n1027), 
	.B1(n3213), 
	.A(n3475));
   NOR2_X1 U3477 (.ZN(n3439), 
	.A2(n3448), 
	.A1(n3447));
   NAND3_X1 U3478 (.ZN(n3448), 
	.A3(n1350), 
	.A2(n3479), 
	.A1(n17122));
   AOI221_X1 U3479 (.ZN(n1350), 
	.C2(n3482), 
	.C1(n1353), 
	.B2(n3481), 
	.B1(n3480), 
	.A(n3483));
   OAI21_X1 U3480 (.ZN(n3483), 
	.B2(n5003), 
	.B1(n3484), 
	.A(n3485));
   OAI211_X1 U3481 (.ZN(n3447), 
	.C2(n3484), 
	.C1(n5162), 
	.B(n3487), 
	.A(n3486));
   AOI22_X1 U3482 (.ZN(n3487), 
	.B2(n3489), 
	.B1(n3482), 
	.A2(n3488), 
	.A1(n3481));
   INV_X1 U3483 (.ZN(n3484), 
	.A(n3490));
   NOR2_X1 U3484 (.ZN(n3446), 
	.A2(n3441), 
	.A1(n3440));
   NAND3_X1 U3485 (.ZN(n3441), 
	.A3(n3491), 
	.A2(n3485), 
	.A1(n3486));
   AOI222_X1 U3486 (.ZN(n3491), 
	.C2(n3493), 
	.C1(n3482), 
	.B2(n3492), 
	.B1(n3481), 
	.A2(n2731), 
	.A1(n3490));
   NAND3_X1 U3487 (.ZN(n3440), 
	.A3(n3494), 
	.A2(n3485), 
	.A1(n3486));
   AOI222_X1 U3488 (.ZN(n3494), 
	.C2(n3496), 
	.C1(n3482), 
	.B2(n3495), 
	.B1(n3481), 
	.A2(n1723), 
	.A1(n3490));
   OAI211_X1 U3489 (.ZN(n3482), 
	.C2(n699), 
	.C1(n16854), 
	.B(n3498), 
	.A(n3497));
   NAND4_X1 U3490 (.ZN(n3498), 
	.A4(FE_OFN72_n16867), 
	.A3(FE_OFN85_n16839), 
	.A2(n757), 
	.A1(n611));
   INV_X1 U3491 (.ZN(n611), 
	.A(n1211));
   NAND2_X1 U3492 (.ZN(n1211), 
	.A2(n16851), 
	.A1(n16845));
   NAND4_X1 U3493 (.ZN(n3497), 
	.A4(n16833), 
	.A3(FE_OFN633_n16868), 
	.A2(n1262), 
	.A1(n998));
   NAND4_X1 U3495 (.ZN(n3481), 
	.A4(n3501), 
	.A3(n3500), 
	.A2(n759), 
	.A1(n3499));
   AOI221_X1 U3496 (.ZN(n3501), 
	.C2(n16847), 
	.C1(n529), 
	.B2(n16854), 
	.B1(n998), 
	.A(n3502));
   AOI21_X1 U3497 (.ZN(n3500), 
	.B2(n16833), 
	.B1(n1868), 
	.A(n3503));
   AOI211_X1 U3498 (.ZN(n3503), 
	.C2(n3504), 
	.C1(n918), 
	.B(n16845), 
	.A(FE_OFN70_n16867));
   NAND2_X1 U3499 (.ZN(n3504), 
	.A2(FE_OFN73_n16806), 
	.A1(n16825));
   INV_X1 U3500 (.ZN(n1868), 
	.A(n723));
   NAND2_X1 U3501 (.ZN(n723), 
	.A2(n16838), 
	.A1(n483));
   NAND2_X1 U3502 (.ZN(n759), 
	.A2(n16855), 
	.A1(n501));
   OAI211_X1 U3503 (.ZN(n3499), 
	.C2(n3506), 
	.C1(n3505), 
	.B(n568), 
	.A(n653));
   NOR2_X1 U3504 (.ZN(n3505), 
	.A2(n16826), 
	.A1(FE_OFN100_n1086));
   OAI221_X1 U3505 (.ZN(n3490), 
	.C2(n1580), 
	.C1(n1519), 
	.B2(n3507), 
	.B1(FE_OFN633_n16868), 
	.A(n3508));
   NOR2_X1 U3506 (.ZN(n3508), 
	.A2(n3510), 
	.A1(n3509));
   NOR3_X1 U3507 (.ZN(n3510), 
	.A3(n16824), 
	.A2(n16845), 
	.A1(FE_OFN103_n715));
   AOI222_X1 U3508 (.ZN(n3507), 
	.C2(n16836), 
	.C1(n563), 
	.B2(n16859), 
	.B1(n751), 
	.A2(FE_OFN72_n16867), 
	.A1(n760));
   INV_X1 U3509 (.ZN(n751), 
	.A(n648));
   NAND2_X1 U3510 (.ZN(n648), 
	.A2(FE_OFN82_n16856), 
	.A1(FE_OFN70_n16867));
   AOI21_X1 U3511 (.ZN(n3485), 
	.B2(n2049), 
	.B1(n16859), 
	.A(n2631));
   INV_X1 U3512 (.ZN(n2631), 
	.A(n1334));
   NAND2_X1 U3513 (.ZN(n1334), 
	.A2(n16831), 
	.A1(n16838));
   INV_X1 U3514 (.ZN(n2049), 
	.A(n3363));
   NAND2_X1 U3515 (.ZN(n3363), 
	.A2(n16870), 
	.A1(n3430));
   AND3_X1 U3516 (.ZN(n3486), 
	.A3(n17122), 
	.A2(n713), 
	.A1(n3479));
   NAND3_X1 U3517 (.ZN(n3479), 
	.A3(n3513), 
	.A2(n3512), 
	.A1(n3511));
   NOR4_X1 U3518 (.ZN(n3513), 
	.A4(n3516), 
	.A3(n784), 
	.A2(n3515), 
	.A1(n3514));
   NOR4_X1 U3519 (.ZN(n3515), 
	.A4(n755), 
	.A3(n568), 
	.A2(n556), 
	.A1(n16808));
   OAI221_X1 U3520 (.ZN(n3514), 
	.C2(n3519), 
	.C1(n3518), 
	.B2(FE_OFN106_n585), 
	.B1(n3517), 
	.A(n3520));
   NAND3_X1 U3521 (.ZN(n3520), 
	.A3(n1042), 
	.A2(n16862), 
	.A1(n909));
   AOI211_X1 U3522 (.ZN(n3519), 
	.C2(n827), 
	.C1(n1042), 
	.B(n3521), 
	.A(n16833));
   NOR3_X1 U3523 (.ZN(n3521), 
	.A3(n1023), 
	.A2(FE_OFN100_n1086), 
	.A1(n617));
   AOI211_X1 U3524 (.ZN(n3518), 
	.C2(n897), 
	.C1(n1605), 
	.B(n16828), 
	.A(n3522));
   OAI33_X1 U3525 (.ZN(n3522), 
	.B3(n16826), 
	.B2(FE_OFN98_n1104), 
	.B1(n849), 
	.A3(FE_OFN17_n16805), 
	.A2(n1519), 
	.A1(n617));
   INV_X1 U3526 (.ZN(n1605), 
	.A(n912));
   NAND2_X1 U3527 (.ZN(n912), 
	.A2(n16851), 
	.A1(n565));
   AOI22_X1 U3528 (.ZN(n3517), 
	.B2(n16824), 
	.B1(n1946), 
	.A2(n3430), 
	.A1(n812));
   INV_X1 U3529 (.ZN(n812), 
	.A(n2689));
   NAND2_X1 U3530 (.ZN(n2689), 
	.A2(n16690), 
	.A1(n16680));
   AOI222_X1 U3531 (.ZN(n3512), 
	.C2(n3525), 
	.C1(n563), 
	.B2(FE_OFN85_n16839), 
	.B1(n3524), 
	.A2(n3523), 
	.A1(n757));
   OAI211_X1 U3532 (.ZN(n3525), 
	.C2(n17096), 
	.C1(n3526), 
	.B(n3528), 
	.A(n3527));
   NAND3_X1 U3533 (.ZN(n3527), 
	.A3(n997), 
	.A2(FE_OFN87_n16848), 
	.A1(n566));
   AOI21_X1 U3534 (.ZN(n3526), 
	.B2(n16680), 
	.B1(n1034), 
	.A(n1803));
   OAI22_X1 U3535 (.ZN(n3524), 
	.B2(n16821), 
	.B1(n3529), 
	.A2(n758), 
	.A1(n917));
   AOI21_X1 U3536 (.ZN(n3529), 
	.B2(FE_OFN81_n16856), 
	.B1(n608), 
	.A(n1207));
   INV_X1 U3537 (.ZN(n1207), 
	.A(n1027));
   OAI221_X1 U3538 (.ZN(n3523), 
	.C2(n673), 
	.C1(FE_OFN70_n16867), 
	.B2(n568), 
	.B1(n16843), 
	.A(n3530));
   AOI221_X1 U3539 (.ZN(n3530), 
	.C2(n16836), 
	.C1(n3531), 
	.B2(n16826), 
	.B1(n3432), 
	.A(n1564));
   NOR2_X1 U3540 (.ZN(n3531), 
	.A2(n16828), 
	.A1(n16845));
   INV_X1 U3541 (.ZN(n3432), 
	.A(n3429));
   NAND2_X1 U3542 (.ZN(n3429), 
	.A2(FE_OFN90_n16849), 
	.A1(n16845));
   AOI222_X1 U3543 (.ZN(n3511), 
	.C2(n3532), 
	.C1(n2661), 
	.B2(n785), 
	.B1(n827), 
	.A2(n565), 
	.A1(n506));
   INV_X1 U3544 (.ZN(n785), 
	.A(n524));
   NAND2_X1 U3545 (.ZN(n524), 
	.A2(n17096), 
	.A1(n16826));
   OAI22_X1 U3546 (.ZN(U229_Z_0), 
	.B2(n2087), 
	.B1(n3533), 
	.A2(n2085), 
	.A1(n4948));
   INV_X1 U3547 (.ZN(n2087), 
	.A(n2085));
   AOI222_X1 U3548 (.ZN(n3533), 
	.C2(n84), 
	.C1(n1510), 
	.B2(n2077), 
	.B1(n86), 
	.A2(n3534), 
	.A1(n88));
   AOI22_X1 U3549 (.ZN(n1510), 
	.B2(n1783), 
	.B1(n1759), 
	.A2(n4947), 
	.A1(n2102));
   INV_X1 U3550 (.ZN(n1783), 
	.A(n3535));
   OAI221_X1 U3551 (.ZN(n3535), 
	.C2(n3477), 
	.C1(n2375), 
	.B2(n2376), 
	.B1(n3092), 
	.A(n3536));
   AOI22_X1 U3552 (.ZN(n3536), 
	.B2(n1787), 
	.B1(n2322), 
	.A2(n3538), 
	.A1(n3537));
   OAI22_X1 U3553 (.ZN(n3537), 
	.B2(n2390), 
	.B1(n1791), 
	.A2(n3539), 
	.A1(n1789));
   INV_X1 U3554 (.ZN(n2102), 
	.A(n2078));
   OAI211_X1 U3555 (.ZN(n2078), 
	.C2(n3540), 
	.C1(n94), 
	.B(n3542), 
	.A(n3541));
   AOI222_X1 U3556 (.ZN(n3542), 
	.C2(FE_OFN2_n2015), 
	.C1(n16688), 
	.B2(n3534), 
	.B1(n17008), 
	.A2(vis_apsr_o[3]), 
	.A1(n2125));
   OAI22_X1 U3557 (.ZN(n2015), 
	.B2(n3544), 
	.B1(n4950), 
	.A2(n3543), 
	.A1(n16957));
   AOI221_X1 U3558 (.ZN(n3544), 
	.C2(n3545), 
	.C1(n16824), 
	.B2(FE_OFN610_n16690), 
	.B1(n1041), 
	.A(n1095));
   OAI211_X1 U3559 (.ZN(n3545), 
	.C2(n3546), 
	.C1(n16828), 
	.B(n1023), 
	.A(n1233));
   INV_X1 U3560 (.ZN(n1041), 
	.A(n1043));
   NAND2_X1 U3561 (.ZN(n1043), 
	.A2(n16860), 
	.A1(n16851));
   OAI21_X1 U3563 (.ZN(n2243), 
	.B2(n3547), 
	.B1(n543), 
	.A(FE_OFN10_n1697));
   NOR2_X1 U3564 (.ZN(n3547), 
	.A2(n532), 
	.A1(n1218));
   NAND2_X1 U3565 (.ZN(n1218), 
	.A2(n16855), 
	.A1(FE_OFN73_n16806));
   NAND2_X2 U3567 (.ZN(n713), 
	.A2(n16831), 
	.A1(n914));
   NOR3_X1 U3569 (.ZN(n2125), 
	.A3(n2168), 
	.A2(FE_OFN15_n16671), 
	.A1(n16656));
   NAND4_X1 U3570 (.ZN(n2168), 
	.A4(FE_OFN10_n1697), 
	.A3(n1574), 
	.A2(FE_OFN633_n16868), 
	.A1(n2662));
   INV_X1 U3571 (.ZN(n2662), 
	.A(n606));
   NAND2_X2 U3572 (.ZN(n606), 
	.A2(FE_OFN82_n16856), 
	.A1(n16862));
   AOI21_X1 U3573 (.ZN(n3541), 
	.B2(n1513), 
	.B1(n3548), 
	.A(n2055));
   NAND3_X2 U3575 (.ZN(n2124), 
	.A3(n1034), 
	.A2(FE_OFN10_n1697), 
	.A1(n16828));
   NOR2_X1 U3576 (.ZN(n3548), 
	.A2(n16992), 
	.A1(U186_Z_0));
   NAND2_X2 U3578 (.ZN(n2127), 
	.A2(n2501), 
	.A1(n3549));
   AOI22_X1 U3579 (.ZN(n3540), 
	.B2(n16994), 
	.B1(n1872), 
	.A2(n2126), 
	.A1(n1513));
   INV_X1 U3582 (.ZN(n1872), 
	.A(n1513));
   OAI221_X1 U3584 (.ZN(n3550), 
	.C2(n16828), 
	.C1(n501), 
	.B2(n515), 
	.B1(n1803), 
	.A(n16845));
   INV_X1 U3585 (.ZN(n3549), 
	.A(n3551));
   OAI22_X1 U3586 (.ZN(n3551), 
	.B2(n3552), 
	.B1(n4950), 
	.A2(n2628), 
	.A1(n16957));
   AOI211_X1 U3587 (.ZN(n3552), 
	.C2(n16826), 
	.C1(n884), 
	.B(n3554), 
	.A(n3553));
   NOR3_X1 U3588 (.ZN(n3554), 
	.A3(n1519), 
	.A2(n16859), 
	.A1(n16826));
   OAI21_X1 U3589 (.ZN(n3553), 
	.B2(n818), 
	.B1(FE_OFN626_n16820), 
	.A(n3555));
   INV_X1 U3590 (.ZN(n3555), 
	.A(n3502));
   OAI21_X1 U3591 (.ZN(n3502), 
	.B2(n3556), 
	.B1(n762), 
	.A(n1541));
   NAND2_X1 U3592 (.ZN(n3556), 
	.A2(n16821), 
	.A1(n998));
   INV_X1 U3593 (.ZN(n998), 
	.A(n860));
   NAND2_X1 U3594 (.ZN(n860), 
	.A2(n16845), 
	.A1(n16825));
   NAND2_X1 U3595 (.ZN(n818), 
	.A2(n16838), 
	.A1(n914));
   NOR2_X1 U3596 (.ZN(n884), 
	.A2(n16862), 
	.A1(n532));
   INV_X1 U3597 (.ZN(n2628), 
	.A(n3543));
   OAI22_X1 U3598 (.ZN(n3543), 
	.B2(n3558), 
	.B1(n5100), 
	.A2(n795), 
	.A1(n3557));
   AOI22_X1 U3599 (.ZN(n3558), 
	.B2(n3560), 
	.B1(n16810), 
	.A2(FE_OFN15_n16671), 
	.A1(n3559));
   OAI33_X1 U3600 (.ZN(n3560), 
	.B3(n3565), 
	.B2(n16809), 
	.B1(n3564), 
	.A3(n3563), 
	.A2(n3562), 
	.A1(n3561));
   AOI221_X1 U3601 (.ZN(n3565), 
	.C2(n3566), 
	.C1(n3348), 
	.B2(n1821), 
	.B1(n3255), 
	.A(n3567));
   INV_X1 U3602 (.ZN(n3255), 
	.A(n2764));
   OAI22_X1 U3603 (.ZN(n3564), 
	.B2(n1820), 
	.B1(n3256), 
	.A2(n1900), 
	.A1(n3349));
   INV_X1 U3604 (.ZN(n3256), 
	.A(n2809));
   NOR2_X1 U3605 (.ZN(n3563), 
	.A2(n1900), 
	.A1(n3346));
   AOI221_X1 U3606 (.ZN(n3562), 
	.C2(n3566), 
	.C1(n3345), 
	.B2(n1821), 
	.B1(n3251), 
	.A(n3567));
   INV_X1 U3607 (.ZN(n3251), 
	.A(n2507));
   OAI21_X1 U3608 (.ZN(n3561), 
	.B2(n1820), 
	.B1(n3252), 
	.A(n16809));
   INV_X1 U3609 (.ZN(n3252), 
	.A(n2705));
   OAI33_X1 U3610 (.ZN(n3559), 
	.B3(n3572), 
	.B2(n16809), 
	.B1(n3571), 
	.A3(n3570), 
	.A2(n3569), 
	.A1(n3568));
   AOI221_X1 U3611 (.ZN(n3572), 
	.C2(n3566), 
	.C1(n3319), 
	.B2(n1821), 
	.B1(n3239), 
	.A(n3567));
   INV_X1 U3612 (.ZN(n3239), 
	.A(FE_OFN543_n2585));
   OAI22_X1 U3613 (.ZN(n3571), 
	.B2(n1820), 
	.B1(n3240), 
	.A2(n1900), 
	.A1(n3280));
   INV_X1 U3614 (.ZN(n3240), 
	.A(FE_OFN560_n3199));
   NOR2_X1 U3615 (.ZN(n3570), 
	.A2(n1900), 
	.A1(n3315));
   AOI221_X1 U3616 (.ZN(n3569), 
	.C2(n3566), 
	.C1(n3314), 
	.B2(n1821), 
	.B1(n3231), 
	.A(n3567));
   INV_X1 U3617 (.ZN(n3231), 
	.A(n3317));
   OAI21_X1 U3618 (.ZN(n3568), 
	.B2(n1820), 
	.B1(n3233), 
	.A(n16809));
   INV_X1 U3619 (.ZN(n3233), 
	.A(n2531));
   AOI22_X1 U3620 (.ZN(n3557), 
	.B2(n3574), 
	.B1(n16810), 
	.A2(FE_OFN15_n16671), 
	.A1(n3573));
   OAI33_X1 U3621 (.ZN(n3574), 
	.B3(n3579), 
	.B2(n16809), 
	.B1(n3578), 
	.A3(n3577), 
	.A2(n3576), 
	.A1(n3575));
   AOI221_X1 U3622 (.ZN(n3579), 
	.C2(n1821), 
	.C1(n3281), 
	.B2(n3566), 
	.B1(n3338), 
	.A(n3567));
   INV_X1 U3623 (.ZN(n3281), 
	.A(n2271));
   OAI22_X1 U3624 (.ZN(n3578), 
	.B2(n1900), 
	.B1(n3339), 
	.A2(n1820), 
	.A1(n3282));
   INV_X1 U3625 (.ZN(n3282), 
	.A(n2452));
   NOR2_X1 U3626 (.ZN(n3577), 
	.A2(n1820), 
	.A1(n3398));
   INV_X1 U3627 (.ZN(n3398), 
	.A(n2297));
   AOI221_X1 U3628 (.ZN(n3576), 
	.C2(n1821), 
	.C1(n2183), 
	.B2(n3566), 
	.B1(n3278), 
	.A(n3567));
   INV_X1 U3629 (.ZN(n2183), 
	.A(n3274));
   OAI21_X1 U3630 (.ZN(n3575), 
	.B2(n1900), 
	.B1(n3341), 
	.A(n16809));
   OAI33_X1 U3631 (.ZN(n3573), 
	.B3(n3584), 
	.B2(n16809), 
	.B1(n3583), 
	.A3(n3582), 
	.A2(n3581), 
	.A1(n3580));
   AOI221_X1 U3632 (.ZN(n3584), 
	.C2(n3566), 
	.C1(n3328), 
	.B2(n1821), 
	.B1(n3261), 
	.A(n3567));
   INV_X1 U3633 (.ZN(n3261), 
	.A(n3041));
   OAI22_X1 U3634 (.ZN(n3583), 
	.B2(n1820), 
	.B1(n3262), 
	.A2(n1900), 
	.A1(n3329));
   INV_X1 U3635 (.ZN(n3262), 
	.A(n3155));
   NOR2_X1 U3636 (.ZN(n3582), 
	.A2(n1900), 
	.A1(n3333));
   INV_X1 U3638 (.ZN(n3333), 
	.A(n3022));
   AOI221_X1 U3639 (.ZN(n3581), 
	.C2(n3566), 
	.C1(n3332), 
	.B2(n1821), 
	.B1(n3264), 
	.A(n3567));
   AND2_X1 U3640 (.ZN(n3567), 
	.A2(n3566), 
	.A1(n1821));
   INV_X1 U3643 (.ZN(n3264), 
	.A(n2856));
   OAI21_X1 U3644 (.ZN(n3580), 
	.B2(n1820), 
	.B1(n3265), 
	.A(n16809));
   NAND4_X1 U3647 (.ZN(n1513), 
	.A4(n3588), 
	.A3(n3587), 
	.A2(n3586), 
	.A1(n3585));
   AOI222_X1 U3648 (.ZN(n3588), 
	.C2(vis_msp_o[29]), 
	.C1(n16975), 
	.B2(vis_psp_o[29]), 
	.B1(n16969), 
	.A2(vis_r12_o[31]), 
	.A1(FE_OFN109_n16964));
   NAND3_X2 U3653 (.ZN(n2182), 
	.A3(n3593), 
	.A2(n5036), 
	.A1(n4978));
   AOI222_X1 U3654 (.ZN(n3587), 
	.C2(vis_r14_o[31]), 
	.C1(n16984), 
	.B2(vis_r11_o[31]), 
	.B1(n16987), 
	.A2(vis_r10_o[31]), 
	.A1(n16961));
   NOR2_X1 U3657 (.ZN(n3593), 
	.A2(n3597), 
	.A1(n2184));
   NAND3_X2 U3661 (.ZN(n2191), 
	.A3(n3598), 
	.A2(n3480), 
	.A1(n4978));
   AOI222_X1 U3662 (.ZN(n3586), 
	.C2(vis_r9_o[31]), 
	.C1(n16979), 
	.B2(vis_r8_o[31]), 
	.B1(n16960), 
	.A2(n3400), 
	.A1(n16970));
   NAND2_X2 U3664 (.ZN(n2637), 
	.A2(n3592), 
	.A1(n3598));
   NAND3_X2 U3667 (.ZN(n2190), 
	.A3(n3598), 
	.A2(n5036), 
	.A1(n4978));
   NOR3_X2 U3668 (.ZN(n3598), 
	.A3(n2184), 
	.A2(n4959), 
	.A1(n3492));
   NAND2_X2 U3670 (.ZN(n2184), 
	.A2(n3601), 
	.A1(n16957));
   AOI22_X1 U3672 (.ZN(n3585), 
	.B2(n874), 
	.B1(n16956), 
	.A2(n867), 
	.A1(n16976));
   NOR4_X2 U3676 (.ZN(n3601), 
	.A4(n3604), 
	.A3(n3603), 
	.A2(n3602), 
	.A1(n727));
   OAI221_X2 U3677 (.ZN(n3604), 
	.C2(FE_OFN100_n1086), 
	.C1(FE_OFN73_n16806), 
	.B2(n3221), 
	.B1(n989), 
	.A(n3605));
   OAI21_X2 U3678 (.ZN(n3605), 
	.B2(n527), 
	.B1(n991), 
	.A(n16845));
   INV_X4 U3679 (.ZN(n3221), 
	.A(n1300));
   NOR2_X2 U3680 (.ZN(n1300), 
	.A2(FE_OFN87_n16848), 
	.A1(FE_OFN84_n16839));
   OAI33_X1 U3681 (.ZN(n3603), 
	.B3(n5036), 
	.B2(n4978), 
	.B1(n3597), 
	.A3(n604), 
	.A2(n16871), 
	.A1(FE_OFN103_n715));
   NAND2_X1 U3682 (.ZN(n3597), 
	.A2(n3495), 
	.A1(n3492));
   NOR3_X1 U3683 (.ZN(n3602), 
	.A3(n16826), 
	.A2(n16836), 
	.A1(n994));
   INV_X4 U3684 (.ZN(n994), 
	.A(n1946));
   NOR2_X2 U3685 (.ZN(n1946), 
	.A2(FE_OFN87_n16848), 
	.A1(n1234));
   INV_X4 U3686 (.ZN(n727), 
	.A(n891));
   OAI21_X2 U3687 (.ZN(n2222), 
	.B2(n1177), 
	.B1(n16821), 
	.A(n3606));
   NAND3_X1 U3688 (.ZN(n3606), 
	.A3(n1034), 
	.A2(n16871), 
	.A1(n3430));
   NAND4_X2 U3689 (.ZN(n1177), 
	.A4(FE_OFN81_n16856), 
	.A3(n991), 
	.A2(n1805), 
	.A1(n597));
   INV_X1 U3690 (.ZN(n94), 
	.A(U186_Z_0));
   INV_X1 U3691 (.ZN(n2077), 
	.A(FE_PHN711_n28));
   AOI221_X1 U3692 (.ZN(n28), 
	.C2(n2072), 
	.C1(FE_PSN5239_n2057), 
	.B2(n2067), 
	.B1(n2061), 
	.A(n3607));
   INV_X2 U3693 (.ZN(n3607), 
	.A(n3608));
   AOI221_X1 U3694 (.ZN(n3608), 
	.C2(n2058), 
	.C1(n2074), 
	.B2(n2062), 
	.B1(n2069), 
	.A(n2076));
   NAND4_X2 U3697 (.ZN(n3209), 
	.A4(n3611), 
	.A3(n3610), 
	.A2(n3092), 
	.A1(1'b1));
   AOI222_X1 U3698 (.ZN(n3611), 
	.C2(FE_OFN514_n2062), 
	.C1(n3614), 
	.B2(n1564), 
	.B1(n3613), 
	.A2(n3612), 
	.A1(n3532));
   OAI21_X1 U3699 (.ZN(n3614), 
	.B2(FE_OFN632_n16859), 
	.B1(n3615), 
	.A(FE_OFN483_n1233));
   AOI21_X1 U3700 (.ZN(n3615), 
	.B2(n5102), 
	.B1(n5227), 
	.A(n16842));
   NOR2_X1 U3701 (.ZN(n3613), 
	.A2(FE_OFN84_n16839), 
	.A1(n3616));
   OAI21_X1 U3702 (.ZN(n3612), 
	.B2(n3616), 
	.B1(n5227), 
	.A(n3617));
   NAND3_X1 U3703 (.ZN(n3617), 
	.A3(n5227), 
	.A2(n3223), 
	.A1(n2061));
   AOI22_X1 U3704 (.ZN(n3616), 
	.B2(n5102), 
	.B1(FE_OFN512_n2058), 
	.A2(FE_OFN511_n2057), 
	.A1(n3223));
   INV_X1 U3706 (.ZN(n3532), 
	.A(n917));
   NAND2_X1 U3707 (.ZN(n917), 
	.A2(n16862), 
	.A1(n16845));
   NAND4_X1 U3708 (.ZN(n3610), 
	.A4(FE_OFN72_n16867), 
	.A3(FE_OFN632_n16859), 
	.A2(n16847), 
	.A1(FE_OFN512_n2058));
   INV_X1 U3709 (.ZN(n3609), 
	.A(n3473));
   OAI211_X1 U3710 (.ZN(n3473), 
	.C2(FE_OFN98_n1104), 
	.C1(n16862), 
	.B(n3618), 
	.A(n3215));
   NOR2_X1 U3711 (.ZN(n3618), 
	.A2(n3620), 
	.A1(1'b0));
   NOR3_X1 U3712 (.ZN(n3620), 
	.A3(n16854), 
	.A2(n16868), 
	.A1(FE_OFN429_n673));
   OR3_X1 U3715 (.ZN(n2376), 
	.A3(n2323), 
	.A2(n2322), 
	.A1(n2359));
   AOI21_X1 U3716 (.ZN(n2323), 
	.B2(n2390), 
	.B1(n3539), 
	.A(n2389));
   INV_X1 U3717 (.ZN(n2359), 
	.A(n3477));
   NAND3_X2 U3718 (.ZN(n2058), 
	.A3(n3623), 
	.A2(n3622), 
	.A1(n3621));
   AOI221_X1 U3719 (.ZN(n3623), 
	.C2(n3624), 
	.C1(n2922), 
	.B2(n2879), 
	.B1(hrdata_i[15]), 
	.A(n3625));
   OAI22_X1 U3720 (.ZN(n3625), 
	.B2(n16685), 
	.B1(FE_PHN2429_n5505), 
	.A2(n282), 
	.A1(n2981));
   INV_X1 U3722 (.ZN(n3624), 
	.A(n1791));
   OAI22_X1 U3723 (.ZN(n1791), 
	.B2(n2354), 
	.B1(n2337), 
	.A2(n2384), 
	.A1(n16788));
   OAI221_X1 U3724 (.ZN(n2354), 
	.C2(n16951), 
	.C1(n3348), 
	.B2(n16948), 
	.B1(n3346), 
	.A(n3626));
   AOI22_X1 U3725 (.ZN(n3626), 
	.B2(n2705), 
	.B1(n16942), 
	.A2(n2764), 
	.A1(n16945));
   NAND3_X1 U3726 (.ZN(n2705), 
	.A3(n3629), 
	.A2(n3628), 
	.A1(n3627));
   AOI221_X1 U3727 (.ZN(n3629), 
	.C2(vis_r0_o[22]), 
	.C1(FE_OFN644_n16936), 
	.B2(vis_r2_o[22]), 
	.B1(FE_OFN645_n16939), 
	.A(n3634));
   OAI22_X1 U3728 (.ZN(n3634), 
	.B2(n16931), 
	.B1(n5436), 
	.A2(n16934), 
	.A1(n5050));
   AOI22_X1 U3730 (.ZN(n3628), 
	.B2(vis_r4_o[22]), 
	.B1(n16924), 
	.A2(vis_r5_o[22]), 
	.A1(n16927));
   AOI22_X1 U3731 (.ZN(n3627), 
	.B2(vis_r1_o[22]), 
	.B1(n16918), 
	.A2(vis_r6_o[22]), 
	.A1(n16921));
   NAND3_X1 U3734 (.ZN(n2764), 
	.A3(n3647), 
	.A2(n3646), 
	.A1(n3645));
   AOI221_X1 U3735 (.ZN(n3647), 
	.C2(vis_r0_o[20]), 
	.C1(FE_OFN644_n16936), 
	.B2(vis_r2_o[20]), 
	.B1(FE_OFN645_n16939), 
	.A(n3650));
   OAI22_X1 U3736 (.ZN(n3650), 
	.B2(n16931), 
	.B1(n5605), 
	.A2(n16934), 
	.A1(n5613));
   AOI22_X1 U3738 (.ZN(n3646), 
	.B2(vis_r4_o[20]), 
	.B1(n16924), 
	.A2(vis_r5_o[20]), 
	.A1(n16927));
   AOI22_X1 U3739 (.ZN(n3645), 
	.B2(vis_r1_o[20]), 
	.B1(n16918), 
	.A2(vis_r6_o[20]), 
	.A1(n16921));
   INV_X1 U3742 (.ZN(n3348), 
	.A(n2787));
   NAND3_X1 U3743 (.ZN(n2787), 
	.A3(n3657), 
	.A2(n3656), 
	.A1(n3655));
   AOI221_X1 U3744 (.ZN(n3657), 
	.C2(vis_r0_o[19]), 
	.C1(FE_OFN644_n16936), 
	.B2(vis_r2_o[19]), 
	.B1(FE_OFN645_n16939), 
	.A(n3660));
   OAI22_X1 U3745 (.ZN(n3660), 
	.B2(n16931), 
	.B1(n5438), 
	.A2(n16934), 
	.A1(n5090));
   AOI22_X1 U3747 (.ZN(n3656), 
	.B2(vis_r4_o[19]), 
	.B1(n16924), 
	.A2(vis_r5_o[19]), 
	.A1(n16927));
   AOI22_X1 U3748 (.ZN(n3655), 
	.B2(vis_r1_o[19]), 
	.B1(n16918), 
	.A2(vis_r6_o[19]), 
	.A1(n16921));
   INV_X1 U3751 (.ZN(n3346), 
	.A(n2738));
   NAND3_X1 U3752 (.ZN(n2738), 
	.A3(n3667), 
	.A2(n3666), 
	.A1(n3665));
   AOI221_X1 U3753 (.ZN(n3667), 
	.C2(vis_r0_o[21]), 
	.C1(FE_OFN644_n16936), 
	.B2(vis_r2_o[21]), 
	.B1(FE_OFN645_n16939), 
	.A(n3670));
   OAI22_X1 U3754 (.ZN(n3670), 
	.B2(n16931), 
	.B1(n5437), 
	.A2(n16934), 
	.A1(n5117));
   AOI22_X1 U3756 (.ZN(n3666), 
	.B2(vis_r4_o[21]), 
	.B1(n16924), 
	.A2(vis_r5_o[21]), 
	.A1(n16927));
   AOI22_X1 U3757 (.ZN(n3665), 
	.B2(vis_r1_o[21]), 
	.B1(n16918), 
	.A2(vis_r6_o[21]), 
	.A1(n16921));
   OAI221_X1 U3760 (.ZN(n2384), 
	.C2(n16951), 
	.C1(n3332), 
	.B2(n16948), 
	.B1(n3349), 
	.A(n3675));
   AOI22_X1 U3761 (.ZN(n3675), 
	.B2(n2809), 
	.B1(n16942), 
	.A2(n2856), 
	.A1(n16945));
   NAND3_X1 U3762 (.ZN(n2809), 
	.A3(n3678), 
	.A2(n3677), 
	.A1(n3676));
   AOI221_X1 U3763 (.ZN(n3678), 
	.C2(vis_r0_o[18]), 
	.C1(FE_OFN644_n16936), 
	.B2(vis_r2_o[18]), 
	.B1(FE_OFN645_n16939), 
	.A(n3681));
   OAI22_X1 U3764 (.ZN(n3681), 
	.B2(n16931), 
	.B1(n5439), 
	.A2(n16934), 
	.A1(n5064));
   AOI22_X1 U3766 (.ZN(n3677), 
	.B2(vis_r4_o[18]), 
	.B1(n16924), 
	.A2(vis_r5_o[18]), 
	.A1(n16927));
   AOI22_X1 U3767 (.ZN(n3676), 
	.B2(vis_r1_o[18]), 
	.B1(n16918), 
	.A2(vis_r6_o[18]), 
	.A1(n16921));
   NAND3_X1 U3770 (.ZN(n2856), 
	.A3(n3688), 
	.A2(n3687), 
	.A1(n3686));
   AOI221_X1 U3771 (.ZN(n3688), 
	.C2(vis_r0_o[16]), 
	.C1(FE_OFN644_n16936), 
	.B2(vis_r2_o[16]), 
	.B1(FE_OFN645_n16939), 
	.A(n3691));
   OAI22_X1 U3772 (.ZN(n3691), 
	.B2(n16931), 
	.B1(n5441), 
	.A2(n16934), 
	.A1(n5071));
   AOI22_X1 U3774 (.ZN(n3687), 
	.B2(vis_r4_o[16]), 
	.B1(n16924), 
	.A2(vis_r5_o[16]), 
	.A1(n16927));
   AOI22_X1 U3775 (.ZN(n3686), 
	.B2(vis_r1_o[16]), 
	.B1(n16918), 
	.A2(vis_r6_o[16]), 
	.A1(n16921));
   INV_X1 U3778 (.ZN(n3332), 
	.A(n3267));
   NAND3_X1 U3779 (.ZN(n3267), 
	.A3(n3698), 
	.A2(n3697), 
	.A1(n3696));
   AOI221_X1 U3780 (.ZN(n3698), 
	.C2(vis_r0_o[15]), 
	.C1(FE_OFN644_n16936), 
	.B2(vis_r2_o[15]), 
	.B1(FE_OFN645_n16939), 
	.A(n3701));
   OAI22_X1 U3781 (.ZN(n3701), 
	.B2(n16931), 
	.B1(n5449), 
	.A2(n16934), 
	.A1(n5110));
   AOI22_X1 U3783 (.ZN(n3697), 
	.B2(vis_r4_o[15]), 
	.B1(n16924), 
	.A2(vis_r5_o[15]), 
	.A1(n16927));
   AOI22_X1 U3784 (.ZN(n3696), 
	.B2(vis_r1_o[15]), 
	.B1(n16918), 
	.A2(vis_r6_o[15]), 
	.A1(n16921));
   INV_X1 U3787 (.ZN(n3349), 
	.A(n2833));
   NAND3_X1 U3788 (.ZN(n2833), 
	.A3(n3708), 
	.A2(n3707), 
	.A1(n3706));
   AOI221_X1 U3789 (.ZN(n3708), 
	.C2(vis_r0_o[17]), 
	.C1(FE_OFN644_n16936), 
	.B2(vis_r2_o[17]), 
	.B1(FE_OFN645_n16939), 
	.A(n3711));
   OAI22_X1 U3790 (.ZN(n3711), 
	.B2(n16931), 
	.B1(n5440), 
	.A2(n16934), 
	.A1(n5085));
   AOI22_X1 U3792 (.ZN(n3707), 
	.B2(vis_r4_o[17]), 
	.B1(n16924), 
	.A2(vis_r5_o[17]), 
	.A1(n16927));
   AOI22_X1 U3793 (.ZN(n3706), 
	.B2(vis_r1_o[17]), 
	.B1(n16918), 
	.A2(vis_r6_o[17]), 
	.A1(n16921));
   AOI221_X1 U3796 (.ZN(n3622), 
	.C2(n3716), 
	.C1(n2882), 
	.B2(n416), 
	.B1(n2895), 
	.A(n2897));
   INV_X1 U3797 (.ZN(n2897), 
	.A(n3247));
   NAND4_X1 U3798 (.ZN(n3247), 
	.A4(n5017), 
	.A3(n2882), 
	.A2(n3717), 
	.A1(FE_OFN573_n4905));
   OAI221_X1 U3799 (.ZN(n3716), 
	.C2(n2899), 
	.C1(n5156), 
	.B2(n2898), 
	.B1(n5150), 
	.A(n3718));
   AOI22_X1 U3800 (.ZN(n3718), 
	.B2(n3720), 
	.B1(n1893), 
	.A2(n3719), 
	.A1(n1897));
   INV_X1 U3801 (.ZN(n416), 
	.A(n424));
   NAND2_X1 U3802 (.ZN(n424), 
	.A2(n3721), 
	.A1(n2905));
   NAND3_X1 U3803 (.ZN(n3721), 
	.A3(n2907), 
	.A2(n1372), 
	.A1(n2908));
   NOR3_X1 U3804 (.ZN(n2905), 
	.A3(n1066), 
	.A2(n1067), 
	.A1(n3066));
   NOR3_X1 U3805 (.ZN(n1067), 
	.A3(n1370), 
	.A2(n2907), 
	.A1(n3722));
   INV_X1 U3806 (.ZN(n1370), 
	.A(n1372));
   OAI21_X1 U3807 (.ZN(n1372), 
	.B2(n209), 
	.B1(n3723), 
	.A(n3724));
   OAI221_X1 U3808 (.ZN(n3724), 
	.C2(n3722), 
	.C1(n2907), 
	.B2(n1371), 
	.B1(n3725), 
	.A(n3726));
   OAI21_X1 U3809 (.ZN(n3726), 
	.B2(n3728), 
	.B1(n3727), 
	.A(n1368));
   OAI22_X1 U3810 (.ZN(n1368), 
	.B2(n3730), 
	.B1(n5098), 
	.A2(n3729), 
	.A1(n3722));
   INV_X1 U3811 (.ZN(n3728), 
	.A(n3725));
   INV_X1 U3812 (.ZN(n1371), 
	.A(n3727));
   AOI22_X1 U3813 (.ZN(n3727), 
	.B2(n3723), 
	.B1(n3732), 
	.A2(n2903), 
	.A1(n3731));
   NOR2_X1 U3814 (.ZN(n3725), 
	.A2(n1369), 
	.A1(n3733));
   OAI22_X1 U3815 (.ZN(n1369), 
	.B2(n3730), 
	.B1(n5097), 
	.A2(n3722), 
	.A1(n3734));
   INV_X1 U3816 (.ZN(n3733), 
	.A(n1373));
   AOI22_X1 U3817 (.ZN(n1373), 
	.B2(n3723), 
	.B1(n5503), 
	.A2(n4826), 
	.A1(n2903));
   INV_X1 U3818 (.ZN(n3723), 
	.A(n2903));
   OAI21_X1 U3819 (.ZN(n2903), 
	.B2(n3735), 
	.B1(n4802), 
	.A(n1053));
   AOI22_X1 U3820 (.ZN(n3735), 
	.B2(n3732), 
	.B1(n4961), 
	.A2(n4826), 
	.A1(n3736));
   AOI21_X1 U3821 (.ZN(n3736), 
	.B2(n3731), 
	.B1(n5504), 
	.A(n5503));
   AND2_X1 U3822 (.ZN(n2907), 
	.A2(n3737), 
	.A1(n3730));
   INV_X1 U3823 (.ZN(n3722), 
	.A(n3730));
   OAI21_X1 U3824 (.ZN(n3730), 
	.B2(n3739), 
	.B1(n3738), 
	.A(n203));
   OAI21_X1 U3826 (.ZN(n3739), 
	.B2(n3740), 
	.B1(n3729), 
	.A(n3737));
   NAND3_X1 U3827 (.ZN(n3737), 
	.A3(n3741), 
	.A2(n2909), 
	.A1(n2911));
   AOI22_X1 U3828 (.ZN(n3738), 
	.B2(n2929), 
	.B1(n3734), 
	.A2(n3740), 
	.A1(n3729));
   AOI22_X1 U3829 (.ZN(n3734), 
	.B2(n2911), 
	.B1(n3743), 
	.A2(n2908), 
	.A1(n3742));
   OAI22_X1 U3830 (.ZN(n3729), 
	.B2(n2911), 
	.B1(n3745), 
	.A2(n3744), 
	.A1(n2908));
   INV_X1 U3831 (.ZN(n2908), 
	.A(n2911));
   OAI21_X1 U3832 (.ZN(n2911), 
	.B2(n2997), 
	.B1(n3746), 
	.A(n3747));
   OAI221_X1 U3833 (.ZN(n3747), 
	.C2(n3749), 
	.C1(n2993), 
	.B2(n3745), 
	.B1(n3748), 
	.A(n3750));
   OAI21_X1 U3834 (.ZN(n3750), 
	.B2(n3752), 
	.B1(n3751), 
	.A(n3744));
   OAI22_X1 U3835 (.ZN(n3744), 
	.B2(n2909), 
	.B1(n3754), 
	.A2(n3753), 
	.A1(n2993));
   INV_X1 U3836 (.ZN(n3752), 
	.A(n3748));
   INV_X1 U3837 (.ZN(n3751), 
	.A(n3745));
   OAI22_X1 U3838 (.ZN(n3745), 
	.B2(n3756), 
	.B1(n3073), 
	.A2(n2910), 
	.A1(n3755));
   NOR2_X1 U3839 (.ZN(n3748), 
	.A2(n3743), 
	.A1(n3757));
   OAI22_X1 U3840 (.ZN(n3743), 
	.B2(n2993), 
	.B1(n3759), 
	.A2(n2909), 
	.A1(n3758));
   INV_X1 U3841 (.ZN(n2993), 
	.A(n2909));
   NAND3_X1 U3843 (.ZN(n3763), 
	.A3(n3765), 
	.A2(n3759), 
	.A1(n3764));
   AOI21_X1 U3844 (.ZN(n3765), 
	.B2(n3754), 
	.B1(n3766), 
	.A(n3741));
   INV_X1 U3845 (.ZN(n3741), 
	.A(n3749));
   INV_X1 U3846 (.ZN(n3766), 
	.A(n3753));
   AOI22_X1 U3847 (.ZN(n3759), 
	.B2(n3086), 
	.B1(n3768), 
	.A2(n3767), 
	.A1(n2995));
   INV_X1 U3848 (.ZN(n3764), 
	.A(n3758));
   INV_X1 U3849 (.ZN(n3761), 
	.A(n2994));
   NAND2_X1 U3850 (.ZN(n3760), 
	.A2(n3753), 
	.A1(n3749));
   OAI22_X1 U3851 (.ZN(n3753), 
	.B2(n2995), 
	.B1(n3770), 
	.A2(n3769), 
	.A1(n3086));
   INV_X1 U3852 (.ZN(n3086), 
	.A(n2995));
   NAND2_X1 U3853 (.ZN(n3749), 
	.A2(n2995), 
	.A1(n3771));
   OAI21_X1 U3854 (.ZN(n2995), 
	.B2(n3772), 
	.B1(n3771), 
	.A(n3774));
   OAI21_X1 U3855 (.ZN(n3774), 
	.B2(n3775), 
	.B1(n244), 
	.A(n3087));
   AOI22_X1 U3856 (.ZN(n3772), 
	.B2(n3768), 
	.B1(n3777), 
	.A2(n3770), 
	.A1(n3776));
   AOI22_X1 U3857 (.ZN(n3768), 
	.B2(n3778), 
	.B1(n1885), 
	.A2(n5151), 
	.A1(n3087));
   AOI21_X1 U3858 (.ZN(n3777), 
	.B2(n3769), 
	.B1(n3779), 
	.A(n3767));
   AOI22_X1 U3859 (.ZN(n3767), 
	.B2(n5152), 
	.B1(n3780), 
	.A2(n5154), 
	.A1(n3088));
   INV_X1 U3860 (.ZN(n3779), 
	.A(n3770));
   OAI22_X1 U3861 (.ZN(n3770), 
	.B2(n3087), 
	.B1(n5521), 
	.A2(n3778), 
	.A1(n5150));
   INV_X1 U3862 (.ZN(n3087), 
	.A(n3778));
   NOR3_X1 U3863 (.ZN(n3778), 
	.A3(n3781), 
	.A2(n4749), 
	.A1(n4795));
   AOI211_X1 U3864 (.ZN(n3781), 
	.C2(n3783), 
	.C1(n3782), 
	.B(n3775), 
	.A(n244));
   NAND2_X1 U3866 (.ZN(n3783), 
	.A2(n5150), 
	.A1(n3784));
   OAI211_X1 U3867 (.ZN(n3782), 
	.C2(n5150), 
	.C1(n3784), 
	.B(n4753), 
	.A(n5151));
   INV_X1 U3868 (.ZN(n3776), 
	.A(n3769));
   OAI22_X1 U3869 (.ZN(n3769), 
	.B2(n3088), 
	.B1(n5153), 
	.A2(n3780), 
	.A1(n5155));
   AOI21_X1 U3870 (.ZN(n3771), 
	.B2(n3786), 
	.B1(n3785), 
	.A(n3780));
   INV_X1 U3871 (.ZN(n3780), 
	.A(n3088));
   OAI211_X1 U3872 (.ZN(n3088), 
	.C2(n3788), 
	.C1(n3787), 
	.B(n2914), 
	.A(n2916));
   NAND2_X1 U3875 (.ZN(n3788), 
	.A2(n3786), 
	.A1(n3785));
   AOI22_X1 U3876 (.ZN(n3787), 
	.B2(n3790), 
	.B1(n5155), 
	.A2(n5154), 
	.A1(n3789));
   AOI21_X1 U3877 (.ZN(n3789), 
	.B2(n3791), 
	.B1(n5153), 
	.A(n5152));
   OAI222_X1 U3878 (.ZN(n3754), 
	.C2(n2994), 
	.C1(n3795), 
	.B2(n3794), 
	.B1(n3793), 
	.A2(n3085), 
	.A1(n3792));
   OAI221_X1 U3879 (.ZN(n3758), 
	.C2(n2994), 
	.C1(n3796), 
	.B2(n3085), 
	.B1(n2932), 
	.A(n3797));
   NAND3_X1 U3880 (.ZN(n3797), 
	.A3(n5158), 
	.A2(n2994), 
	.A1(n3798));
   NAND2_X1 U3881 (.ZN(n3085), 
	.A2(n3794), 
	.A1(n2994));
   NAND3_X1 U3882 (.ZN(n2994), 
	.A3(n3801), 
	.A2(n3800), 
	.A1(n3799));
   OAI21_X1 U3883 (.ZN(n3801), 
	.B2(n5011), 
	.B1(n5578), 
	.A(n3802));
   NAND3_X1 U3884 (.ZN(n3800), 
	.A3(n3803), 
	.A2(n3795), 
	.A1(n3762));
   NAND2_X1 U3885 (.ZN(n3762), 
	.A2(n3804), 
	.A1(n3794));
   OAI21_X1 U3886 (.ZN(n3799), 
	.B2(n3795), 
	.B1(n3803), 
	.A(n3805));
   OAI22_X1 U3887 (.ZN(n3805), 
	.B2(n3804), 
	.B1(n3792), 
	.A2(n3794), 
	.A1(n3793));
   INV_X1 U3888 (.ZN(n3804), 
	.A(n3806));
   OAI22_X1 U3889 (.ZN(n3795), 
	.B2(n3802), 
	.B1(n5522), 
	.A2(n3084), 
	.A1(n5156));
   INV_X1 U3890 (.ZN(n3803), 
	.A(n3807));
   OAI221_X1 U3891 (.ZN(n3807), 
	.C2(n3798), 
	.C1(n5160), 
	.B2(n3794), 
	.B1(n5158), 
	.A(n3796));
   AOI22_X1 U3892 (.ZN(n3796), 
	.B2(n5518), 
	.B1(n3084), 
	.A2(n5157), 
	.A1(n3802));
   INV_X1 U3893 (.ZN(n3802), 
	.A(n3084));
   AOI211_X1 U3894 (.ZN(n3084), 
	.C2(n3809), 
	.C1(n3808), 
	.B(n4747), 
	.A(n4796));
   NOR2_X1 U3895 (.ZN(n3809), 
	.A2(n5011), 
	.A1(n5578));
   INV_X1 U3896 (.ZN(n3808), 
	.A(n3810));
   AOI22_X1 U3897 (.ZN(n3810), 
	.B2(n3812), 
	.B1(n5156), 
	.A2(n5157), 
	.A1(n3811));
   AOI21_X1 U3898 (.ZN(n3811), 
	.B2(n3813), 
	.B1(n5522), 
	.A(n5518));
   INV_X1 U3899 (.ZN(n3794), 
	.A(n3798));
   AOI211_X1 U3900 (.ZN(n3798), 
	.C2(n3806), 
	.C1(n3814), 
	.B(n4748), 
	.A(n5537));
   NOR2_X1 U3901 (.ZN(n3806), 
	.A2(n5572), 
	.A1(n5570));
   OAI22_X1 U3902 (.ZN(n3814), 
	.B2(n5159), 
	.B1(n3792), 
	.A2(n2932), 
	.A1(n3815));
   OAI21_X1 U3903 (.ZN(n3815), 
	.B2(n5161), 
	.B1(n3793), 
	.A(n2888));
   INV_X1 U3905 (.ZN(n3757), 
	.A(n3742));
   AOI22_X1 U3906 (.ZN(n3742), 
	.B2(n3817), 
	.B1(n2910), 
	.A2(n3073), 
	.A1(n3816));
   INV_X1 U3907 (.ZN(n3073), 
	.A(n2910));
   NAND2_X1 U3908 (.ZN(n2997), 
	.A2(n2910), 
	.A1(n3076));
   OAI21_X1 U3909 (.ZN(n2910), 
	.B2(n3818), 
	.B1(n2996), 
	.A(n3819));
   OAI221_X1 U3910 (.ZN(n3819), 
	.C2(n3746), 
	.C1(n3821), 
	.B2(n3756), 
	.B1(n3820), 
	.A(n3822));
   OAI22_X1 U3911 (.ZN(n3822), 
	.B2(n3816), 
	.B1(n3824), 
	.A2(n3755), 
	.A1(n3823));
   OAI221_X1 U3912 (.ZN(n3816), 
	.C2(n3079), 
	.C1(n3825), 
	.B2(n3080), 
	.B1(n2933), 
	.A(n3826));
   NAND3_X1 U3913 (.ZN(n3826), 
	.A3(n3827), 
	.A2(n1896), 
	.A1(n3079));
   INV_X1 U3914 (.ZN(n3825), 
	.A(n3828));
   INV_X1 U3915 (.ZN(n3824), 
	.A(n3817));
   OAI22_X1 U3916 (.ZN(n3817), 
	.B2(n3076), 
	.B1(n3830), 
	.A2(n3821), 
	.A1(n3829));
   INV_X1 U3917 (.ZN(n3823), 
	.A(n3756));
   OAI22_X1 U3918 (.ZN(n3756), 
	.B2(n3076), 
	.B1(n3832), 
	.A2(n3821), 
	.A1(n3831));
   INV_X1 U3919 (.ZN(n3821), 
	.A(n3076));
   INV_X1 U3920 (.ZN(n3820), 
	.A(n3755));
   OAI222_X1 U3921 (.ZN(n3755), 
	.C2(n3079), 
	.C1(n3836), 
	.B2(n3835), 
	.B1(n3834), 
	.A2(n3080), 
	.A1(n3833));
   NAND2_X1 U3922 (.ZN(n3080), 
	.A2(n3835), 
	.A1(n3079));
   INV_X1 U3923 (.ZN(n2996), 
	.A(n3079));
   NAND3_X1 U3924 (.ZN(n3079), 
	.A3(n3839), 
	.A2(n3838), 
	.A1(n3837));
   OAI21_X1 U3925 (.ZN(n3839), 
	.B2(n5534), 
	.B1(n5535), 
	.A(n3840));
   NAND3_X1 U3926 (.ZN(n3838), 
	.A3(n3841), 
	.A2(n3836), 
	.A1(n3818));
   NAND2_X1 U3927 (.ZN(n3818), 
	.A2(n3835), 
	.A1(n3842));
   OAI21_X1 U3928 (.ZN(n3837), 
	.B2(n3836), 
	.B1(n3841), 
	.A(n3843));
   OAI22_X1 U3929 (.ZN(n3843), 
	.B2(n3842), 
	.B1(n3833), 
	.A2(n3835), 
	.A1(n3834));
   OAI22_X1 U3930 (.ZN(n3836), 
	.B2(n3840), 
	.B1(n5549), 
	.A2(n3078), 
	.A1(n5547));
   AOI221_X1 U3931 (.ZN(n3841), 
	.C2(n3835), 
	.C1(n2933), 
	.B2(n3827), 
	.B1(n4752), 
	.A(n3828));
   OAI22_X1 U3932 (.ZN(n3828), 
	.B2(n2951), 
	.B1(n3840), 
	.A2(n2901), 
	.A1(n3078));
   INV_X1 U3933 (.ZN(n3840), 
	.A(n3078));
   AOI211_X1 U3934 (.ZN(n3078), 
	.C2(n3845), 
	.C1(n3844), 
	.B(n5005), 
	.A(n5540));
   NOR2_X1 U3935 (.ZN(n3845), 
	.A2(n5534), 
	.A1(n5535));
   OAI22_X1 U3936 (.ZN(n3844), 
	.B2(n5549), 
	.B1(n3719), 
	.A2(n2901), 
	.A1(n3846));
   OAI21_X1 U3939 (.ZN(n3846), 
	.B2(n5547), 
	.B1(n3847), 
	.A(n2951));
   INV_X1 U3941 (.ZN(n3827), 
	.A(n3835));
   OAI211_X1 U3942 (.ZN(n3835), 
	.C2(n3842), 
	.C1(n3848), 
	.B(n217), 
	.A(n3238));
   NAND2_X1 U3944 (.ZN(n3842), 
	.A2(n3107), 
	.A1(n220));
   AOI22_X1 U3947 (.ZN(n3848), 
	.B2(n3834), 
	.B1(n5553), 
	.A2(n5552), 
	.A1(n3849));
   AOI21_X1 U3949 (.ZN(n3849), 
	.B2(n3833), 
	.B1(n5551), 
	.A(n1896));
   OAI21_X1 U3951 (.ZN(n3076), 
	.B2(n3851), 
	.B1(n3850), 
	.A(n3852));
   OAI21_X1 U3952 (.ZN(n3852), 
	.B2(n3010), 
	.B1(n5533), 
	.A(n3853));
   AOI22_X1 U3954 (.ZN(n3851), 
	.B2(n3855), 
	.B1(n3832), 
	.A2(n3830), 
	.A1(n3854));
   AOI22_X1 U3955 (.ZN(n3830), 
	.B2(n5519), 
	.B1(n3077), 
	.A2(n5046), 
	.A1(n3853));
   AOI21_X1 U3956 (.ZN(n3854), 
	.B2(n3856), 
	.B1(n3831), 
	.A(n3829));
   AOI22_X1 U3957 (.ZN(n3829), 
	.B2(n5053), 
	.B1(n3857), 
	.A2(n5009), 
	.A1(n3072));
   INV_X1 U3958 (.ZN(n3856), 
	.A(n3832));
   OAI22_X1 U3959 (.ZN(n3832), 
	.B2(n3853), 
	.B1(n5523), 
	.A2(n3077), 
	.A1(n5023));
   INV_X1 U3960 (.ZN(n3077), 
	.A(n3853));
   NAND3_X1 U3961 (.ZN(n3853), 
	.A3(n3858), 
	.A2(n3060), 
	.A1(n223));
   OAI211_X1 U3962 (.ZN(n3858), 
	.C2(n3860), 
	.C1(n3859), 
	.B(n4799), 
	.A(n3861));
   NOR2_X1 U3964 (.ZN(n3860), 
	.A2(n3720), 
	.A1(n5523));
   AOI211_X1 U3965 (.ZN(n3859), 
	.C2(n3720), 
	.C1(n5523), 
	.B(n5519), 
	.A(n2902));
   INV_X1 U3969 (.ZN(n3831), 
	.A(n3855));
   OAI22_X1 U3970 (.ZN(n3855), 
	.B2(n3072), 
	.B1(n3863), 
	.A2(n3862), 
	.A1(n3857));
   INV_X1 U3971 (.ZN(n3857), 
	.A(n3072));
   INV_X1 U3972 (.ZN(n3850), 
	.A(n3746));
   OAI21_X1 U3973 (.ZN(n3746), 
	.B2(n4797), 
	.B1(n5530), 
	.A(n3072));
   OAI211_X1 U3974 (.ZN(n3072), 
	.C2(n3865), 
	.C1(n3864), 
	.B(n228), 
	.A(n2953));
   OR2_X1 U3977 (.ZN(n3865), 
	.A2(n4797), 
	.A1(n5530));
   AOI22_X1 U3978 (.ZN(n3864), 
	.B2(n3863), 
	.B1(n5010), 
	.A2(n5009), 
	.A1(n3866));
   AOI21_X1 U3979 (.ZN(n3866), 
	.B2(n3862), 
	.B1(n5008), 
	.A(n5053));
   AOI22_X1 U3980 (.ZN(n3621), 
	.B2(n3785), 
	.B1(n2915), 
	.A2(n3786), 
	.A1(n2913));
   INV_X1 U3983 (.ZN(n2913), 
	.A(n3011));
   NAND2_X1 U3985 (.ZN(n2723), 
	.A2(n3538), 
	.A1(n3214));
   INV_X1 U3986 (.ZN(n3214), 
	.A(n3243));
   NAND2_X1 U3987 (.ZN(n3243), 
	.A2(n3213), 
	.A1(n2340));
   INV_X1 U3988 (.ZN(n2340), 
	.A(n2390));
   NAND3_X1 U3989 (.ZN(n2390), 
	.A3(n1773), 
	.A2(n1774), 
	.A1(n3867));
   INV_X1 U3990 (.ZN(n1773), 
	.A(n1780));
   NAND2_X1 U3991 (.ZN(n2062), 
	.A2(n3869), 
	.A1(n3868));
   AOI221_X1 U3992 (.ZN(n3869), 
	.C2(n2879), 
	.C1(hrdata_i[7]), 
	.B2(n231), 
	.B1(n2915), 
	.A(n3870));
   OAI22_X1 U3993 (.ZN(n3870), 
	.B2(n2926), 
	.B1(n3871), 
	.A2(n3011), 
	.A1(n5530));
   AOI221_X1 U3994 (.ZN(n3871), 
	.C2(n3812), 
	.C1(n1890), 
	.B2(n3784), 
	.B1(n1887), 
	.A(n3872));
   OAI22_X1 U3995 (.ZN(n3872), 
	.B2(n2885), 
	.B1(n5549), 
	.A2(n2886), 
	.A1(n5523));
   INV_X1 U3999 (.ZN(n2915), 
	.A(n2948));
   NOR4_X1 U4001 (.ZN(n252), 
	.A4(n5502), 
	.A3(n1110), 
	.A2(n3875), 
	.A1(n3874));
   INV_X1 U4002 (.ZN(n3868), 
	.A(n3876));
   OAI222_X1 U4003 (.ZN(n3876), 
	.C2(FE_PHN2430_n5520), 
	.C1(n16685), 
	.B2(n2998), 
	.B1(n1789), 
	.A2(n2981), 
	.A1(n298));
   OAI22_X1 U4004 (.ZN(n1789), 
	.B2(n2338), 
	.B1(n16788), 
	.A2(n2386), 
	.A1(n2337));
   OAI221_X1 U4005 (.ZN(n2338), 
	.C2(n16951), 
	.C1(n3314), 
	.B2(n16948), 
	.B1(n3329), 
	.A(n3877));
   AOI22_X1 U4006 (.ZN(n3877), 
	.B2(n3155), 
	.B1(n16942), 
	.A2(n3317), 
	.A1(n16945));
   NAND3_X1 U4007 (.ZN(n3155), 
	.A3(n3880), 
	.A2(n3879), 
	.A1(n3878));
   AOI221_X1 U4008 (.ZN(n3880), 
	.C2(vis_r0_o[10]), 
	.C1(n16936), 
	.B2(vis_r2_o[10]), 
	.B1(n16939), 
	.A(n3883));
   OAI22_X1 U4009 (.ZN(n3883), 
	.B2(n16931), 
	.B1(n5445), 
	.A2(n16934), 
	.A1(n5146));
   AOI22_X1 U4011 (.ZN(n3879), 
	.B2(vis_r4_o[10]), 
	.B1(n16924), 
	.A2(vis_r5_o[10]), 
	.A1(n16927));
   AOI22_X1 U4012 (.ZN(n3878), 
	.B2(vis_r1_o[10]), 
	.B1(n16918), 
	.A2(vis_r6_o[10]), 
	.A1(n16921));
   NAND3_X1 U4015 (.ZN(n3317), 
	.A3(n3890), 
	.A2(n3889), 
	.A1(n3888));
   AOI221_X1 U4016 (.ZN(n3890), 
	.C2(vis_r0_o[8]), 
	.C1(FE_OFN644_n16936), 
	.B2(vis_r2_o[8]), 
	.B1(FE_OFN645_n16939), 
	.A(n3893));
   OAI22_X1 U4017 (.ZN(n3893), 
	.B2(n16931), 
	.B1(n5448), 
	.A2(n16934), 
	.A1(n5137));
   AOI22_X1 U4019 (.ZN(n3889), 
	.B2(vis_r4_o[8]), 
	.B1(n16924), 
	.A2(vis_r5_o[8]), 
	.A1(n16927));
   AOI22_X1 U4020 (.ZN(n3888), 
	.B2(vis_r1_o[8]), 
	.B1(n16918), 
	.A2(vis_r6_o[8]), 
	.A1(n16921));
   INV_X1 U4023 (.ZN(n3314), 
	.A(n2209));
   NAND3_X1 U4024 (.ZN(n2209), 
	.A3(n3900), 
	.A2(n3899), 
	.A1(n3898));
   AOI221_X1 U4025 (.ZN(n3900), 
	.C2(vis_r0_o[7]), 
	.C1(n16936), 
	.B2(vis_r2_o[7]), 
	.B1(n16939), 
	.A(n3903));
   OAI22_X1 U4026 (.ZN(n3903), 
	.B2(n16931), 
	.B1(n5423), 
	.A2(n16934), 
	.A1(n5020));
   AOI22_X1 U4029 (.ZN(n3899), 
	.B2(vis_r4_o[7]), 
	.B1(n16925), 
	.A2(vis_r5_o[7]), 
	.A1(n16927));
   AOI22_X1 U4030 (.ZN(n3898), 
	.B2(vis_r1_o[7]), 
	.B1(n16919), 
	.A2(vis_r6_o[7]), 
	.A1(n16922));
   INV_X1 U4033 (.ZN(n3329), 
	.A(n3237));
   NAND3_X1 U4034 (.ZN(n3237), 
	.A3(n3910), 
	.A2(n3909), 
	.A1(n3908));
   AOI221_X1 U4035 (.ZN(n3910), 
	.C2(vis_r0_o[9]), 
	.C1(n16936), 
	.B2(vis_r2_o[9]), 
	.B1(n16939), 
	.A(n3913));
   OAI22_X1 U4036 (.ZN(n3913), 
	.B2(n16931), 
	.B1(n5447), 
	.A2(n16934), 
	.A1(n5143));
   AOI22_X1 U4038 (.ZN(n3909), 
	.B2(vis_r4_o[9]), 
	.B1(n16925), 
	.A2(vis_r5_o[9]), 
	.A1(n16927));
   AOI22_X1 U4039 (.ZN(n3908), 
	.B2(vis_r1_o[9]), 
	.B1(n16919), 
	.A2(vis_r6_o[9]), 
	.A1(n16922));
   OAI221_X1 U4042 (.ZN(n2386), 
	.C2(n16951), 
	.C1(n3328), 
	.B2(n3279), 
	.B1(n3265), 
	.A(n3918));
   AOI22_X1 U4043 (.ZN(n3918), 
	.B2(n3022), 
	.B1(n3275), 
	.A2(n3041), 
	.A1(n16945));
   NAND3_X1 U4044 (.ZN(n3022), 
	.A3(n3921), 
	.A2(n3920), 
	.A1(n3919));
   AOI221_X1 U4045 (.ZN(n3921), 
	.C2(vis_r0_o[13]), 
	.C1(n16936), 
	.B2(vis_r2_o[13]), 
	.B1(n16939), 
	.A(n3924));
   OAI22_X1 U4046 (.ZN(n3924), 
	.B2(n16931), 
	.B1(n5443), 
	.A2(n16934), 
	.A1(n5134));
   AOI22_X1 U4048 (.ZN(n3920), 
	.B2(vis_r4_o[13]), 
	.B1(n16925), 
	.A2(vis_r5_o[13]), 
	.A1(n16927));
   AOI22_X1 U4049 (.ZN(n3919), 
	.B2(vis_r1_o[13]), 
	.B1(n16919), 
	.A2(vis_r6_o[13]), 
	.A1(n16922));
   NAND3_X1 U4052 (.ZN(n3041), 
	.A3(n3931), 
	.A2(n3930), 
	.A1(n3929));
   AOI221_X1 U4053 (.ZN(n3931), 
	.C2(vis_r0_o[12]), 
	.C1(n16936), 
	.B2(vis_r2_o[12]), 
	.B1(n16939), 
	.A(n3934));
   OAI22_X1 U4054 (.ZN(n3934), 
	.B2(n16931), 
	.B1(n5444), 
	.A2(n16934), 
	.A1(n5129));
   AOI22_X1 U4056 (.ZN(n3930), 
	.B2(vis_r4_o[12]), 
	.B1(n16925), 
	.A2(vis_r5_o[12]), 
	.A1(n16927));
   AOI22_X1 U4057 (.ZN(n3929), 
	.B2(vis_r1_o[12]), 
	.B1(n16919), 
	.A2(vis_r6_o[12]), 
	.A1(n16922));
   INV_X1 U4060 (.ZN(n3328), 
	.A(n3134));
   NAND3_X1 U4061 (.ZN(n3134), 
	.A3(n3941), 
	.A2(n3940), 
	.A1(n3939));
   AOI221_X1 U4062 (.ZN(n3941), 
	.C2(vis_r0_o[11]), 
	.C1(n16936), 
	.B2(vis_r2_o[11]), 
	.B1(n16939), 
	.A(n3944));
   OAI22_X1 U4063 (.ZN(n3944), 
	.B2(n16931), 
	.B1(n5557), 
	.A2(n16934), 
	.A1(n5565));
   AOI22_X1 U4065 (.ZN(n3940), 
	.B2(vis_r4_o[11]), 
	.B1(n16925), 
	.A2(vis_r5_o[11]), 
	.A1(n16927));
   AOI22_X1 U4066 (.ZN(n3939), 
	.B2(vis_r1_o[11]), 
	.B1(n16919), 
	.A2(vis_r6_o[11]), 
	.A1(n16922));
   INV_X1 U4069 (.ZN(n3265), 
	.A(n2964));
   NAND3_X1 U4070 (.ZN(n2964), 
	.A3(n3951), 
	.A2(n3950), 
	.A1(n3949));
   AOI221_X1 U4071 (.ZN(n3951), 
	.C2(vis_r0_o[14]), 
	.C1(n16936), 
	.B2(vis_r2_o[14]), 
	.B1(n16939), 
	.A(n3954));
   OAI22_X1 U4072 (.ZN(n3954), 
	.B2(n16931), 
	.B1(n5442), 
	.A2(n16934), 
	.A1(n5105));
   AOI22_X1 U4074 (.ZN(n3950), 
	.B2(vis_r4_o[14]), 
	.B1(n16925), 
	.A2(vis_r5_o[14]), 
	.A1(n16927));
   AOI22_X1 U4075 (.ZN(n3949), 
	.B2(vis_r1_o[14]), 
	.B1(n16919), 
	.A2(vis_r6_o[14]), 
	.A1(n16922));
   OAI21_X1 U4078 (.ZN(n2069), 
	.B2(n3475), 
	.B1(n2389), 
	.A(n3285));
   NAND2_X1 U4079 (.ZN(n3285), 
	.A2(n1574), 
	.A1(n3215));
   NAND2_X1 U4080 (.ZN(n3475), 
	.A2(n3213), 
	.A1(n2358));
   INV_X1 U4081 (.ZN(n2358), 
	.A(n3539));
   NAND3_X1 U4082 (.ZN(n3539), 
	.A3(n1790), 
	.A2(n3867), 
	.A1(n1780));
   OAI21_X1 U4083 (.ZN(n2072), 
	.B2(n3477), 
	.B1(n3215), 
	.A(n3476));
   OAI21_X1 U4084 (.ZN(n3476), 
	.B2(n3959), 
	.B1(n16868), 
	.A(n3215));
   AOI21_X1 U4085 (.ZN(n3959), 
	.B2(n16842), 
	.B1(n16826), 
	.A(n760));
   NAND3_X1 U4086 (.ZN(n3477), 
	.A3(n1780), 
	.A2(n1774), 
	.A1(n3867));
   OAI211_X1 U4088 (.ZN(n2057), 
	.C2(n2375), 
	.C1(n2998), 
	.B(n3960), 
	.A(n2919));
   AOI222_X1 U4089 (.ZN(n3960), 
	.C2(n1066), 
	.C1(n2895), 
	.B2(n3961), 
	.B1(n2882), 
	.A2(n2879), 
	.A1(hrdata_i[31]));
   NAND2_X1 U4092 (.ZN(n3961), 
	.A2(n3964), 
	.A1(n3963));
   AOI222_X1 U4093 (.ZN(n3964), 
	.C2(n3740), 
	.C1(n1191), 
	.B2(n1189), 
	.B1(n3965), 
	.A2(n3791), 
	.A1(n1887));
   NOR2_X1 U4095 (.ZN(n3965), 
	.A2(n2930), 
	.A1(n5504));
   AOI222_X1 U4096 (.ZN(n3963), 
	.C2(n3833), 
	.C1(n1897), 
	.B2(n3792), 
	.B1(n1890), 
	.A2(n3862), 
	.A1(n1893));
   INV_X1 U4097 (.ZN(n1897), 
	.A(n2885));
   INV_X1 U4098 (.ZN(n1893), 
	.A(n2886));
   AND2_X1 U4099 (.ZN(n2919), 
	.A2(n3966), 
	.A1(n3003));
   NAND3_X1 U4100 (.ZN(n3966), 
	.A3(n3967), 
	.A2(n5502), 
	.A1(n3318));
   NOR3_X1 U4101 (.ZN(n3967), 
	.A3(n5017), 
	.A2(n4905), 
	.A1(n5096));
   NOR2_X1 U4102 (.ZN(n3318), 
	.A2(FE_PHN1894_n5149), 
	.A1(n2926));
   NAND2_X1 U4103 (.ZN(n3003), 
	.A2(n14), 
	.A1(n2882));
   NOR3_X1 U4104 (.ZN(n14), 
	.A3(n3875), 
	.A2(n5502), 
	.A1(n2930));
   OAI22_X1 U4105 (.ZN(n2375), 
	.B2(n3969), 
	.B1(n1786), 
	.A2(n3968), 
	.A1(n2313));
   INV_X1 U4106 (.ZN(n3969), 
	.A(n3968));
   INV_X1 U4107 (.ZN(n1786), 
	.A(n3970));
   OAI22_X1 U4108 (.ZN(n3970), 
	.B2(n2334), 
	.B1(n2337), 
	.A2(n2369), 
	.A1(n16788));
   OAI221_X1 U4109 (.ZN(n2334), 
	.C2(n16951), 
	.C1(n3319), 
	.B2(n16948), 
	.B1(n3315), 
	.A(n3971));
   AOI22_X1 U4110 (.ZN(n3971), 
	.B2(n2531), 
	.B1(n16942), 
	.A2(FE_OFN543_n2585), 
	.A1(n16945));
   NAND3_X1 U4111 (.ZN(n2531), 
	.A3(n3974), 
	.A2(n3973), 
	.A1(n3972));
   AOI221_X1 U4112 (.ZN(n3974), 
	.C2(vis_r0_o[6]), 
	.C1(n16936), 
	.B2(vis_r2_o[6]), 
	.B1(n16939), 
	.A(n3977));
   OAI22_X1 U4113 (.ZN(n3977), 
	.B2(n16931), 
	.B1(n5432), 
	.A2(n16934), 
	.A1(n5043));
   AOI22_X1 U4116 (.ZN(n3973), 
	.B2(vis_r4_o[6]), 
	.B1(n16925), 
	.A2(vis_r5_o[6]), 
	.A1(n16927));
   AOI22_X1 U4117 (.ZN(n3972), 
	.B2(vis_r1_o[6]), 
	.B1(n16919), 
	.A2(vis_r6_o[6]), 
	.A1(n16922));
   NAND3_X1 U4120 (.ZN(n2585), 
	.A3(n3984), 
	.A2(n3983), 
	.A1(n3982));
   AOI221_X1 U4121 (.ZN(n3984), 
	.C2(vis_r0_o[4]), 
	.C1(n16936), 
	.B2(vis_r2_o[4]), 
	.B1(n16939), 
	.A(n3987));
   OAI22_X1 U4122 (.ZN(n3987), 
	.B2(n16931), 
	.B1(n5434), 
	.A2(n16934), 
	.A1(n5123));
   AOI22_X1 U4125 (.ZN(n3983), 
	.B2(vis_r4_o[4]), 
	.B1(n16925), 
	.A2(vis_r5_o[4]), 
	.A1(n16927));
   AOI22_X1 U4126 (.ZN(n3982), 
	.B2(vis_r1_o[4]), 
	.B1(n16919), 
	.A2(vis_r6_o[4]), 
	.A1(n16922));
   INV_X1 U4129 (.ZN(n3319), 
	.A(FE_OFN544_n2612));
   NAND3_X1 U4130 (.ZN(n2612), 
	.A3(n3994), 
	.A2(n3993), 
	.A1(n3992));
   AOI221_X1 U4131 (.ZN(n3994), 
	.C2(vis_r0_o[3]), 
	.C1(n16936), 
	.B2(vis_r2_o[3]), 
	.B1(n16939), 
	.A(n3997));
   OAI22_X1 U4132 (.ZN(n3997), 
	.B2(n16931), 
	.B1(n5435), 
	.A2(n16934), 
	.A1(n5030));
   AOI22_X1 U4135 (.ZN(n3993), 
	.B2(vis_r4_o[3]), 
	.B1(n16925), 
	.A2(vis_r5_o[3]), 
	.A1(n16927));
   AOI22_X1 U4136 (.ZN(n3992), 
	.B2(vis_r1_o[3]), 
	.B1(n16919), 
	.A2(vis_r6_o[3]), 
	.A1(n16922));
   INV_X1 U4139 (.ZN(n3315), 
	.A(FE_OFN542_n2562));
   NAND3_X1 U4140 (.ZN(n2562), 
	.A3(n4004), 
	.A2(n4003), 
	.A1(n4002));
   AOI221_X1 U4141 (.ZN(n4004), 
	.C2(vis_r0_o[5]), 
	.C1(n16936), 
	.B2(vis_r2_o[5]), 
	.B1(n16939), 
	.A(n4007));
   OAI22_X1 U4142 (.ZN(n4007), 
	.B2(n16931), 
	.B1(n5433), 
	.A2(n16934), 
	.A1(n5093));
   AOI22_X1 U4145 (.ZN(n4003), 
	.B2(vis_r4_o[5]), 
	.B1(n16925), 
	.A2(vis_r5_o[5]), 
	.A1(n16927));
   AOI22_X1 U4146 (.ZN(n4002), 
	.B2(vis_r1_o[5]), 
	.B1(n16919), 
	.A2(vis_r6_o[5]), 
	.A1(n16922));
   OAI221_X1 U4149 (.ZN(n2369), 
	.C2(n16951), 
	.C1(n3278), 
	.B2(n16948), 
	.B1(n3280), 
	.A(n4012));
   AOI22_X1 U4150 (.ZN(n4012), 
	.B2(FE_OFN560_n3199), 
	.B1(n16942), 
	.A2(n3274), 
	.A1(n16945));
   NAND3_X1 U4151 (.ZN(n3199), 
	.A3(n4015), 
	.A2(n4014), 
	.A1(n4013));
   AOI221_X1 U4152 (.ZN(n4015), 
	.C2(vis_r0_o[2]), 
	.C1(n16936), 
	.B2(vis_r2_o[2]), 
	.B1(n16939), 
	.A(n4018));
   OAI22_X1 U4153 (.ZN(n4018), 
	.B2(n16931), 
	.B1(n5446), 
	.A2(n16934), 
	.A1(n5058));
   AOI22_X1 U4156 (.ZN(n4014), 
	.B2(vis_r4_o[2]), 
	.B1(n16925), 
	.A2(vis_r5_o[2]), 
	.A1(n16927));
   AOI22_X1 U4157 (.ZN(n4013), 
	.B2(vis_r1_o[2]), 
	.B1(n16919), 
	.A2(vis_r6_o[2]), 
	.A1(n16922));
   NAND3_X2 U4160 (.ZN(n3274), 
	.A3(n4025), 
	.A2(n4024), 
	.A1(n4023));
   AOI221_X2 U4161 (.ZN(n4025), 
	.C2(vis_r0_o[0]), 
	.C1(n16936), 
	.B2(vis_r2_o[0]), 
	.B1(n16939), 
	.A(n4028));
   OAI22_X2 U4162 (.ZN(n4028), 
	.B2(n16930), 
	.B1(n5425), 
	.A2(n16933), 
	.A1(n5038));
   AOI22_X2 U4165 (.ZN(n4024), 
	.B2(vis_r4_o[0]), 
	.B1(n16924), 
	.A2(vis_r5_o[0]), 
	.A1(n16927));
   AOI22_X2 U4166 (.ZN(n4023), 
	.B2(vis_r1_o[0]), 
	.B1(n16918), 
	.A2(vis_r6_o[0]), 
	.A1(n16921));
   INV_X1 U4169 (.ZN(n3278), 
	.A(n3400));
   INV_X1 U4170 (.ZN(n3280), 
	.A(n2639));
   NAND3_X1 U4171 (.ZN(n2639), 
	.A3(n4035), 
	.A2(n4034), 
	.A1(n4033));
   AOI221_X1 U4172 (.ZN(n4035), 
	.C2(vis_r0_o[1]), 
	.C1(n16936), 
	.B2(vis_r2_o[1]), 
	.B1(n16939), 
	.A(n4038));
   OAI22_X1 U4173 (.ZN(n4038), 
	.B2(n16930), 
	.B1(n5424), 
	.A2(n16933), 
	.A1(n4985));
   AOI22_X1 U4176 (.ZN(n4034), 
	.B2(vis_r4_o[1]), 
	.B1(n16924), 
	.A2(vis_r5_o[1]), 
	.A1(n16927));
   AOI22_X1 U4177 (.ZN(n4033), 
	.B2(vis_r1_o[1]), 
	.B1(n16918), 
	.A2(vis_r6_o[1]), 
	.A1(n16921));
   AOI22_X1 U4180 (.ZN(n3968), 
	.B2(n2941), 
	.B1(n16951), 
	.A2(n2940), 
	.A1(n3118));
   NOR2_X1 U4181 (.ZN(n2941), 
	.A2(FE_OFN631_n16851), 
	.A1(n3120));
   INV_X1 U4182 (.ZN(n2940), 
	.A(n3091));
   OAI211_X1 U4183 (.ZN(n3091), 
	.C2(n16788), 
	.C1(n3120), 
	.B(FE_OFN87_n16848), 
	.A(n3119));
   NAND2_X1 U4184 (.ZN(n3119), 
	.A2(n16788), 
	.A1(n3120));
   INV_X1 U4185 (.ZN(n3120), 
	.A(n3343));
   NAND2_X1 U4186 (.ZN(n3343), 
	.A2(n3478), 
	.A1(n3538));
   NAND4_X1 U4187 (.ZN(n3478), 
	.A4(n1774), 
	.A3(n1780), 
	.A2(n2337), 
	.A1(n3118));
   INV_X1 U4188 (.ZN(n2313), 
	.A(n3092));
   NAND3_X1 U4189 (.ZN(n3092), 
	.A3(n4043), 
	.A2(n1759), 
	.A1(n3400));
   OAI21_X1 U4190 (.ZN(n4043), 
	.B2(FE_OFN100_n1086), 
	.B1(n16828), 
	.A(n1784));
   NAND3_X1 U4191 (.ZN(n3400), 
	.A3(n4046), 
	.A2(n4045), 
	.A1(n4044));
   AOI221_X1 U4192 (.ZN(n4046), 
	.C2(vis_r0_o[31]), 
	.C1(n16936), 
	.B2(vis_r2_o[31]), 
	.B1(n16939), 
	.A(n4049));
   OAI22_X1 U4193 (.ZN(n4049), 
	.B2(n16930), 
	.B1(n5421), 
	.A2(n16933), 
	.A1(n4962));
   AOI22_X1 U4195 (.ZN(n4045), 
	.B2(vis_r4_o[31]), 
	.B1(n16924), 
	.A2(vis_r5_o[31]), 
	.A1(n16927));
   AOI22_X1 U4196 (.ZN(n4044), 
	.B2(vis_r1_o[31]), 
	.B1(n16918), 
	.A2(vis_r6_o[31]), 
	.A1(n16921));
   OAI21_X1 U4199 (.ZN(n2067), 
	.B2(n1027), 
	.B1(n3213), 
	.A(n3472));
   NAND2_X1 U4200 (.ZN(n3472), 
	.A2(n3213), 
	.A1(n2322));
   NOR2_X1 U4201 (.ZN(n2322), 
	.A2(n2389), 
	.A1(n3217));
   INV_X1 U4202 (.ZN(n2389), 
	.A(n3538));
   NAND2_X1 U4203 (.ZN(n3538), 
	.A2(n918), 
	.A1(FE_OFN79_n16834));
   NAND2_X1 U4205 (.ZN(n3867), 
	.A2(FE_OFN89_n16849), 
	.A1(n1793));
   OAI21_X1 U4206 (.ZN(n1793), 
	.B2(n1519), 
	.B1(n4054), 
	.A(n4055));
   NAND4_X1 U4207 (.ZN(n4055), 
	.A4(n4057), 
	.A3(n4056), 
	.A2(n16833), 
	.A1(n563));
   NOR3_X1 U4208 (.ZN(n4057), 
	.A3(n795), 
	.A2(FE_OFN15_n16671), 
	.A1(n16656));
   INV_X1 U4209 (.ZN(n4056), 
	.A(n3566));
   NOR3_X1 U4211 (.ZN(n4054), 
	.A3(n1795), 
	.A2(FE_OFN565_n4058), 
	.A1(n1794));
   NOR2_X1 U4212 (.ZN(n1777), 
	.A2(n1780), 
	.A1(n1774));
   OAI21_X1 U4213 (.ZN(n1780), 
	.B2(n4059), 
	.B1(n16828), 
	.A(n4060));
   OAI21_X1 U4214 (.ZN(n4060), 
	.B2(n1763), 
	.B1(n4061), 
	.A(n16831));
   AND3_X1 U4215 (.ZN(n1763), 
	.A3(n4064), 
	.A2(n4063), 
	.A1(n4062));
   AOI21_X1 U4216 (.ZN(n4061), 
	.B2(n4063), 
	.B1(n4062), 
	.A(n4064));
   INV_X1 U4217 (.ZN(n4059), 
	.A(n4064));
   AOI22_X1 U4218 (.ZN(n4064), 
	.B2(n529), 
	.B1(FE_OFN566_n4065), 
	.A2(n563), 
	.A1(FE_OFN15_n16671));
   INV_X1 U4219 (.ZN(n1774), 
	.A(n1790));
   AOI22_X1 U4220 (.ZN(n1790), 
	.B2(n4066), 
	.B1(n16828), 
	.A2(n4063), 
	.A1(n16833));
   XNOR2_X1 U4221 (.ZN(n4066), 
	.B(n4062), 
	.A(n4063));
   AND2_X1 U4222 (.ZN(n4062), 
	.A2(n4068), 
	.A1(n4067));
   AOI22_X1 U4223 (.ZN(n4063), 
	.B2(n529), 
	.B1(FE_OFN567_n4069), 
	.A2(n563), 
	.A1(n795));
   NAND2_X2 U4225 (.ZN(n1027), 
	.A2(n16842), 
	.A1(n195));
   NAND2_X1 U4227 (.ZN(n4070), 
	.A2(n616), 
	.A1(n624));
   OAI221_X1 U4228 (.ZN(n2061), 
	.C2(n264), 
	.C1(n2981), 
	.B2(n262), 
	.B1(n16685), 
	.A(n4071));
   AOI222_X1 U4229 (.ZN(n4071), 
	.C2(n2879), 
	.C1(hrdata_i[23]), 
	.B2(n4072), 
	.B1(n2882), 
	.A2(n2922), 
	.A1(n1787));
   AND3_X1 U4232 (.ZN(n1111), 
	.A3(n1189), 
	.A2(n5096), 
	.A1(n4905));
   NOR2_X1 U4233 (.ZN(n1189), 
	.A2(n3875), 
	.A1(n4073));
   OAI221_X1 U4234 (.ZN(n4072), 
	.C2(n2886), 
	.C1(n5008), 
	.B2(n2885), 
	.B1(n5551), 
	.A(n4074));
   AOI222_X1 U4235 (.ZN(n4074), 
	.C2(n3790), 
	.C1(n1887), 
	.B2(n3731), 
	.B1(n1191), 
	.A2(n3793), 
	.A1(n1890));
   INV_X1 U4237 (.ZN(n1887), 
	.A(n2898));
   NAND3_X1 U4238 (.ZN(n2898), 
	.A3(n1188), 
	.A2(n3875), 
	.A1(n4073));
   INV_X1 U4239 (.ZN(n1188), 
	.A(n2930));
   NAND3_X1 U4240 (.ZN(n2930), 
	.A3(FE_PHN1894_n5149), 
	.A2(n251), 
	.A1(n3874));
   AND3_X1 U4242 (.ZN(n1191), 
	.A3(n4075), 
	.A2(n4073), 
	.A1(n5017));
   INV_X1 U4244 (.ZN(n1890), 
	.A(n2899));
   NAND3_X1 U4245 (.ZN(n2899), 
	.A3(n4076), 
	.A2(FE_PHN1894_n5149), 
	.A1(n4905));
   NOR3_X1 U4246 (.ZN(n4076), 
	.A3(n5096), 
	.A2(n5017), 
	.A1(n5502));
   NAND3_X1 U4247 (.ZN(n2886), 
	.A3(n3717), 
	.A2(n251), 
	.A1(n3875));
   NAND3_X1 U4248 (.ZN(n2885), 
	.A3(n4905), 
	.A2(n3875), 
	.A1(n3717));
   OAI211_X1 U4251 (.ZN(n4077), 
	.C2(n526), 
	.C1(n16845), 
	.B(n3546), 
	.A(FE_OFN483_n1233));
   NAND2_X1 U4252 (.ZN(n3546), 
	.A2(FE_OFN70_n16867), 
	.A1(FE_OFN73_n16806));
   INV_X1 U4253 (.ZN(n1787), 
	.A(n2346));
   OAI22_X1 U4254 (.ZN(n2346), 
	.B2(n3117), 
	.B1(n2337), 
	.A2(n2356), 
	.A1(n16788));
   OAI221_X1 U4255 (.ZN(n3117), 
	.C2(n16951), 
	.C1(n3338), 
	.B2(n16948), 
	.B1(n3341), 
	.A(n4078));
   AOI22_X1 U4256 (.ZN(n4078), 
	.B2(n2297), 
	.B1(n16942), 
	.A2(n2271), 
	.A1(n16945));
   NAND3_X1 U4257 (.ZN(n2297), 
	.A3(n4081), 
	.A2(n4080), 
	.A1(n4079));
   AOI221_X1 U4258 (.ZN(n4081), 
	.C2(vis_r0_o[30]), 
	.C1(n16936), 
	.B2(vis_r2_o[30]), 
	.B1(n16939), 
	.A(n4084));
   OAI22_X1 U4259 (.ZN(n4084), 
	.B2(n16930), 
	.B1(n5426), 
	.A2(n16933), 
	.A1(n5082));
   AOI22_X1 U4261 (.ZN(n4080), 
	.B2(vis_r4_o[30]), 
	.B1(n16924), 
	.A2(vis_r5_o[30]), 
	.A1(n16927));
   AOI22_X1 U4262 (.ZN(n4079), 
	.B2(vis_r1_o[30]), 
	.B1(n16918), 
	.A2(vis_r6_o[30]), 
	.A1(n16921));
   NAND3_X1 U4265 (.ZN(n2271), 
	.A3(n4091), 
	.A2(n4090), 
	.A1(n4089));
   AOI221_X1 U4266 (.ZN(n4091), 
	.C2(vis_r0_o[28]), 
	.C1(n16936), 
	.B2(vis_r2_o[28]), 
	.B1(n16939), 
	.A(n4094));
   OAI22_X1 U4267 (.ZN(n4094), 
	.B2(n16930), 
	.B1(n5422), 
	.A2(n16933), 
	.A1(n4996));
   AOI22_X1 U4269 (.ZN(n4090), 
	.B2(vis_r4_o[28]), 
	.B1(n16924), 
	.A2(vis_r5_o[28]), 
	.A1(n16927));
   AOI22_X1 U4270 (.ZN(n4089), 
	.B2(vis_r1_o[28]), 
	.B1(n16918), 
	.A2(vis_r6_o[28]), 
	.A1(n16921));
   INV_X1 U4273 (.ZN(n3338), 
	.A(n2433));
   NAND3_X1 U4274 (.ZN(n2433), 
	.A3(n4101), 
	.A2(n4100), 
	.A1(n4099));
   AOI221_X1 U4275 (.ZN(n4101), 
	.C2(vis_r0_o[27]), 
	.C1(n16936), 
	.B2(vis_r2_o[27]), 
	.B1(n16939), 
	.A(n4104));
   OAI22_X1 U4276 (.ZN(n4104), 
	.B2(n16930), 
	.B1(n5428), 
	.A2(n16933), 
	.A1(n5113));
   AOI22_X1 U4278 (.ZN(n4100), 
	.B2(vis_r4_o[27]), 
	.B1(n16924), 
	.A2(vis_r5_o[27]), 
	.A1(n16927));
   AOI22_X1 U4279 (.ZN(n4099), 
	.B2(vis_r1_o[27]), 
	.B1(n16918), 
	.A2(vis_r6_o[27]), 
	.A1(n16921));
   INV_X1 U4282 (.ZN(n3341), 
	.A(n2402));
   NAND3_X1 U4283 (.ZN(n2402), 
	.A3(n4111), 
	.A2(n4110), 
	.A1(n4109));
   AOI221_X1 U4284 (.ZN(n4111), 
	.C2(vis_r0_o[29]), 
	.C1(n16936), 
	.B2(vis_r2_o[29]), 
	.B1(n16939), 
	.A(n4114));
   OAI22_X1 U4285 (.ZN(n4114), 
	.B2(n16930), 
	.B1(n5427), 
	.A2(n16933), 
	.A1(n5077));
   AOI22_X1 U4287 (.ZN(n4110), 
	.B2(vis_r4_o[29]), 
	.B1(n16924), 
	.A2(vis_r5_o[29]), 
	.A1(n16927));
   AOI22_X1 U4288 (.ZN(n4109), 
	.B2(vis_r1_o[29]), 
	.B1(n16918), 
	.A2(vis_r6_o[29]), 
	.A1(n16921));
   OAI221_X1 U4292 (.ZN(n2356), 
	.C2(n16951), 
	.C1(n3345), 
	.B2(n16948), 
	.B1(n3339), 
	.A(n4119));
   AOI22_X1 U4293 (.ZN(n4119), 
	.B2(n2452), 
	.B1(n16942), 
	.A2(n2507), 
	.A1(n16945));
   NAND3_X1 U4294 (.ZN(n2452), 
	.A3(n4122), 
	.A2(n4121), 
	.A1(n4120));
   AOI221_X1 U4295 (.ZN(n4122), 
	.C2(vis_r0_o[26]), 
	.C1(n16936), 
	.B2(vis_r2_o[26]), 
	.B1(n16939), 
	.A(n4125));
   OAI22_X1 U4296 (.ZN(n4125), 
	.B2(n16930), 
	.B1(n5429), 
	.A2(n16933), 
	.A1(n4991));
   AOI22_X1 U4298 (.ZN(n4121), 
	.B2(vis_r4_o[26]), 
	.B1(n16924), 
	.A2(vis_r5_o[26]), 
	.A1(n16927));
   AOI22_X1 U4299 (.ZN(n4120), 
	.B2(vis_r1_o[26]), 
	.B1(n16918), 
	.A2(vis_r6_o[26]), 
	.A1(n16921));
   NAND2_X1 U4303 (.ZN(n3279), 
	.A2(n4131), 
	.A1(n4130));
   NAND3_X1 U4304 (.ZN(n2507), 
	.A3(n4134), 
	.A2(n4133), 
	.A1(n4132));
   AOI221_X1 U4305 (.ZN(n4134), 
	.C2(vis_r0_o[24]), 
	.C1(n16936), 
	.B2(vis_r2_o[24]), 
	.B1(n16939), 
	.A(n4137));
   OAI22_X1 U4306 (.ZN(n4137), 
	.B2(n16930), 
	.B1(n5431), 
	.A2(n16933), 
	.A1(n4972));
   AOI22_X1 U4308 (.ZN(n4133), 
	.B2(vis_r4_o[24]), 
	.B1(n16924), 
	.A2(vis_r5_o[24]), 
	.A1(n16927));
   AOI22_X1 U4309 (.ZN(n4132), 
	.B2(vis_r1_o[24]), 
	.B1(n16918), 
	.A2(vis_r6_o[24]), 
	.A1(n16921));
   NAND2_X1 U4313 (.ZN(n3277), 
	.A2(n4142), 
	.A1(n4131));
   INV_X1 U4316 (.ZN(n3345), 
	.A(n3254));
   NAND3_X1 U4317 (.ZN(n3254), 
	.A3(n4145), 
	.A2(n4144), 
	.A1(n4143));
   AOI221_X1 U4318 (.ZN(n4145), 
	.C2(vis_r0_o[23]), 
	.C1(n16936), 
	.B2(vis_r2_o[23]), 
	.B1(n16939), 
	.A(n4148));
   OAI22_X1 U4319 (.ZN(n4148), 
	.B2(n16930), 
	.B1(n5585), 
	.A2(n16933), 
	.A1(n4960));
   AOI22_X1 U4321 (.ZN(n4144), 
	.B2(vis_r4_o[23]), 
	.B1(n16924), 
	.A2(vis_r5_o[23]), 
	.A1(n16927));
   AOI22_X1 U4322 (.ZN(n4143), 
	.B2(vis_r1_o[23]), 
	.B1(n16918), 
	.A2(vis_r6_o[23]), 
	.A1(n16921));
   INV_X1 U4327 (.ZN(n4142), 
	.A(n4130));
   AOI221_X1 U4328 (.ZN(n4130), 
	.C2(n4155), 
	.C1(n16833), 
	.B2(n4154), 
	.B1(n4153), 
	.A(n4067));
   INV_X1 U4329 (.ZN(n4155), 
	.A(n4153));
   AND2_X1 U4330 (.ZN(n4154), 
	.A2(n16828), 
	.A1(n4131));
   INV_X1 U4331 (.ZN(n3339), 
	.A(n2484));
   NAND3_X1 U4332 (.ZN(n2484), 
	.A3(n4158), 
	.A2(n4157), 
	.A1(n4156));
   AOI221_X1 U4333 (.ZN(n4158), 
	.C2(vis_r0_o[25]), 
	.C1(n16936), 
	.B2(vis_r2_o[25]), 
	.B1(n16939), 
	.A(n4161));
   OAI22_X1 U4334 (.ZN(n4161), 
	.B2(n16930), 
	.B1(n5430), 
	.A2(n16933), 
	.A1(n5014));
   NOR3_X1 U4337 (.ZN(n4162), 
	.A3(n3495), 
	.A2(n4978), 
	.A1(FE_OFN583_n5036));
   NOR3_X1 U4341 (.ZN(n4163), 
	.A3(n3492), 
	.A2(n3495), 
	.A1(n3488));
   AOI22_X1 U4342 (.ZN(n4157), 
	.B2(vis_r4_o[25]), 
	.B1(n16924), 
	.A2(vis_r5_o[25]), 
	.A1(n16927));
   AOI22_X1 U4346 (.ZN(n4156), 
	.B2(vis_r1_o[25]), 
	.B1(n16918), 
	.A2(vis_r6_o[25]), 
	.A1(n16921));
   NOR2_X1 U4349 (.ZN(n3592), 
	.A2(n4978), 
	.A1(n3480));
   NOR2_X1 U4356 (.ZN(n4168), 
	.A2(n16833), 
	.A1(n4067));
   NOR2_X1 U4357 (.ZN(n4067), 
	.A2(n4153), 
	.A1(n4131));
   OAI22_X1 U4358 (.ZN(n4153), 
	.B2(n1519), 
	.B1(n4169), 
	.A2(n1234), 
	.A1(n5027));
   OAI22_X1 U4359 (.ZN(n4131), 
	.B2(n1519), 
	.B1(n4170), 
	.A2(n1234), 
	.A1(n5120));
   AOI22_X1 U4360 (.ZN(n4068), 
	.B2(n529), 
	.B1(n4171), 
	.A2(n563), 
	.A1(n16656));
   NAND2_X1 U4361 (.ZN(n2981), 
	.A2(n2882), 
	.A1(n316));
   AND3_X1 U4363 (.ZN(n316), 
	.A3(n4075), 
	.A2(n3875), 
	.A1(n5502));
   NOR3_X1 U4364 (.ZN(n4075), 
	.A3(n251), 
	.A2(n5096), 
	.A1(FE_PHN1894_n5149));
   NAND4_X1 U4368 (.ZN(n261), 
	.A4(n3875), 
	.A3(FE_PHN1894_n5149), 
	.A2(n5096), 
	.A1(n5502));
   OAI211_X1 U4371 (.ZN(n4172), 
	.C2(n1964), 
	.C1(n16845), 
	.B(n4174), 
	.A(n4173));
   AOI21_X1 U4372 (.ZN(n4174), 
	.B2(n16868), 
	.B1(n1262), 
	.A(n17096));
   INV_X1 U4373 (.ZN(n1262), 
	.A(n616));
   NAND3_X1 U4375 (.ZN(n4173), 
	.A3(n757), 
	.A2(FE_OFN95_n16864), 
	.A1(n16845));
   INV_X1 U4376 (.ZN(n757), 
	.A(n624));
   NAND2_X1 U4377 (.ZN(n624), 
	.A2(n16871), 
	.A1(n16680));
   NAND2_X1 U4378 (.ZN(n1964), 
	.A2(n16838), 
	.A1(n526));
   AOI21_X1 U4380 (.ZN(n2085), 
	.B2(n1508), 
	.B1(n84), 
	.A(FE_PHN674_n17127));
   AOI21_X1 U4382 (.ZN(n1508), 
	.B2(n16871), 
	.B1(n4175), 
	.A(n3516));
   NOR2_X1 U4383 (.ZN(n3516), 
	.A2(n1519), 
	.A1(n758));
   OR4_X1 U4384 (.ZN(n4175), 
	.A4(n4177), 
	.A3(n4176), 
	.A2(n1803), 
	.A1(n1801));
   OAI222_X1 U4385 (.ZN(n4177), 
	.C2(FE_OFN98_n1104), 
	.C1(n653), 
	.B2(n16859), 
	.B1(n849), 
	.A2(n1579), 
	.A1(FE_OFN91_n16864));
   OAI21_X1 U4386 (.ZN(n4176), 
	.B2(n16824), 
	.B1(n4178), 
	.A(n1230));
   NAND2_X1 U4387 (.ZN(n1230), 
	.A2(n16851), 
	.A1(FE_OFN70_n16867));
   NOR2_X1 U4388 (.ZN(n1803), 
	.A2(FE_OFN79_n16834), 
	.A1(FE_OFN91_n16864));
   AND3_X1 U4389 (.ZN(n1801), 
	.A3(n4179), 
	.A2(n16828), 
	.A1(n4178));
   INV_X1 U4390 (.ZN(n4178), 
	.A(n1606));
   NOR2_X1 U4391 (.ZN(n1606), 
	.A2(FE_OFN100_n1086), 
	.A1(n16842));
   NOR2_X1 U4392 (.ZN(n84), 
	.A2(n86), 
	.A1(n88));
   NOR2_X1 U4393 (.ZN(n86), 
	.A2(n1040), 
	.A1(n499));
   NOR3_X1 U4394 (.ZN(n88), 
	.A3(n16656), 
	.A2(n1348), 
	.A1(FE_OFN15_n16671));
   INV_X1 U4396 (.ZN(n1348), 
	.A(n2027));
   OAI21_X1 U4397 (.ZN(n2027), 
	.B2(n891), 
	.B1(n16851), 
	.A(n4180));
   NAND3_X1 U4398 (.ZN(n4180), 
	.A3(n563), 
	.A2(n16862), 
	.A1(n566));
   NOR2_X1 U4399 (.ZN(n566), 
	.A2(FE_OFN79_n16834), 
	.A1(n851));
   NAND2_X2 U4400 (.ZN(n891), 
	.A2(n17096), 
	.A1(n760));
   OAI22_X1 U4401 (.ZN(U227_Z_0), 
	.B2(n1096), 
	.B1(n4182), 
	.A2(n4181), 
	.A1(n4956));
   NOR4_X1 U4403 (.ZN(n4182), 
	.A4(txev_o), 
	.A3(rxev_i), 
	.A2(n17092), 
	.A1(n4183));
   OAI21_X1 U4405 (.ZN(n4183), 
	.B2(n4184), 
	.B1(n5168), 
	.A(n1314));
   NOR2_X2 U4407 (.ZN(n1125), 
	.A2(n605), 
	.A1(n1092));
   NAND2_X2 U4408 (.ZN(n605), 
	.A2(n16855), 
	.A1(n16851));
   NAND2_X1 U4409 (.ZN(n1092), 
	.A2(n527), 
	.A1(n997));
   NOR4_X1 U4410 (.ZN(n4184), 
	.A4(n4188), 
	.A3(n4187), 
	.A2(n4186), 
	.A1(n4185));
   INV_X1 U4411 (.ZN(n4188), 
	.A(n4189));
   AOI222_X1 U4412 (.ZN(n4189), 
	.C2(n11929), 
	.C1(n5005), 
	.B2(n4893), 
	.B1(n5526), 
	.A2(FE_PHN1502_n11928), 
	.A1(n4965));
   AOI21_X1 U4413 (.ZN(n11929), 
	.B2(n17092), 
	.B1(n1318), 
	.A(FE_PHN1354_n4190));
   AOI21_X1 U4414 (.ZN(n4190), 
	.B2(FE_PHN2985_IRQ_0_), 
	.B1(n1310), 
	.A(n4191));
   AOI22_X1 U4415 (.ZN(n4191), 
	.B2(n4192), 
	.B1(hwdata_o[0]), 
	.A2(n5005), 
	.A1(n1316));
   NAND2_X1 U4416 (.ZN(n1316), 
	.A2(n1124), 
	.A1(hwdata_o[0]));
   AOI21_X1 U4420 (.ZN(n4893), 
	.B2(n17092), 
	.B1(n1392), 
	.A(FE_PHN1344_n4193));
   AOI21_X1 U4421 (.ZN(n4193), 
	.B2(n5525), 
	.B1(FE_PHN2991_IRQ_3_), 
	.A(n4194));
   AOI22_X1 U4422 (.ZN(n4194), 
	.B2(n4192), 
	.B1(hwdata_o[3]), 
	.A2(n5526), 
	.A1(n1390));
   NAND2_X1 U4423 (.ZN(n1390), 
	.A2(n1124), 
	.A1(hwdata_o[3]));
   AOI21_X1 U4426 (.ZN(n11928), 
	.B2(n4195), 
	.B1(n4965), 
	.A(n1429));
   NOR2_X1 U4427 (.ZN(n1429), 
	.A2(n183), 
	.A1(n200));
   NAND2_X1 U4428 (.ZN(n183), 
	.A2(n186), 
	.A1(n1343));
   AOI21_X1 U4429 (.ZN(n4195), 
	.B2(FE_PHN4631_NMI), 
	.B1(n4964), 
	.A(n1428));
   NOR2_X1 U4430 (.ZN(n1428), 
	.A2(n3962), 
	.A1(n1187));
   OAI221_X1 U4431 (.ZN(n4187), 
	.C2(n4196), 
	.C1(n3238), 
	.B2(n3066), 
	.B1(n1012), 
	.A(n4197));
   OAI21_X1 U4432 (.ZN(n4197), 
	.B2(n4199), 
	.B1(n4198), 
	.A(n1124));
   NAND4_X1 U4433 (.ZN(n4199), 
	.A4(n4201), 
	.A3(n4200), 
	.A2(n1190), 
	.A1(n19));
   NOR3_X1 U4434 (.ZN(n4201), 
	.A3(hwdata_o[21]), 
	.A2(hwdata_o[19]), 
	.A1(hwdata_o[30]));
   NAND4_X2 U4437 (.ZN(n21), 
	.A4(n4207), 
	.A3(n4206), 
	.A2(n4205), 
	.A1(n4204));
   AOI221_X1 U4438 (.ZN(n4207), 
	.C2(vis_r5_o[21]), 
	.C1(n16913), 
	.B2(vis_r4_o[21]), 
	.B1(n16916), 
	.A(n4210));
   OAI222_X1 U4439 (.ZN(n4210), 
	.C2(n16905), 
	.C1(n5466), 
	.B2(n16908), 
	.B1(n5185), 
	.A2(n16910), 
	.A1(n4765));
   AOI221_X1 U4442 (.ZN(n4206), 
	.C2(vis_r10_o[21]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[19]), 
	.B1(n16902), 
	.A(n4216));
   OAI22_X1 U4443 (.ZN(n4216), 
	.B2(n16893), 
	.B1(n5623), 
	.A2(n16895), 
	.A1(n5622));
   AOI221_X1 U4446 (.ZN(n4205), 
	.C2(vis_r12_o[21]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[21]), 
	.B1(FE_OFN638_n16891), 
	.A(n4221));
   OAI22_X1 U4447 (.ZN(n4221), 
	.B2(n16882), 
	.B1(n5408), 
	.A2(n16885), 
	.A1(n5115));
   AOI221_X1 U4450 (.ZN(n4204), 
	.C2(vis_r3_o[21]), 
	.C1(FE_OFN635_n16877), 
	.B2(vis_r0_o[21]), 
	.B1(n4224), 
	.A(n4227));
   OAI22_X1 U4451 (.ZN(n4227), 
	.B2(n16873), 
	.B1(n5321), 
	.A2(n16875), 
	.A1(n5117));
   NAND4_X2 U4456 (.ZN(n22), 
	.A4(n4233), 
	.A3(n4232), 
	.A2(n4231), 
	.A1(n4230));
   AOI221_X1 U4457 (.ZN(n4233), 
	.C2(vis_r5_o[19]), 
	.C1(n16913), 
	.B2(vis_r4_o[19]), 
	.B1(n16916), 
	.A(n4234));
   OAI222_X1 U4458 (.ZN(n4234), 
	.C2(n16905), 
	.C1(n5467), 
	.B2(n16908), 
	.B1(n5186), 
	.A2(n16910), 
	.A1(n4767));
   AOI221_X1 U4461 (.ZN(n4232), 
	.C2(vis_r10_o[19]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[17]), 
	.B1(n16902), 
	.A(n4235));
   OAI22_X1 U4462 (.ZN(n4235), 
	.B2(n16893), 
	.B1(n5637), 
	.A2(n16895), 
	.A1(n5636));
   AOI221_X1 U4465 (.ZN(n4231), 
	.C2(vis_r12_o[19]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[19]), 
	.B1(FE_OFN638_n16891), 
	.A(n4236));
   OAI22_X1 U4466 (.ZN(n4236), 
	.B2(n16882), 
	.B1(n5409), 
	.A2(n16885), 
	.A1(n5088));
   AOI221_X1 U4469 (.ZN(n4230), 
	.C2(vis_r3_o[19]), 
	.C1(FE_OFN635_n16877), 
	.B2(vis_r0_o[19]), 
	.B1(n4224), 
	.A(n4238));
   OAI22_X1 U4470 (.ZN(n4238), 
	.B2(n16873), 
	.B1(n5322), 
	.A2(n16875), 
	.A1(n5090));
   INV_X1 U4475 (.ZN(n4200), 
	.A(n18));
   NAND3_X1 U4476 (.ZN(n18), 
	.A3(n4241), 
	.A2(n1115), 
	.A1(n1187));
   NOR3_X1 U4477 (.ZN(n4241), 
	.A3(hwdata_o[27]), 
	.A2(hwdata_o[28]), 
	.A1(hwdata_o[25]));
   AOI222_X1 U4479 (.ZN(n208), 
	.C2(n4203), 
	.C1(n2427), 
	.B2(n4240), 
	.B1(n2246), 
	.A2(n4239), 
	.A1(n2257));
   AOI222_X1 U4482 (.ZN(n201), 
	.C2(n4239), 
	.C1(n2028), 
	.B2(n4203), 
	.B1(n2248), 
	.A2(n4240), 
	.A1(n3287));
   NAND4_X1 U4483 (.ZN(n2248), 
	.A4(n4245), 
	.A3(n4244), 
	.A2(n4243), 
	.A1(n4242));
   AOI221_X1 U4484 (.ZN(n4245), 
	.C2(vis_r5_o[25]), 
	.C1(n16913), 
	.B2(vis_r4_o[25]), 
	.B1(n16916), 
	.A(n4246));
   OAI222_X1 U4485 (.ZN(n4246), 
	.C2(n16905), 
	.C1(n5459), 
	.B2(n16908), 
	.B1(n5178), 
	.A2(n16910), 
	.A1(n4763));
   AOI221_X1 U4488 (.ZN(n4244), 
	.C2(vis_r10_o[25]), 
	.C1(n16897), 
	.B2(vis_psp_o[23]), 
	.B1(n16902), 
	.A(n4247));
   OAI22_X1 U4489 (.ZN(n4247), 
	.B2(n16893), 
	.B1(n5015), 
	.A2(n16895), 
	.A1(n5291));
   AOI221_X1 U4492 (.ZN(n4243), 
	.C2(vis_r12_o[25]), 
	.C1(n16886), 
	.B2(vis_r9_o[25]), 
	.B1(n16891), 
	.A(n4248));
   OAI22_X1 U4493 (.ZN(n4248), 
	.B2(n16882), 
	.B1(n5401), 
	.A2(n16885), 
	.A1(n5012));
   AOI221_X1 U4496 (.ZN(n4242), 
	.C2(vis_r3_o[25]), 
	.C1(n16877), 
	.B2(vis_r0_o[25]), 
	.B1(n4224), 
	.A(n4250));
   OAI22_X1 U4497 (.ZN(n4250), 
	.B2(n16873), 
	.B1(n5314), 
	.A2(n16875), 
	.A1(n5014));
   NAND4_X2 U4501 (.ZN(n2249), 
	.A4(n4254), 
	.A3(n4253), 
	.A2(n4252), 
	.A1(n4251));
   AOI221_X1 U4502 (.ZN(n4254), 
	.C2(vis_r5_o[18]), 
	.C1(n16913), 
	.B2(vis_r4_o[18]), 
	.B1(n16916), 
	.A(n4255));
   OAI222_X1 U4503 (.ZN(n4255), 
	.C2(n16905), 
	.C1(n5468), 
	.B2(n16908), 
	.B1(n5187), 
	.A2(n16910), 
	.A1(n4768));
   AOI221_X1 U4506 (.ZN(n4253), 
	.C2(vis_r10_o[18]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[16]), 
	.B1(n16902), 
	.A(n4256));
   OAI22_X1 U4507 (.ZN(n4256), 
	.B2(n16893), 
	.B1(n5065), 
	.A2(n16895), 
	.A1(n5297));
   AOI221_X1 U4510 (.ZN(n4252), 
	.C2(vis_r12_o[18]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[18]), 
	.B1(FE_OFN638_n16891), 
	.A(n4257));
   OAI22_X1 U4511 (.ZN(n4257), 
	.B2(n16882), 
	.B1(n5410), 
	.A2(n16885), 
	.A1(n5062));
   AOI221_X1 U4514 (.ZN(n4251), 
	.C2(vis_r3_o[18]), 
	.C1(FE_OFN635_n16877), 
	.B2(vis_r0_o[18]), 
	.B1(n4224), 
	.A(n4259));
   OAI22_X1 U4515 (.ZN(n4259), 
	.B2(n16873), 
	.B1(n5323), 
	.A2(n16875), 
	.A1(n5064));
   NAND2_X2 U4518 (.ZN(n1187), 
	.A2(hwdata_o[31]), 
	.A1(n253));
   AOI222_X1 U4520 (.ZN(n4260), 
	.C2(n4203), 
	.C1(n3534), 
	.B2(n4240), 
	.B1(n2254), 
	.A2(n4239), 
	.A1(n2196));
   INV_X4 U4521 (.ZN(n1190), 
	.A(n13));
   NOR2_X1 U4522 (.ZN(n13), 
	.A2(n4261), 
	.A1(FE_PHN1037_n5007));
   NAND4_X2 U4524 (.ZN(n2251), 
	.A4(n4265), 
	.A3(n4264), 
	.A2(n4263), 
	.A1(n4262));
   AOI221_X1 U4525 (.ZN(n4265), 
	.C2(vis_r5_o[22]), 
	.C1(n16913), 
	.B2(vis_r4_o[22]), 
	.B1(n16916), 
	.A(n4266));
   OAI222_X1 U4526 (.ZN(n4266), 
	.C2(n16905), 
	.C1(n5465), 
	.B2(n16908), 
	.B1(n5184), 
	.A2(n16910), 
	.A1(n4764));
   AOI221_X1 U4529 (.ZN(n4264), 
	.C2(vis_r10_o[22]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[20]), 
	.B1(n16902), 
	.A(n4267));
   OAI22_X1 U4530 (.ZN(n4267), 
	.B2(n16893), 
	.B1(n5051), 
	.A2(n16895), 
	.A1(n5296));
   AOI221_X1 U4533 (.ZN(n4263), 
	.C2(vis_r12_o[22]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[22]), 
	.B1(FE_OFN638_n16891), 
	.A(n4268));
   OAI22_X1 U4534 (.ZN(n4268), 
	.B2(n16882), 
	.B1(n5407), 
	.A2(n16885), 
	.A1(n5048));
   AOI221_X1 U4537 (.ZN(n4262), 
	.C2(vis_r3_o[22]), 
	.C1(FE_OFN635_n16877), 
	.B2(vis_r0_o[22]), 
	.B1(n4224), 
	.A(n4270));
   OAI22_X1 U4538 (.ZN(n4270), 
	.B2(n16873), 
	.B1(n5320), 
	.A2(n16875), 
	.A1(n5050));
   NAND4_X1 U4541 (.ZN(n4198), 
	.A4(n4271), 
	.A3(n1117), 
	.A2(n1118), 
	.A1(n1112));
   NOR3_X1 U4542 (.ZN(n4271), 
	.A3(hwdata_o[26]), 
	.A2(hwdata_o[29]), 
	.A1(hwdata_o[24]));
   AOI222_X1 U4545 (.ZN(n4272), 
	.C2(n4203), 
	.C1(n1755), 
	.B2(n4240), 
	.B1(n2259), 
	.A2(n4239), 
	.A1(n2556));
   AOI222_X1 U4547 (.ZN(n25), 
	.C2(n4203), 
	.C1(n2496), 
	.B2(n4240), 
	.B1(n2261), 
	.A2(n4239), 
	.A1(n1354));
   NAND4_X2 U4549 (.ZN(n20), 
	.A4(n4276), 
	.A3(n4275), 
	.A2(n4274), 
	.A1(n4273));
   AOI221_X1 U4550 (.ZN(n4276), 
	.C2(vis_r5_o[20]), 
	.C1(n16913), 
	.B2(vis_r4_o[20]), 
	.B1(n16916), 
	.A(n4277));
   OAI222_X1 U4551 (.ZN(n4277), 
	.C2(n16905), 
	.C1(n5604), 
	.B2(n16908), 
	.B1(n5612), 
	.A2(n16910), 
	.A1(n4766));
   AOI221_X1 U4554 (.ZN(n4275), 
	.C2(vis_r10_o[20]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[18]), 
	.B1(n16902), 
	.A(n4278));
   OAI22_X1 U4555 (.ZN(n4278), 
	.B2(n16893), 
	.B1(n5616), 
	.A2(n16895), 
	.A1(n5615));
   AOI221_X1 U4558 (.ZN(n4274), 
	.C2(vis_r12_o[20]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[20]), 
	.B1(FE_OFN638_n16891), 
	.A(n4279));
   OAI22_X1 U4559 (.ZN(n4279), 
	.B2(n16882), 
	.B1(n5606), 
	.A2(n16885), 
	.A1(n5603));
   AOI221_X1 U4562 (.ZN(n4273), 
	.C2(vis_r3_o[20]), 
	.C1(FE_OFN635_n16877), 
	.B2(vis_r0_o[20]), 
	.B1(n4224), 
	.A(n4281));
   OAI22_X1 U4563 (.ZN(n4281), 
	.B2(n16873), 
	.B1(n5609), 
	.A2(n16875), 
	.A1(n5613));
   NAND4_X2 U4567 (.ZN(n17), 
	.A4(n4285), 
	.A3(n4284), 
	.A2(n4283), 
	.A1(n4282));
   AOI221_X1 U4568 (.ZN(n4285), 
	.C2(vis_r5_o[16]), 
	.C1(n16913), 
	.B2(vis_r4_o[16]), 
	.B1(n16916), 
	.A(n4286));
   OAI222_X1 U4569 (.ZN(n4286), 
	.C2(n16905), 
	.C1(n5470), 
	.B2(n16908), 
	.B1(n5189), 
	.A2(n16910), 
	.A1(n4770));
   AOI221_X1 U4572 (.ZN(n4284), 
	.C2(vis_r10_o[16]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[14]), 
	.B1(n16902), 
	.A(n4287));
   OAI22_X1 U4573 (.ZN(n4287), 
	.B2(n16893), 
	.B1(n5072), 
	.A2(n16895), 
	.A1(n5299));
   AOI221_X1 U4576 (.ZN(n4283), 
	.C2(vis_r12_o[16]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[16]), 
	.B1(FE_OFN638_n16891), 
	.A(n4288));
   OAI22_X1 U4577 (.ZN(n4288), 
	.B2(n16882), 
	.B1(n5412), 
	.A2(n16885), 
	.A1(n5069));
   AOI221_X1 U4580 (.ZN(n4282), 
	.C2(vis_r3_o[16]), 
	.C1(FE_OFN635_n16877), 
	.B2(vis_r0_o[16]), 
	.B1(n4224), 
	.A(n4290));
   OAI22_X1 U4581 (.ZN(n4290), 
	.B2(n16873), 
	.B1(n5325), 
	.A2(n16875), 
	.A1(n5071));
   NAND4_X2 U4585 (.ZN(n2258), 
	.A4(n4294), 
	.A3(n4293), 
	.A2(n4292), 
	.A1(n4291));
   AOI221_X1 U4586 (.ZN(n4294), 
	.C2(vis_r5_o[17]), 
	.C1(n16913), 
	.B2(vis_r4_o[17]), 
	.B1(n16916), 
	.A(n4295));
   OAI222_X1 U4587 (.ZN(n4295), 
	.C2(n16905), 
	.C1(n5469), 
	.B2(n16908), 
	.B1(n5188), 
	.A2(n16910), 
	.A1(n4769));
   AOI221_X1 U4590 (.ZN(n4293), 
	.C2(vis_r10_o[17]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[15]), 
	.B1(n16902), 
	.A(n4296));
   OAI22_X1 U4591 (.ZN(n4296), 
	.B2(n16893), 
	.B1(n5086), 
	.A2(n16895), 
	.A1(n5298));
   AOI221_X1 U4594 (.ZN(n4292), 
	.C2(vis_r12_o[17]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[17]), 
	.B1(FE_OFN638_n16891), 
	.A(n4297));
   OAI22_X1 U4595 (.ZN(n4297), 
	.B2(n16882), 
	.B1(n5411), 
	.A2(n16885), 
	.A1(n5083));
   AOI221_X1 U4598 (.ZN(n4291), 
	.C2(vis_r3_o[17]), 
	.C1(FE_OFN635_n16877), 
	.B2(vis_r0_o[17]), 
	.B1(n4224), 
	.A(n4299));
   OAI22_X1 U4599 (.ZN(n4299), 
	.B2(n16873), 
	.B1(n5324), 
	.A2(n16875), 
	.A1(n5085));
   INV_X1 U4602 (.ZN(n4196), 
	.A(n4894));
   AOI21_X1 U4603 (.ZN(n4894), 
	.B2(n17092), 
	.B1(n1398), 
	.A(FE_PHN1348_n4300));
   AOI21_X1 U4604 (.ZN(n4300), 
	.B2(n5527), 
	.B1(FE_PHN2992_IRQ_2_), 
	.A(n4301));
   AOI22_X1 U4605 (.ZN(n4301), 
	.B2(n4192), 
	.B1(hwdata_o[2]), 
	.A2(n5528), 
	.A1(n1396));
   NAND2_X1 U4606 (.ZN(n1396), 
	.A2(n1124), 
	.A1(hwdata_o[2]));
   INV_X1 U4611 (.ZN(n1012), 
	.A(n4302));
   OAI221_X1 U4612 (.ZN(n4302), 
	.C2(n4305), 
	.C1(n559), 
	.B2(n4304), 
	.B1(n4303), 
	.A(n4306));
   OAI21_X1 U4613 (.ZN(n4306), 
	.B2(n4307), 
	.B1(n1866), 
	.A(n5228));
   OAI33_X1 U4614 (.ZN(n4307), 
	.B3(n532), 
	.B2(FE_OFN107_n585), 
	.B1(n4309), 
	.A3(n4308), 
	.A2(n16802), 
	.A1(n4179));
   OR2_X1 U4615 (.ZN(n4309), 
	.A2(n918), 
	.A1(n1856));
   NAND2_X1 U4616 (.ZN(n1856), 
	.A2(n16842), 
	.A1(n16825));
   NAND2_X1 U4617 (.ZN(n4179), 
	.A2(FE_OFN610_n16690), 
	.A1(n1574));
   OAI211_X1 U4618 (.ZN(n1866), 
	.C2(n4310), 
	.C1(n559), 
	.B(n4312), 
	.A(n4311));
   NOR2_X1 U4619 (.ZN(n4312), 
	.A2(n4313), 
	.A1(n1839));
   NOR4_X1 U4620 (.ZN(n4313), 
	.A4(n604), 
	.A3(n1469), 
	.A2(n532), 
	.A1(n4314));
   AOI21_X1 U4621 (.ZN(n1469), 
	.B2(FE_OFN426_n659), 
	.B1(n781), 
	.A(n669));
   NAND2_X1 U4623 (.ZN(n4314), 
	.A2(n466), 
	.A1(n760));
   INV_X1 U4624 (.ZN(n1839), 
	.A(n2658));
   OAI21_X1 U4625 (.ZN(n2658), 
	.B2(n991), 
	.B1(n667), 
	.A(n909));
   INV_X4 U4626 (.ZN(n909), 
	.A(n1541));
   NAND2_X1 U4627 (.ZN(n1541), 
	.A2(n16808), 
	.A1(FE_OFN73_n16806));
   NAND3_X1 U4628 (.ZN(n4311), 
	.A3(n4316), 
	.A2(n16826), 
	.A1(n4315));
   INV_X1 U4629 (.ZN(n4316), 
	.A(n4308));
   NAND3_X1 U4630 (.ZN(n4308), 
	.A3(n501), 
	.A2(n1094), 
	.A1(n592));
   OAI21_X1 U4631 (.ZN(n4315), 
	.B2(n603), 
	.B1(n16725), 
	.A(n2673));
   NOR2_X1 U4632 (.ZN(n2673), 
	.A2(n475), 
	.A1(n602));
   OAI21_X1 U4633 (.ZN(n602), 
	.B2(n16659), 
	.B1(n16802), 
	.A(n711));
   NAND2_X1 U4634 (.ZN(n711), 
	.A2(n16725), 
	.A1(n16804));
   NAND2_X1 U4635 (.ZN(n603), 
	.A2(n16802), 
	.A1(n4974));
   INV_X1 U4636 (.ZN(n559), 
	.A(n930));
   NAND2_X1 U4637 (.ZN(n4304), 
	.A2(n16808), 
	.A1(n17096));
   AOI22_X1 U4639 (.ZN(n4303), 
	.B2(FE_OFN19_n1063), 
	.B1(n5228), 
	.A2(n4317), 
	.A1(n5167));
   NAND2_X1 U4640 (.ZN(n4317), 
	.A2(n1343), 
	.A1(n1040));
   INV_X1 U4641 (.ZN(n1343), 
	.A(n181));
   INV_X1 U4642 (.ZN(n1040), 
	.A(n1058));
   NAND4_X1 U4643 (.ZN(n1058), 
	.A4(n4320), 
	.A3(n4319), 
	.A2(n1860), 
	.A1(n4318));
   AOI22_X1 U4644 (.ZN(n4320), 
	.B2(n529), 
	.B1(n528), 
	.A2(n16862), 
	.A1(n1173));
   INV_X1 U4645 (.ZN(n528), 
	.A(n692));
   AND3_X1 U4646 (.ZN(n1173), 
	.A3(FE_OFN469_n1034), 
	.A2(FE_OFN627_n16828), 
	.A1(n563));
   NOR2_X1 U4647 (.ZN(n1034), 
	.A2(FE_OFN85_n16839), 
	.A1(n16826));
   NAND4_X1 U4648 (.ZN(n4319), 
	.A4(FE_OFN81_n16856), 
	.A3(n16821), 
	.A2(n760), 
	.A1(n809));
   INV_X1 U4649 (.ZN(n1860), 
	.A(n1473));
   NOR3_X1 U4650 (.ZN(n1473), 
	.A3(FE_OFN422_n641), 
	.A2(n5165), 
	.A1(n745));
   INV_X1 U4651 (.ZN(n4186), 
	.A(n4321));
   AOI221_X1 U4652 (.ZN(n4321), 
	.C2(n4749), 
	.C1(n4900), 
	.B2(n5572), 
	.B1(n11971), 
	.A(n4322));
   INV_X1 U4653 (.ZN(n4322), 
	.A(n4323));
   AOI222_X1 U4654 (.ZN(n4323), 
	.C2(n5533), 
	.C1(n11945), 
	.B2(n5534), 
	.B1(n11939), 
	.A2(n11957), 
	.A1(n5011));
   AOI21_X1 U4655 (.ZN(n11945), 
	.B2(n17092), 
	.B1(n1419), 
	.A(FE_PHN1900_n4324));
   AOI21_X1 U4656 (.ZN(n4324), 
	.B2(FE_PHN2984_IRQ_5_), 
	.B1(n1411), 
	.A(n4325));
   AOI22_X1 U4657 (.ZN(n4325), 
	.B2(n4192), 
	.B1(hwdata_o[5]), 
	.A2(n5533), 
	.A1(n1416));
   NAND2_X1 U4658 (.ZN(n1416), 
	.A2(n1124), 
	.A1(hwdata_o[5]));
   AOI21_X1 U4662 (.ZN(n11939), 
	.B2(n17092), 
	.B1(n1453), 
	.A(FE_PHN1899_n4326));
   AOI21_X1 U4663 (.ZN(n4326), 
	.B2(FE_PHN4634_IRQ_1_), 
	.B1(n1447), 
	.A(n4327));
   AOI22_X1 U4664 (.ZN(n4327), 
	.B2(n4192), 
	.B1(hwdata_o[1]), 
	.A2(n5534), 
	.A1(n1452));
   NAND2_X1 U4665 (.ZN(n1452), 
	.A2(n1124), 
	.A1(hwdata_o[1]));
   NOR2_X1 U4669 (.ZN(n11957), 
	.A2(n1128), 
	.A1(FE_PHN1598_n4328));
   NOR2_X1 U4670 (.ZN(n1128), 
	.A2(n4329), 
	.A1(n200));
   AOI221_X1 U4671 (.ZN(n4328), 
	.C2(FE_PHN4637_IRQ_9_), 
	.C1(n5580), 
	.B2(n1124), 
	.B1(hwdata_o[9]), 
	.A(n4330));
   AOI21_X1 U4672 (.ZN(n4330), 
	.B2(n4192), 
	.B1(hwdata_o[9]), 
	.A(n5011));
   AOI21_X1 U4673 (.ZN(n4900), 
	.B2(n17092), 
	.B1(n1446), 
	.A(FE_PHN1512_n4331));
   INV_X1 U4674 (.ZN(n4331), 
	.A(n4332));
   OAI221_X1 U4675 (.ZN(n4332), 
	.C2(n4333), 
	.C1(FE_PHN2970_n1444), 
	.B2(n1385), 
	.B1(n240), 
	.A(n4334));
   OAI21_X1 U4676 (.ZN(n4334), 
	.B2(n4335), 
	.B1(n240), 
	.A(n3089));
   INV_X1 U4679 (.ZN(n1444), 
	.A(irq_i[12]));
   NOR2_X1 U4680 (.ZN(n11971), 
	.A2(n1432), 
	.A1(FE_PHN1356_n4336));
   NOR2_X1 U4681 (.ZN(n1432), 
	.A2(n4337), 
	.A1(n200));
   AOI221_X1 U4682 (.ZN(n4336), 
	.C2(FE_PHN5177_IRQ_11_), 
	.C1(n4338), 
	.B2(n1124), 
	.B1(hwdata_o[11]), 
	.A(n4339));
   AOI21_X1 U4683 (.ZN(n4339), 
	.B2(n4192), 
	.B1(hwdata_o[11]), 
	.A(n5572));
   NAND4_X1 U4685 (.ZN(n4185), 
	.A4(n4343), 
	.A3(n4342), 
	.A2(n4341), 
	.A1(n4340));
   AOI21_X1 U4686 (.ZN(n4343), 
	.B2(n4344), 
	.B1(n4748), 
	.A(n4345));
   OAI33_X1 U4687 (.ZN(n4345), 
	.B3(n930), 
	.B2(n1050), 
	.B1(n1053), 
	.A3(n209), 
	.A2(n205), 
	.A1(n202));
   OAI211_X1 U4688 (.ZN(n930), 
	.C2(n4347), 
	.C1(n4346), 
	.B(n1045), 
	.A(n181));
   NAND4_X1 U4690 (.ZN(n181), 
	.A4(n170), 
	.A3(n4348), 
	.A2(n176), 
	.A1(vis_ipsr_o[1]));
   AOI22_X1 U4691 (.ZN(n4347), 
	.B2(n4350), 
	.B1(n1355), 
	.A2(n3732), 
	.A1(n4349));
   OR2_X1 U4692 (.ZN(n4349), 
	.A2(n1355), 
	.A1(n4350));
   NOR4_X1 U4693 (.ZN(n1355), 
	.A4(n4354), 
	.A3(n4353), 
	.A2(n4352), 
	.A1(n4351));
   OAI221_X1 U4694 (.ZN(n4354), 
	.C2(n199), 
	.C1(n5098), 
	.B2(n1456), 
	.B1(n5153), 
	.A(n4355));
   AOI222_X1 U4695 (.ZN(n4355), 
	.C2(n3862), 
	.C1(n1404), 
	.B2(n4356), 
	.B1(n1386), 
	.A2(n3791), 
	.A1(n1378));
   OAI221_X1 U4699 (.ZN(n4353), 
	.C2(n1451), 
	.C1(n5547), 
	.B2(n1415), 
	.B1(n5023), 
	.A(n4357));
   AOI222_X1 U4700 (.ZN(n4357), 
	.C2(n3792), 
	.C1(n1430), 
	.B2(n3732), 
	.B1(n4358), 
	.A2(n3793), 
	.A1(n1122));
   OAI221_X1 U4704 (.ZN(n4352), 
	.C2(n1423), 
	.C1(n5523), 
	.B2(n1441), 
	.B1(n5522), 
	.A(n4359));
   AOI22_X1 U4705 (.ZN(n4359), 
	.B2(n3833), 
	.B1(n1392), 
	.A2(n3847), 
	.A1(n1318));
   INV_X1 U4707 (.ZN(n1392), 
	.A(n1391));
   OAI221_X1 U4709 (.ZN(n4351), 
	.C2(n207), 
	.C1(n4961), 
	.B2(n1397), 
	.B1(n5551), 
	.A(n4360));
   AOI222_X1 U4710 (.ZN(n4360), 
	.C2(n3813), 
	.C1(n1126), 
	.B2(n3784), 
	.B1(n1446), 
	.A2(n3863), 
	.A1(n1410));
   INV_X1 U4712 (.ZN(n1126), 
	.A(n4329));
   INV_X1 U4714 (.ZN(n1446), 
	.A(n1445));
   NAND2_X1 U4716 (.ZN(n4350), 
	.A2(n4361), 
	.A1(n5503));
   NAND4_X1 U4717 (.ZN(n4361), 
	.A4(n1367), 
	.A3(n1365), 
	.A2(n1363), 
	.A1(n1362));
   AOI221_X1 U4718 (.ZN(n1367), 
	.C2(n1122), 
	.C1(n2888), 
	.B2(n1404), 
	.B1(n2931), 
	.A(n4362));
   OAI22_X1 U4719 (.ZN(n4362), 
	.B2(n5151), 
	.B1(n1384), 
	.A2(n5160), 
	.A1(n4337));
   INV_X1 U4722 (.ZN(n1365), 
	.A(n4363));
   OAI221_X1 U4723 (.ZN(n4363), 
	.C2(n1885), 
	.C1(n1445), 
	.B2(n1456), 
	.B1(n5152), 
	.A(n4364));
   AOI222_X1 U4724 (.ZN(n4364), 
	.C2(n2889), 
	.C1(n4366), 
	.B2(n2929), 
	.B1(n4365), 
	.A2(n2927), 
	.A1(n1378));
   AOI221_X1 U4729 (.ZN(n1363), 
	.C2(n1419), 
	.C1(n2902), 
	.B2(n1410), 
	.B1(n4367), 
	.A(n4368));
   OAI222_X1 U4730 (.ZN(n4368), 
	.C2(n5157), 
	.C1(n4329), 
	.B2(n5518), 
	.B1(n1441), 
	.A2(n5519), 
	.A1(n1423));
   INV_X1 U4731 (.ZN(n1419), 
	.A(n1415));
   AOI221_X1 U4734 (.ZN(n1362), 
	.C2(n1318), 
	.C1(n2951), 
	.B2(n4752), 
	.B1(n1398), 
	.A(n4369));
   OAI22_X1 U4735 (.ZN(n4369), 
	.B2(n5552), 
	.B1(n1391), 
	.A2(n5550), 
	.A1(n1451));
   INV_X1 U4737 (.ZN(n4346), 
	.A(n1358));
   NAND4_X1 U4738 (.ZN(n1358), 
	.A4(n4373), 
	.A3(n4372), 
	.A2(n4371), 
	.A1(n4370));
   NOR4_X1 U4739 (.ZN(n4373), 
	.A4(n4365), 
	.A3(n4366), 
	.A2(n1453), 
	.A1(n4374));
   INV_X1 U4740 (.ZN(n4365), 
	.A(n199));
   NAND2_X1 U4741 (.ZN(n199), 
	.A2(n4376), 
	.A1(n4375));
   INV_X1 U4742 (.ZN(n4366), 
	.A(n207));
   NAND2_X1 U4743 (.ZN(n207), 
	.A2(n4376), 
	.A1(n4377));
   INV_X1 U4744 (.ZN(n1453), 
	.A(n1451));
   NAND2_X1 U4745 (.ZN(n1451), 
	.A2(n4379), 
	.A1(n4378));
   NAND2_X1 U4746 (.ZN(n4374), 
	.A2(n1415), 
	.A1(n1391));
   NAND2_X1 U4747 (.ZN(n1415), 
	.A2(n4375), 
	.A1(n4379));
   NAND2_X1 U4748 (.ZN(n1391), 
	.A2(n4378), 
	.A1(n4380));
   NOR4_X1 U4749 (.ZN(n4372), 
	.A4(n1398), 
	.A3(n1318), 
	.A2(n1410), 
	.A1(n4381));
   INV_X1 U4750 (.ZN(n1398), 
	.A(n1397));
   NAND2_X1 U4751 (.ZN(n1397), 
	.A2(n4380), 
	.A1(n4382));
   INV_X1 U4752 (.ZN(n1318), 
	.A(n1315));
   NAND2_X1 U4753 (.ZN(n1315), 
	.A2(n4379), 
	.A1(n4382));
   NAND2_X1 U4754 (.ZN(n4381), 
	.A2(n1423), 
	.A1(n4329));
   NAND2_X1 U4755 (.ZN(n4329), 
	.A2(n4378), 
	.A1(n4383));
   NOR3_X1 U4756 (.ZN(n4371), 
	.A3(n1122), 
	.A2(n1378), 
	.A1(n4384));
   INV_X1 U4757 (.ZN(n1122), 
	.A(n1436));
   NAND2_X1 U4758 (.ZN(n1436), 
	.A2(n4382), 
	.A1(n4385));
   NAND3_X1 U4759 (.ZN(n4384), 
	.A3(n1456), 
	.A2(n1441), 
	.A1(n1445));
   NAND2_X1 U4760 (.ZN(n1441), 
	.A2(n4382), 
	.A1(n4383));
   NAND2_X1 U4761 (.ZN(n1445), 
	.A2(n4377), 
	.A1(n4383));
   NOR4_X1 U4762 (.ZN(n4370), 
	.A4(n4358), 
	.A3(n1430), 
	.A2(n1386), 
	.A1(n1404));
   INV_X1 U4763 (.ZN(n4358), 
	.A(n1052));
   NAND2_X1 U4764 (.ZN(n1052), 
	.A2(n4376), 
	.A1(n4378));
   NOR4_X1 U4765 (.ZN(n4376), 
	.A4(vis_ipsr_o[5]), 
	.A3(vis_ipsr_o[4]), 
	.A2(n191), 
	.A1(n170));
   INV_X1 U4766 (.ZN(n1430), 
	.A(n4337));
   NAND2_X1 U4767 (.ZN(n4337), 
	.A2(n4378), 
	.A1(n4385));
   NOR2_X1 U4768 (.ZN(n4378), 
	.A2(vis_ipsr_o[2]), 
	.A1(n186));
   AND2_X1 U4769 (.ZN(n1050), 
	.A2(n4310), 
	.A1(n4305));
   NAND3_X1 U4770 (.ZN(n4310), 
	.A3(n542), 
	.A2(n914), 
	.A1(n827));
   NOR2_X1 U4771 (.ZN(n542), 
	.A2(FE_OFN81_n16856), 
	.A1(n16842));
   INV_X1 U4772 (.ZN(n914), 
	.A(n762));
   NAND2_X1 U4773 (.ZN(n762), 
	.A2(n16870), 
	.A1(FE_OFN73_n16806));
   NAND4_X1 U4775 (.ZN(n4305), 
	.A4(n3509), 
	.A3(n16820), 
	.A2(n16824), 
	.A1(n563));
   INV_X1 U4776 (.ZN(n3509), 
	.A(n1088));
   NAND3_X1 U4777 (.ZN(n1088), 
	.A3(n16862), 
	.A2(n1574), 
	.A1(n991));
   NAND2_X2 U4781 (.ZN(n1234), 
	.A2(n16694), 
	.A1(n16845));
   AOI222_X1 U4784 (.ZN(n205), 
	.C2(n4203), 
	.C1(n89), 
	.B2(n4240), 
	.B1(n2247), 
	.A2(n4239), 
	.A1(n2578));
   INV_X1 U4785 (.ZN(n4344), 
	.A(n1123));
   AOI221_X1 U4786 (.ZN(n1123), 
	.C2(n5061), 
	.C1(FE_PHN2989_IRQ_10_), 
	.B2(n1124), 
	.B1(hwdata_o[10]), 
	.A(n4386));
   AOI21_X1 U4787 (.ZN(n4386), 
	.B2(n4192), 
	.B1(hwdata_o[10]), 
	.A(n4748));
   AOI222_X1 U4788 (.ZN(n4342), 
	.C2(n4387), 
	.C1(n4747), 
	.B2(n5530), 
	.B1(n4899), 
	.A2(n5532), 
	.A1(n4898));
   INV_X1 U4789 (.ZN(n4387), 
	.A(n1121));
   AOI221_X1 U4790 (.ZN(n1121), 
	.C2(n5582), 
	.C1(FE_PHN2995_IRQ_8_), 
	.B2(n1124), 
	.B1(hwdata_o[8]), 
	.A(n4388));
   AOI21_X1 U4791 (.ZN(n4388), 
	.B2(n4192), 
	.B1(hwdata_o[8]), 
	.A(n4747));
   AOI21_X1 U4792 (.ZN(n4899), 
	.B2(n17092), 
	.B1(n1404), 
	.A(FE_PHN1668_n4389));
   AOI21_X1 U4793 (.ZN(n4389), 
	.B2(n5529), 
	.B1(FE_PHN2990_IRQ_7_), 
	.A(n4390));
   AOI22_X1 U4794 (.ZN(n4390), 
	.B2(n4192), 
	.B1(hwdata_o[7]), 
	.A2(n5530), 
	.A1(n1403));
   NAND2_X1 U4795 (.ZN(n1403), 
	.A2(n1124), 
	.A1(hwdata_o[7]));
   INV_X1 U4798 (.ZN(n1404), 
	.A(n1402));
   NAND2_X1 U4799 (.ZN(n1402), 
	.A2(n4375), 
	.A1(n4380));
   AOI21_X1 U4800 (.ZN(n4898), 
	.B2(n17092), 
	.B1(n1410), 
	.A(FE_PHN1352_n4391));
   AOI21_X1 U4801 (.ZN(n4391), 
	.B2(n5531), 
	.B1(FE_PHN2987_IRQ_6_), 
	.A(n4392));
   AOI22_X1 U4802 (.ZN(n4392), 
	.B2(n4192), 
	.B1(hwdata_o[6]), 
	.A2(n5532), 
	.A1(n1409));
   NAND2_X1 U4803 (.ZN(n1409), 
	.A2(n1124), 
	.A1(hwdata_o[6]));
   INV_X1 U4806 (.ZN(n1410), 
	.A(n1408));
   NAND2_X1 U4807 (.ZN(n1408), 
	.A2(n4377), 
	.A1(n4380));
   AND2_X1 U4808 (.ZN(n4380), 
	.A2(vis_ipsr_o[1]), 
	.A1(n4393));
   AOI222_X1 U4809 (.ZN(n4341), 
	.C2(n3775), 
	.C1(n4897), 
	.B2(n4750), 
	.B1(n4901), 
	.A2(n4896), 
	.A1(n5047));
   AOI21_X1 U4810 (.ZN(n4897), 
	.B2(n17092), 
	.B1(n1386), 
	.A(FE_PHN1358_n4394));
   AOI221_X1 U4811 (.ZN(n4394), 
	.C2(n5118), 
	.C1(FE_PHN2993_IRQ_13_), 
	.B2(n1124), 
	.B1(hwdata_o[13]), 
	.A(n4395));
   AOI21_X1 U4812 (.ZN(n4395), 
	.B2(n4192), 
	.B1(hwdata_o[13]), 
	.A(n3775));
   INV_X1 U4814 (.ZN(n1386), 
	.A(n1384));
   NAND2_X1 U4815 (.ZN(n1384), 
	.A2(n4375), 
	.A1(n4383));
   AND2_X1 U4816 (.ZN(n4383), 
	.A2(n191), 
	.A1(n4396));
   AOI21_X1 U4817 (.ZN(n4901), 
	.B2(n17092), 
	.B1(n1425), 
	.A(FE_PHN1362_n4397));
   AOI21_X1 U4818 (.ZN(n4397), 
	.B2(n5524), 
	.B1(FE_PHN2986_IRQ_4_), 
	.A(n4398));
   AOI22_X1 U4819 (.ZN(n4398), 
	.B2(n4750), 
	.B1(n1424), 
	.A2(n4192), 
	.A1(hwdata_o[4]));
   NAND2_X1 U4820 (.ZN(n1424), 
	.A2(n1124), 
	.A1(hwdata_o[4]));
   INV_X1 U4823 (.ZN(n1425), 
	.A(n1423));
   NAND2_X1 U4824 (.ZN(n1423), 
	.A2(n4377), 
	.A1(n4379));
   AND2_X1 U4825 (.ZN(n4379), 
	.A2(n191), 
	.A1(n4393));
   NOR3_X1 U4826 (.ZN(n4393), 
	.A3(n165), 
	.A2(vis_ipsr_o[5]), 
	.A1(vis_ipsr_o[3]));
   AOI21_X1 U4827 (.ZN(n4896), 
	.B2(n17092), 
	.B1(n1459), 
	.A(n4399));
   AOI221_X1 U4828 (.ZN(n4399), 
	.C2(n5619), 
	.C1(FE_PHN4641_IRQ_14_), 
	.B2(hwdata_o[14]), 
	.B1(n1124), 
	.A(n4400));
   AOI21_X1 U4829 (.ZN(n4400), 
	.B2(n4192), 
	.B1(hwdata_o[14]), 
	.A(n5047));
   NAND4_X1 U4832 (.ZN(n2253), 
	.A4(n4405), 
	.A3(n4404), 
	.A2(n4403), 
	.A1(n4402));
   AOI221_X1 U4833 (.ZN(n4405), 
	.C2(vis_r5_o[14]), 
	.C1(n16913), 
	.B2(vis_r4_o[14]), 
	.B1(n16916), 
	.A(n4406));
   OAI222_X1 U4834 (.ZN(n4406), 
	.C2(n16905), 
	.C1(n5471), 
	.B2(n16908), 
	.B1(n5190), 
	.A2(n16910), 
	.A1(n4850));
   AOI221_X1 U4837 (.ZN(n4404), 
	.C2(vis_r10_o[14]), 
	.C1(n16897), 
	.B2(vis_psp_o[12]), 
	.B1(n16902), 
	.A(n4407));
   OAI22_X1 U4838 (.ZN(n4407), 
	.B2(n16893), 
	.B1(n5106), 
	.A2(n16895), 
	.A1(n5300));
   AOI221_X1 U4841 (.ZN(n4403), 
	.C2(vis_r12_o[14]), 
	.C1(n16886), 
	.B2(vis_r9_o[14]), 
	.B1(n16891), 
	.A(n4408));
   OAI22_X1 U4842 (.ZN(n4408), 
	.B2(n16882), 
	.B1(n5413), 
	.A2(n16885), 
	.A1(n5103));
   AOI221_X1 U4845 (.ZN(n4402), 
	.C2(vis_r3_o[14]), 
	.C1(n16877), 
	.B2(vis_r0_o[14]), 
	.B1(n4224), 
	.A(n4410));
   OAI22_X1 U4846 (.ZN(n4410), 
	.B2(n16873), 
	.B1(n5326), 
	.A2(n16875), 
	.A1(n5105));
   NAND4_X2 U4849 (.ZN(n2250), 
	.A4(n4414), 
	.A3(n4413), 
	.A2(n4412), 
	.A1(n4411));
   AOI222_X1 U4850 (.ZN(n4414), 
	.C2(vis_msp_o[4]), 
	.C1(n16651), 
	.B2(n1152), 
	.B1(n16911), 
	.A2(vis_r14_o[6]), 
	.A1(n16652));
   AOI22_X1 U4854 (.ZN(n4413), 
	.B2(vis_r10_o[6]), 
	.B1(n16897), 
	.A2(vis_psp_o[4]), 
	.A1(n16902));
   AOI222_X1 U4857 (.ZN(n4412), 
	.C2(vis_r9_o[6]), 
	.C1(n16891), 
	.B2(vis_r8_o[6]), 
	.B1(n16648), 
	.A2(vis_r12_o[6]), 
	.A1(n16886));
   AOI21_X1 U4861 (.ZN(n4411), 
	.B2(vis_r11_o[6]), 
	.B1(n16650), 
	.A(n1794));
   NAND2_X1 U4862 (.ZN(n1794), 
	.A2(n4421), 
	.A1(n4420));
   AOI221_X1 U4863 (.ZN(n4421), 
	.C2(vis_r5_o[6]), 
	.C1(FE_OFN642_n16913), 
	.B2(vis_r4_o[6]), 
	.B1(FE_OFN643_n16916), 
	.A(n4422));
   OAI22_X1 U4864 (.ZN(n4422), 
	.B2(n16908), 
	.B1(n5180), 
	.A2(n16905), 
	.A1(n5461));
   AOI221_X1 U4867 (.ZN(n4420), 
	.C2(vis_r7_o[6]), 
	.C1(n16649), 
	.B2(vis_r3_o[6]), 
	.B1(n16877), 
	.A(n4426));
   OAI22_X1 U4868 (.ZN(n4426), 
	.B2(n16885), 
	.B1(n5041), 
	.A2(n4427), 
	.A1(n5485));
   INV_X1 U4872 (.ZN(n1459), 
	.A(n1456));
   NAND2_X1 U4873 (.ZN(n1456), 
	.A2(n4377), 
	.A1(n4385));
   NOR2_X1 U4874 (.ZN(n4377), 
	.A2(vis_ipsr_o[0]), 
	.A1(n176));
   AOI22_X1 U4875 (.ZN(n4340), 
	.B2(n204), 
	.B1(n4988), 
	.A2(FE_PHN1367_n4895), 
	.A1(n5024));
   OAI21_X1 U4876 (.ZN(n204), 
	.B2(n202), 
	.B1(n24), 
	.A(n4428));
   OR4_X1 U4877 (.ZN(n4428), 
	.A4(n4833), 
	.A3(FE_PHN3501_n5516), 
	.A2(n260), 
	.A1(n259));
   NAND4_X1 U4879 (.ZN(n259), 
	.A4(n4432), 
	.A3(n4431), 
	.A2(n4430), 
	.A1(n4429));
   NOR4_X1 U4880 (.ZN(n4432), 
	.A4(sub_2068_A_5_), 
	.A3(sub_2068_A_6_), 
	.A2(sub_2068_A_4_), 
	.A1(n4433));
   NAND3_X1 U4881 (.ZN(n4433), 
	.A3(n298), 
	.A2(n294), 
	.A1(n296));
   NOR4_X1 U4885 (.ZN(n4431), 
	.A4(sub_2068_A_21_), 
	.A3(sub_2068_A_22_), 
	.A2(sub_2068_A_20_), 
	.A1(n4434));
   NAND3_X1 U4886 (.ZN(n4434), 
	.A3(n264), 
	.A2(n306), 
	.A1(n308));
   NOR4_X1 U4890 (.ZN(n4430), 
	.A4(sub_2068_A_16_), 
	.A3(sub_2068_A_17_), 
	.A2(sub_2068_A_15_), 
	.A1(n4435));
   NAND3_X1 U4891 (.ZN(n4435), 
	.A3(n276), 
	.A2(n310), 
	.A1(n274));
   NOR3_X1 U4895 (.ZN(n4429), 
	.A3(sub_2068_A_10_), 
	.A2(sub_2068_A_11_), 
	.A1(n4436));
   NAND3_X1 U4896 (.ZN(n4436), 
	.A3(n288), 
	.A2(n284), 
	.A1(n286));
   OR2_X1 U4900 (.ZN(n202), 
	.A2(FE_PHN1037_n5007), 
	.A1(n3962));
   NAND3_X1 U4901 (.ZN(n3962), 
	.A3(n3717), 
	.A2(n251), 
	.A1(n5017));
   NOR3_X1 U4902 (.ZN(n3717), 
	.A3(n3874), 
	.A2(FE_PHN1894_n5149), 
	.A1(n5502));
   AOI222_X1 U4904 (.ZN(n24), 
	.C2(n4239), 
	.C1(n3177), 
	.B2(n4203), 
	.B1(n2260), 
	.A2(n4240), 
	.A1(n3145));
   NAND4_X1 U4905 (.ZN(n2260), 
	.A4(n4440), 
	.A3(n4439), 
	.A2(n4438), 
	.A1(n4437));
   AOI221_X1 U4906 (.ZN(n4440), 
	.C2(vis_r5_o[26]), 
	.C1(n16913), 
	.B2(vis_r4_o[26]), 
	.B1(n16916), 
	.A(n4441));
   OAI222_X1 U4907 (.ZN(n4441), 
	.C2(n16905), 
	.C1(n5458), 
	.B2(n16908), 
	.B1(n5177), 
	.A2(n16910), 
	.A1(n4762));
   AOI221_X1 U4910 (.ZN(n4439), 
	.C2(vis_r10_o[26]), 
	.C1(n16897), 
	.B2(vis_psp_o[24]), 
	.B1(n16902), 
	.A(n4442));
   OAI22_X1 U4911 (.ZN(n4442), 
	.B2(n16893), 
	.B1(n4992), 
	.A2(n16895), 
	.A1(n5290));
   AOI221_X1 U4914 (.ZN(n4438), 
	.C2(vis_r12_o[26]), 
	.C1(n16886), 
	.B2(vis_r9_o[26]), 
	.B1(n16891), 
	.A(n4443));
   OAI22_X1 U4915 (.ZN(n4443), 
	.B2(n16882), 
	.B1(n5400), 
	.A2(n16885), 
	.A1(n4989));
   AOI221_X1 U4918 (.ZN(n4437), 
	.C2(vis_r3_o[26]), 
	.C1(n16877), 
	.B2(vis_r0_o[26]), 
	.B1(n4224), 
	.A(n4445));
   OAI22_X1 U4919 (.ZN(n4445), 
	.B2(n16873), 
	.B1(n5313), 
	.A2(n16875), 
	.A1(n4991));
   INV_X1 U4923 (.ZN(n1614), 
	.A(n1670));
   AOI21_X1 U4924 (.ZN(n4895), 
	.B2(n17092), 
	.B1(n1378), 
	.A(n4446));
   AOI221_X1 U4925 (.ZN(n4446), 
	.C2(n5620), 
	.C1(FE_PHN5178_IRQ_15_), 
	.B2(hwdata_o[15]), 
	.B1(n1124), 
	.A(n4447));
   AOI21_X1 U4926 (.ZN(n4447), 
	.B2(n4192), 
	.B1(hwdata_o[15]), 
	.A(n5024));
   NAND3_X1 U4928 (.ZN(n4335), 
	.A3(n3873), 
	.A2(n253), 
	.A1(n1385));
   NAND4_X2 U4931 (.ZN(n2254), 
	.A4(n4451), 
	.A3(n4450), 
	.A2(n4449), 
	.A1(n4448));
   AOI221_X1 U4932 (.ZN(n4451), 
	.C2(vis_r5_o[15]), 
	.C1(n16913), 
	.B2(vis_r4_o[15]), 
	.B1(n16916), 
	.A(n4452));
   OAI222_X1 U4933 (.ZN(n4452), 
	.C2(n16905), 
	.C1(n5478), 
	.B2(n16908), 
	.B1(n5197), 
	.A2(n16910), 
	.A1(n4827));
   AOI221_X1 U4936 (.ZN(n4450), 
	.C2(vis_r10_o[15]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[13]), 
	.B1(FE_OFN641_n16902), 
	.A(n4453));
   OAI22_X1 U4937 (.ZN(n4453), 
	.B2(n16893), 
	.B1(n5633), 
	.A2(n16895), 
	.A1(n5632));
   AOI221_X1 U4940 (.ZN(n4449), 
	.C2(vis_r12_o[15]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[15]), 
	.B1(FE_OFN638_n16891), 
	.A(n4454));
   OAI22_X1 U4941 (.ZN(n4454), 
	.B2(n16882), 
	.B1(n5420), 
	.A2(n16885), 
	.A1(n5108));
   AOI221_X1 U4944 (.ZN(n4448), 
	.C2(vis_r3_o[15]), 
	.C1(FE_OFN635_n16877), 
	.B2(vis_r0_o[15]), 
	.B1(n4224), 
	.A(n4456));
   OAI22_X1 U4945 (.ZN(n4456), 
	.B2(n16873), 
	.B1(n5333), 
	.A2(n16875), 
	.A1(n5110));
   NAND3_X1 U4949 (.ZN(n1385), 
	.A3(n3873), 
	.A2(n253), 
	.A1(n4905));
   NOR4_X1 U4950 (.ZN(n3873), 
	.A4(n5017), 
	.A3(n5502), 
	.A2(n1110), 
	.A1(n3874));
   INV_X4 U4956 (.ZN(n760), 
	.A(n568));
   INV_X4 U4957 (.ZN(n809), 
	.A(n813));
   NAND2_X1 U4958 (.ZN(n813), 
	.A2(n16831), 
	.A1(n608));
   AND2_X1 U4959 (.ZN(n1378), 
	.A2(n4375), 
	.A1(n4385));
   NOR2_X1 U4960 (.ZN(n4375), 
	.A2(n176), 
	.A1(n186));
   AND2_X1 U4963 (.ZN(n4385), 
	.A2(vis_ipsr_o[1]), 
	.A1(n4396));
   NOR3_X1 U4964 (.ZN(n4396), 
	.A3(n165), 
	.A2(vis_ipsr_o[5]), 
	.A1(n170));
   NOR4_X1 U4966 (.ZN(n4181), 
	.A4(n1583), 
	.A3(FE_OFN629_n16850), 
	.A2(n1784), 
	.A1(n4457));
   NOR3_X1 U4967 (.ZN(n1583), 
	.A3(n604), 
	.A2(n16821), 
	.A1(n16871));
   NAND2_X1 U4968 (.ZN(n4457), 
	.A2(n2661), 
	.A1(n1097));
   INV_X1 U4969 (.ZN(n2661), 
	.A(n849));
   INV_X1 U4970 (.ZN(n1097), 
	.A(n989));
   NAND2_X2 U4971 (.ZN(n989), 
	.A2(FE_OFN79_n16834), 
	.A1(n997));
   NAND4_X2 U4974 (.ZN(n2261), 
	.A4(n4461), 
	.A3(n4460), 
	.A2(n4459), 
	.A1(n4458));
   AOI221_X1 U4975 (.ZN(n4461), 
	.C2(vis_r5_o[8]), 
	.C1(n16913), 
	.B2(vis_r4_o[8]), 
	.B1(n16916), 
	.A(n4462));
   OAI222_X1 U4976 (.ZN(n4462), 
	.C2(n16905), 
	.C1(n5477), 
	.B2(n16908), 
	.B1(n5196), 
	.A2(n16910), 
	.A1(n4851));
   AOI221_X1 U4979 (.ZN(n4460), 
	.C2(vis_r10_o[8]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[6]), 
	.B1(n16902), 
	.A(n4463));
   OAI22_X1 U4980 (.ZN(n4463), 
	.B2(n16893), 
	.B1(n5138), 
	.A2(n16895), 
	.A1(n5304));
   AOI221_X1 U4983 (.ZN(n4459), 
	.C2(vis_r12_o[8]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[8]), 
	.B1(FE_OFN638_n16891), 
	.A(n4464));
   OAI22_X1 U4984 (.ZN(n4464), 
	.B2(n16882), 
	.B1(n5419), 
	.A2(n16885), 
	.A1(n5135));
   AOI221_X1 U4987 (.ZN(n4458), 
	.C2(vis_r3_o[8]), 
	.C1(FE_OFN635_n16877), 
	.B2(vis_r0_o[8]), 
	.B1(n4224), 
	.A(n4466));
   OAI22_X1 U4988 (.ZN(n4466), 
	.B2(n16873), 
	.B1(n5332), 
	.A2(n16875), 
	.A1(n5137));
   NAND4_X2 U4991 (.ZN(n1354), 
	.A4(n4469), 
	.A3(n4468), 
	.A2(n4467), 
	.A1(n4170));
   AOI221_X1 U4992 (.ZN(n4469), 
	.C2(vis_r8_o[0]), 
	.C1(n16648), 
	.B2(vis_r10_o[0]), 
	.B1(n16897), 
	.A(n4472));
   OAI22_X1 U4993 (.ZN(n4472), 
	.B2(n4211), 
	.B1(n5101), 
	.A2(n16895), 
	.A1(n5288));
   AOI22_X1 U4996 (.ZN(n4468), 
	.B2(vis_r12_o[0]), 
	.B1(n16886), 
	.A2(vis_r9_o[0]), 
	.A1(n16891));
   NAND2_X1 U4999 (.ZN(n4467), 
	.A2(vis_r11_o[0]), 
	.A1(n16650));
   AND2_X4 U5001 (.ZN(n4170), 
	.A2(n4475), 
	.A1(n4474));
   AOI221_X1 U5002 (.ZN(n4475), 
	.C2(vis_r5_o[0]), 
	.C1(n16913), 
	.B2(vis_r4_o[0]), 
	.B1(n16916), 
	.A(n4476));
   OAI22_X2 U5003 (.ZN(n4476), 
	.B2(n16908), 
	.B1(n5173), 
	.A2(n16905), 
	.A1(n5454));
   AOI221_X2 U5006 (.ZN(n4474), 
	.C2(vis_r7_o[0]), 
	.C1(n16649), 
	.B2(vis_r3_o[0]), 
	.B1(n16877), 
	.A(n4479));
   OAI22_X2 U5007 (.ZN(n4479), 
	.B2(n16885), 
	.B1(n5039), 
	.A2(n4427), 
	.A1(n5040));
   NAND4_X2 U5012 (.ZN(n2028), 
	.A4(n4482), 
	.A3(n4481), 
	.A2(n4480), 
	.A1(n4169));
   AOI221_X1 U5013 (.ZN(n4482), 
	.C2(vis_r8_o[1]), 
	.C1(n16648), 
	.B2(vis_r10_o[1]), 
	.B1(n16897), 
	.A(n4484));
   OAI22_X1 U5014 (.ZN(n4484), 
	.B2(n4211), 
	.B1(n5255), 
	.A2(n16895), 
	.A1(n5287));
   AOI22_X1 U5017 (.ZN(n4481), 
	.B2(vis_r12_o[1]), 
	.B1(n16886), 
	.A2(vis_r9_o[1]), 
	.A1(n16891));
   NAND2_X1 U5020 (.ZN(n4480), 
	.A2(vis_r11_o[1]), 
	.A1(n16650));
   AND2_X1 U5022 (.ZN(n4169), 
	.A2(n4487), 
	.A1(n4486));
   AOI221_X1 U5023 (.ZN(n4487), 
	.C2(vis_r5_o[1]), 
	.C1(n16913), 
	.B2(vis_r4_o[1]), 
	.B1(n16916), 
	.A(n4488));
   OAI22_X1 U5024 (.ZN(n4488), 
	.B2(n16908), 
	.B1(n5172), 
	.A2(n16905), 
	.A1(n5453));
   AOI221_X1 U5027 (.ZN(n4486), 
	.C2(vis_r7_o[1]), 
	.C1(n16649), 
	.B2(vis_r3_o[1]), 
	.B1(n16877), 
	.A(n4491));
   OAI22_X1 U5028 (.ZN(n4491), 
	.B2(n16885), 
	.B1(n4986), 
	.A2(n4427), 
	.A1(n4987));
   NAND4_X2 U5031 (.ZN(n3287), 
	.A4(n4495), 
	.A3(n4494), 
	.A2(n4493), 
	.A1(n4492));
   AOI221_X1 U5032 (.ZN(n4495), 
	.C2(vis_r5_o[9]), 
	.C1(FE_OFN642_n16913), 
	.B2(vis_r4_o[9]), 
	.B1(n16916), 
	.A(n4496));
   OAI222_X1 U5033 (.ZN(n4496), 
	.C2(n16905), 
	.C1(n5476), 
	.B2(n16908), 
	.B1(n5195), 
	.A2(n16910), 
	.A1(n5140));
   AOI221_X1 U5036 (.ZN(n4494), 
	.C2(vis_r10_o[9]), 
	.C1(n16897), 
	.B2(vis_psp_o[7]), 
	.B1(n16902), 
	.A(n4497));
   OAI22_X1 U5037 (.ZN(n4497), 
	.B2(n16893), 
	.B1(n5576), 
	.A2(n16895), 
	.A1(n5575));
   AOI221_X1 U5040 (.ZN(n4493), 
	.C2(vis_r12_o[9]), 
	.C1(n16886), 
	.B2(vis_r9_o[9]), 
	.B1(n16891), 
	.A(n4498));
   OAI22_X1 U5041 (.ZN(n4498), 
	.B2(n16882), 
	.B1(n5418), 
	.A2(n16885), 
	.A1(n5141));
   AOI221_X1 U5044 (.ZN(n4492), 
	.C2(vis_r3_o[9]), 
	.C1(n16877), 
	.B2(vis_r0_o[9]), 
	.B1(n4224), 
	.A(n4500));
   OAI22_X1 U5045 (.ZN(n4500), 
	.B2(n16873), 
	.B1(n5331), 
	.A2(n16875), 
	.A1(n5143));
   NAND4_X2 U5050 (.ZN(n3145), 
	.A4(n4504), 
	.A3(n4503), 
	.A2(n4502), 
	.A1(n4501));
   AOI221_X1 U5051 (.ZN(n4504), 
	.C2(vis_r5_o[10]), 
	.C1(n16913), 
	.B2(vis_r4_o[10]), 
	.B1(n16916), 
	.A(n4505));
   OAI222_X1 U5052 (.ZN(n4505), 
	.C2(n16905), 
	.C1(n5474), 
	.B2(n16908), 
	.B1(n5193), 
	.A2(n16910), 
	.A1(n4771));
   AOI221_X1 U5055 (.ZN(n4503), 
	.C2(vis_r10_o[10]), 
	.C1(n16897), 
	.B2(vis_psp_o[8]), 
	.B1(n16902), 
	.A(n4506));
   OAI22_X1 U5056 (.ZN(n4506), 
	.B2(n16893), 
	.B1(n5147), 
	.A2(n16895), 
	.A1(n5302));
   AOI221_X1 U5059 (.ZN(n4502), 
	.C2(vis_r12_o[10]), 
	.C1(n16886), 
	.B2(vis_r9_o[10]), 
	.B1(n16891), 
	.A(n4507));
   OAI22_X1 U5060 (.ZN(n4507), 
	.B2(n16882), 
	.B1(n5416), 
	.A2(n16885), 
	.A1(n5144));
   AOI221_X1 U5063 (.ZN(n4501), 
	.C2(vis_r3_o[10]), 
	.C1(n16877), 
	.B2(vis_r0_o[10]), 
	.B1(n4224), 
	.A(n4509));
   OAI22_X1 U5064 (.ZN(n4509), 
	.B2(n16873), 
	.B1(n5329), 
	.A2(n16875), 
	.A1(n5146));
   NAND4_X2 U5067 (.ZN(n3177), 
	.A4(n4513), 
	.A3(n4512), 
	.A2(n4511), 
	.A1(n4510));
   AOI222_X1 U5068 (.ZN(n4513), 
	.C2(vis_msp_o[0]), 
	.C1(n16651), 
	.B2(n2620), 
	.B1(n16911), 
	.A2(vis_r14_o[2]), 
	.A1(n16652));
   AOI22_X1 U5072 (.ZN(n4512), 
	.B2(vis_r10_o[2]), 
	.B1(n16897), 
	.A2(vis_psp_o[0]), 
	.A1(n16902));
   AOI222_X1 U5075 (.ZN(n4511), 
	.C2(vis_r9_o[2]), 
	.C1(n16891), 
	.B2(vis_r8_o[2]), 
	.B1(n16648), 
	.A2(vis_r12_o[2]), 
	.A1(n16886));
   AOI21_X1 U5079 (.ZN(n4510), 
	.B2(vis_r11_o[2]), 
	.B1(n16650), 
	.A(n4171));
   NAND2_X2 U5080 (.ZN(n4171), 
	.A2(n4515), 
	.A1(n4514));
   AOI221_X2 U5081 (.ZN(n4515), 
	.C2(vis_r5_o[2]), 
	.C1(FE_OFN642_n16913), 
	.B2(vis_r4_o[2]), 
	.B1(FE_OFN643_n16916), 
	.A(n4516));
   OAI22_X1 U5082 (.ZN(n4516), 
	.B2(n16908), 
	.B1(n5194), 
	.A2(n16905), 
	.A1(n5475));
   AOI221_X2 U5085 (.ZN(n4514), 
	.C2(vis_r7_o[2]), 
	.C1(n16649), 
	.B2(vis_r3_o[2]), 
	.B1(n16877), 
	.A(n4519));
   OAI22_X1 U5086 (.ZN(n4519), 
	.B2(n16885), 
	.B1(n5056), 
	.A2(n4427), 
	.A1(n5499));
   NAND4_X2 U5092 (.ZN(n2246), 
	.A4(n4523), 
	.A3(n4522), 
	.A2(n4521), 
	.A1(n4520));
   AOI221_X1 U5093 (.ZN(n4523), 
	.C2(vis_r5_o[11]), 
	.C1(FE_OFN642_n16913), 
	.B2(vis_r4_o[11]), 
	.B1(FE_OFN643_n16916), 
	.A(n4524));
   OAI222_X1 U5094 (.ZN(n4524), 
	.C2(n16905), 
	.C1(n5556), 
	.B2(n16908), 
	.B1(n5564), 
	.A2(n16910), 
	.A1(n4831));
   AOI221_X1 U5097 (.ZN(n4522), 
	.C2(vis_r10_o[11]), 
	.C1(n16897), 
	.B2(vis_psp_o[9]), 
	.B1(n16902), 
	.A(n4525));
   OAI22_X1 U5098 (.ZN(n4525), 
	.B2(n16893), 
	.B1(n5568), 
	.A2(n16895), 
	.A1(n5567));
   AOI221_X1 U5101 (.ZN(n4521), 
	.C2(vis_r12_o[11]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[11]), 
	.B1(FE_OFN638_n16891), 
	.A(n4526));
   OAI22_X1 U5102 (.ZN(n4526), 
	.B2(n16882), 
	.B1(n5558), 
	.A2(n16885), 
	.A1(n5555));
   AOI221_X1 U5105 (.ZN(n4520), 
	.C2(vis_r3_o[11]), 
	.C1(n16877), 
	.B2(vis_r0_o[11]), 
	.B1(n4224), 
	.A(n4528));
   OAI22_X1 U5106 (.ZN(n4528), 
	.B2(n16873), 
	.B1(n5561), 
	.A2(n16875), 
	.A1(n5565));
   NAND4_X2 U5109 (.ZN(n2257), 
	.A4(n4532), 
	.A3(n4531), 
	.A2(n4530), 
	.A1(n4529));
   AOI222_X1 U5110 (.ZN(n4532), 
	.C2(vis_msp_o[1]), 
	.C1(n16651), 
	.B2(n2593), 
	.B1(n16911), 
	.A2(vis_r14_o[3]), 
	.A1(n16652));
   AOI22_X1 U5114 (.ZN(n4531), 
	.B2(vis_r10_o[3]), 
	.B1(n16897), 
	.A2(vis_psp_o[1]), 
	.A1(n16902));
   AOI222_X1 U5117 (.ZN(n4530), 
	.C2(vis_r9_o[3]), 
	.C1(n16891), 
	.B2(vis_r8_o[3]), 
	.B1(n16648), 
	.A2(vis_r12_o[3]), 
	.A1(n16886));
   AOI21_X1 U5121 (.ZN(n4529), 
	.B2(vis_r11_o[3]), 
	.B1(n16650), 
	.A(n4069));
   NAND2_X1 U5122 (.ZN(n4069), 
	.A2(n4534), 
	.A1(n4533));
   AOI221_X1 U5123 (.ZN(n4534), 
	.C2(vis_r5_o[3]), 
	.C1(FE_OFN642_n16913), 
	.B2(vis_r4_o[3]), 
	.B1(FE_OFN643_n16916), 
	.A(n4535));
   OAI22_X1 U5124 (.ZN(n4535), 
	.B2(n16908), 
	.B1(n5183), 
	.A2(n16905), 
	.A1(n5464));
   AOI221_X1 U5127 (.ZN(n4533), 
	.C2(vis_r7_o[3]), 
	.C1(n16649), 
	.B2(vis_r3_o[3]), 
	.B1(n16877), 
	.A(n4538));
   OAI22_X1 U5128 (.ZN(n4538), 
	.B2(n16885), 
	.B1(n5028), 
	.A2(n4427), 
	.A1(n5488));
   NAND4_X2 U5134 (.ZN(n2247), 
	.A4(n4542), 
	.A3(n4541), 
	.A2(n4540), 
	.A1(n4539));
   AOI221_X1 U5135 (.ZN(n4542), 
	.C2(vis_r5_o[12]), 
	.C1(FE_OFN642_n16913), 
	.B2(vis_r4_o[12]), 
	.B1(FE_OFN643_n16916), 
	.A(n4543));
   OAI222_X1 U5136 (.ZN(n4543), 
	.C2(n16905), 
	.C1(n5473), 
	.B2(n16908), 
	.B1(n5192), 
	.A2(n16910), 
	.A1(n4830));
   AOI221_X1 U5139 (.ZN(n4541), 
	.C2(vis_r10_o[12]), 
	.C1(FE_OFN639_n16897), 
	.B2(vis_psp_o[10]), 
	.B1(n16902), 
	.A(n4544));
   OAI22_X1 U5140 (.ZN(n4544), 
	.B2(n16893), 
	.B1(n5130), 
	.A2(n16895), 
	.A1(n5301));
   AOI221_X1 U5143 (.ZN(n4540), 
	.C2(vis_r12_o[12]), 
	.C1(FE_OFN636_n16886), 
	.B2(vis_r9_o[12]), 
	.B1(n16891), 
	.A(n4545));
   OAI22_X1 U5144 (.ZN(n4545), 
	.B2(n16882), 
	.B1(n5415), 
	.A2(n16885), 
	.A1(n5127));
   AOI221_X1 U5147 (.ZN(n4539), 
	.C2(vis_r3_o[12]), 
	.C1(n16877), 
	.B2(vis_r0_o[12]), 
	.B1(n4224), 
	.A(n4547));
   OAI22_X1 U5148 (.ZN(n4547), 
	.B2(n16873), 
	.B1(n5328), 
	.A2(n16875), 
	.A1(n5129));
   NAND4_X2 U5151 (.ZN(n2578), 
	.A4(n4551), 
	.A3(n4550), 
	.A2(n4549), 
	.A1(n4548));
   AOI222_X1 U5152 (.ZN(n4551), 
	.C2(vis_msp_o[2]), 
	.C1(n16651), 
	.B2(n2570), 
	.B1(n16911), 
	.A2(vis_r14_o[4]), 
	.A1(n16652));
   AOI22_X1 U5156 (.ZN(n4550), 
	.B2(vis_r10_o[4]), 
	.B1(n16897), 
	.A2(vis_psp_o[2]), 
	.A1(n16902));
   AOI222_X1 U5159 (.ZN(n4549), 
	.C2(vis_r9_o[4]), 
	.C1(n16891), 
	.B2(vis_r8_o[4]), 
	.B1(n16648), 
	.A2(vis_r12_o[4]), 
	.A1(n16886));
   AOI21_X1 U5163 (.ZN(n4548), 
	.B2(vis_r11_o[4]), 
	.B1(n16650), 
	.A(n4065));
   NAND2_X1 U5164 (.ZN(n4065), 
	.A2(n4553), 
	.A1(n4552));
   AOI221_X1 U5165 (.ZN(n4553), 
	.C2(vis_r5_o[4]), 
	.C1(FE_OFN642_n16913), 
	.B2(vis_r4_o[4]), 
	.B1(FE_OFN643_n16916), 
	.A(n4554));
   OAI22_X1 U5166 (.ZN(n4554), 
	.B2(n16908), 
	.B1(n5182), 
	.A2(n16905), 
	.A1(n5463));
   AOI221_X1 U5169 (.ZN(n4552), 
	.C2(vis_r7_o[4]), 
	.C1(n16649), 
	.B2(vis_r3_o[4]), 
	.B1(n16877), 
	.A(n4557));
   OAI22_X1 U5170 (.ZN(n4557), 
	.B2(n16885), 
	.B1(n5121), 
	.A2(n4427), 
	.A1(n5487));
   NAND4_X2 U5176 (.ZN(n2259), 
	.A4(n4561), 
	.A3(n4560), 
	.A2(n4559), 
	.A1(n4558));
   AOI221_X1 U5177 (.ZN(n4561), 
	.C2(vis_r5_o[13]), 
	.C1(n16913), 
	.B2(vis_r4_o[13]), 
	.B1(n16916), 
	.A(n4562));
   OAI222_X1 U5178 (.ZN(n4562), 
	.C2(n16905), 
	.C1(n5472), 
	.B2(n16908), 
	.B1(n5191), 
	.A2(n16910), 
	.A1(n4832));
   AOI221_X1 U5181 (.ZN(n4560), 
	.C2(vis_r10_o[13]), 
	.C1(n16897), 
	.B2(vis_psp_o[11]), 
	.B1(n16902), 
	.A(n4563));
   OAI22_X1 U5182 (.ZN(n4563), 
	.B2(n16893), 
	.B1(n5598), 
	.A2(n16895), 
	.A1(n5597));
   AOI221_X1 U5185 (.ZN(n4559), 
	.C2(vis_r12_o[13]), 
	.C1(n16886), 
	.B2(vis_r9_o[13]), 
	.B1(n16891), 
	.A(n4564));
   OAI22_X1 U5186 (.ZN(n4564), 
	.B2(n16882), 
	.B1(n5414), 
	.A2(n16885), 
	.A1(n5132));
   AOI221_X1 U5189 (.ZN(n4558), 
	.C2(vis_r3_o[13]), 
	.C1(n16877), 
	.B2(vis_r0_o[13]), 
	.B1(n4224), 
	.A(n4566));
   OAI22_X1 U5190 (.ZN(n4566), 
	.B2(n16873), 
	.B1(n5327), 
	.A2(n16875), 
	.A1(n5134));
   INV_X1 U5193 (.ZN(n4401), 
	.A(n4239));
   NOR3_X2 U5194 (.ZN(n4239), 
	.A3(n1612), 
	.A2(n5167), 
	.A1(FE_OFN495_n1670));
   AOI21_X1 U5195 (.ZN(n1670), 
	.B2(n4567), 
	.B1(n3362), 
	.A(n1612));
   OAI21_X1 U5196 (.ZN(n4567), 
	.B2(n632), 
	.B1(FE_OFN81_n16856), 
	.A(n556));
   NAND2_X2 U5197 (.ZN(n556), 
	.A2(FE_OFN82_n16856), 
	.A1(FE_OFN78_n16834));
   INV_X1 U5198 (.ZN(n632), 
	.A(n604));
   NAND2_X2 U5199 (.ZN(n604), 
	.A2(n16860), 
	.A1(FE_OFN79_n16834));
   NAND2_X1 U5200 (.ZN(n3362), 
	.A2(n16855), 
	.A1(n16837));
   NAND4_X2 U5201 (.ZN(n2556), 
	.A4(n4571), 
	.A3(n4570), 
	.A2(n4569), 
	.A1(n4568));
   AOI222_X1 U5202 (.ZN(n4571), 
	.C2(vis_msp_o[3]), 
	.C1(n16651), 
	.B2(n2539), 
	.B1(n16911), 
	.A2(vis_r14_o[5]), 
	.A1(n16652));
   AOI22_X1 U5206 (.ZN(n4570), 
	.B2(vis_r10_o[5]), 
	.B1(n16897), 
	.A2(vis_psp_o[3]), 
	.A1(n16902));
   AOI222_X1 U5209 (.ZN(n4569), 
	.C2(vis_r9_o[5]), 
	.C1(n16891), 
	.B2(vis_r8_o[5]), 
	.B1(n16648), 
	.A2(vis_r12_o[5]), 
	.A1(n16886));
   AOI21_X1 U5213 (.ZN(n4568), 
	.B2(vis_r11_o[5]), 
	.B1(n16650), 
	.A(n4058));
   NAND2_X1 U5214 (.ZN(n4058), 
	.A2(n4573), 
	.A1(n4572));
   AOI221_X1 U5215 (.ZN(n4573), 
	.C2(vis_r5_o[5]), 
	.C1(FE_OFN642_n16913), 
	.B2(vis_r4_o[5]), 
	.B1(FE_OFN643_n16916), 
	.A(n4574));
   OAI22_X1 U5216 (.ZN(n4574), 
	.B2(n16908), 
	.B1(n5181), 
	.A2(n16905), 
	.A1(n5462));
   AOI221_X1 U5219 (.ZN(n4572), 
	.C2(vis_r7_o[5]), 
	.C1(n16649), 
	.B2(vis_r3_o[5]), 
	.B1(n16877), 
	.A(n4577));
   OAI22_X1 U5220 (.ZN(n4577), 
	.B2(n16885), 
	.B1(n5091), 
	.A2(n4427), 
	.A1(n5486));
   NAND4_X2 U5226 (.ZN(n2196), 
	.A4(n4581), 
	.A3(n4580), 
	.A2(n4579), 
	.A1(n4578));
   AOI222_X1 U5227 (.ZN(n4581), 
	.C2(vis_msp_o[5]), 
	.C1(n16651), 
	.B2(n2221), 
	.B1(n16911), 
	.A2(vis_r14_o[7]), 
	.A1(n16652));
   AOI22_X1 U5234 (.ZN(n4580), 
	.B2(vis_r10_o[7]), 
	.B1(n16897), 
	.A2(vis_psp_o[5]), 
	.A1(n16902));
   AOI222_X1 U5237 (.ZN(n4579), 
	.C2(vis_r9_o[7]), 
	.C1(n16891), 
	.B2(vis_r8_o[7]), 
	.B1(n16648), 
	.A2(vis_r12_o[7]), 
	.A1(n16886));
   AOI21_X1 U5242 (.ZN(n4578), 
	.B2(vis_r11_o[7]), 
	.B1(n16650), 
	.A(n1795));
   NAND2_X1 U5243 (.ZN(n1795), 
	.A2(n4583), 
	.A1(n4582));
   AOI221_X1 U5244 (.ZN(n4583), 
	.C2(vis_r5_o[7]), 
	.C1(FE_OFN642_n16913), 
	.B2(vis_r4_o[7]), 
	.B1(FE_OFN643_n16916), 
	.A(n4584));
   OAI22_X1 U5245 (.ZN(n4584), 
	.B2(n16908), 
	.B1(n5171), 
	.A2(n16905), 
	.A1(n5452));
   AOI221_X1 U5248 (.ZN(n4582), 
	.C2(vis_r7_o[7]), 
	.C1(n16649), 
	.B2(vis_r3_o[7]), 
	.B1(n16877), 
	.A(n4587));
   OAI22_X1 U5249 (.ZN(n4587), 
	.B2(n16885), 
	.B1(n5021), 
	.A2(n4427), 
	.A1(n5022));
   NAND3_X1 U5258 (.ZN(n4589), 
	.A3(n3430), 
	.A2(FE_OFN632_n16859), 
	.A1(FE_OFN84_n16839));
   NAND2_X1 U5259 (.ZN(n4588), 
	.A2(n1094), 
	.A1(n1805));
   INV_X1 U5260 (.ZN(n1094), 
	.A(n1023));
   NAND2_X1 U5261 (.ZN(n1023), 
	.A2(n16867), 
	.A1(n16854));
   NAND2_X1 U5262 (.ZN(n1603), 
	.A2(n16838), 
	.A1(n16845));
   NAND4_X2 U5264 (.ZN(n3450), 
	.A4(n4594), 
	.A3(n4593), 
	.A2(n4592), 
	.A1(n4591));
   AOI221_X1 U5265 (.ZN(n4594), 
	.C2(vis_r5_o[23]), 
	.C1(n16913), 
	.B2(vis_r4_o[23]), 
	.B1(n16916), 
	.A(n4595));
   OAI222_X1 U5266 (.ZN(n4595), 
	.C2(n16905), 
	.C1(n5584), 
	.B2(n16908), 
	.B1(n5592), 
	.A2(n16910), 
	.A1(n4772));
   AOI221_X1 U5269 (.ZN(n4593), 
	.C2(vis_r10_o[23]), 
	.C1(n16897), 
	.B2(vis_psp_o[21]), 
	.B1(n16902), 
	.A(n4596));
   OAI22_X1 U5270 (.ZN(n4596), 
	.B2(n16893), 
	.B1(n4970), 
	.A2(n16895), 
	.A1(n5594));
   AOI221_X1 U5273 (.ZN(n4592), 
	.C2(vis_r12_o[23]), 
	.C1(n16886), 
	.B2(vis_r9_o[23]), 
	.B1(n16891), 
	.A(n4597));
   OAI22_X1 U5274 (.ZN(n4597), 
	.B2(n16882), 
	.B1(n5586), 
	.A2(n16885), 
	.A1(n4983));
   AOI221_X1 U5277 (.ZN(n4591), 
	.C2(vis_r3_o[23]), 
	.C1(n16877), 
	.B2(vis_r0_o[23]), 
	.B1(n4224), 
	.A(n4599));
   OAI22_X1 U5278 (.ZN(n4599), 
	.B2(n16873), 
	.B1(n5589), 
	.A2(n16875), 
	.A1(n4960));
   OAI22_X1 U5281 (.ZN(U189_Z_0), 
	.B2(n89), 
	.B1(n2462), 
	.A2(n4600), 
	.A1(n2461));
   INV_X1 U5282 (.ZN(n4600), 
	.A(n89));
   NAND4_X2 U5283 (.ZN(n89), 
	.A4(n4604), 
	.A3(n4603), 
	.A2(n4602), 
	.A1(n4601));
   AOI221_X1 U5284 (.ZN(n4604), 
	.C2(vis_r5_o[28]), 
	.C1(n16913), 
	.B2(vis_r4_o[28]), 
	.B1(n16916), 
	.A(n4605));
   OAI222_X1 U5285 (.ZN(n4605), 
	.C2(n16905), 
	.C1(n5451), 
	.B2(n16908), 
	.B1(n5170), 
	.A2(n16910), 
	.A1(n5626));
   AOI221_X1 U5288 (.ZN(n4603), 
	.C2(vis_r10_o[28]), 
	.C1(n16897), 
	.B2(vis_psp_o[26]), 
	.B1(n16902), 
	.A(n4606));
   OAI22_X1 U5289 (.ZN(n4606), 
	.B2(n16893), 
	.B1(n4994), 
	.A2(n16895), 
	.A1(n5285));
   AOI221_X1 U5292 (.ZN(n4602), 
	.C2(vis_r12_o[28]), 
	.C1(n16886), 
	.B2(vis_r9_o[28]), 
	.B1(n16891), 
	.A(n4607));
   OAI22_X1 U5293 (.ZN(n4607), 
	.B2(n16882), 
	.B1(n5393), 
	.A2(n16885), 
	.A1(n4997));
   AOI221_X1 U5296 (.ZN(n4601), 
	.C2(vis_r3_o[28]), 
	.C1(n16877), 
	.B2(vis_r0_o[28]), 
	.B1(n4224), 
	.A(n4609));
   OAI22_X1 U5297 (.ZN(n4609), 
	.B2(n16873), 
	.B1(n5306), 
	.A2(n16875), 
	.A1(n4996));
   INV_X1 U5301 (.ZN(n4610), 
	.A(n3534));
   NAND4_X2 U5302 (.ZN(n3534), 
	.A4(n4614), 
	.A3(n4613), 
	.A2(n4612), 
	.A1(n4611));
   AOI221_X1 U5303 (.ZN(n4614), 
	.C2(vis_r5_o[31]), 
	.C1(n16913), 
	.B2(vis_r4_o[31]), 
	.B1(n16916), 
	.A(n4615));
   OAI222_X1 U5304 (.ZN(n4615), 
	.C2(n16905), 
	.C1(n5450), 
	.B2(n16908), 
	.B1(n5169), 
	.A2(n16910), 
	.A1(n4774));
   AOI221_X1 U5307 (.ZN(n4613), 
	.C2(vis_r10_o[31]), 
	.C1(n16897), 
	.B2(vis_psp_o[29]), 
	.B1(n16902), 
	.A(n4616));
   OAI22_X1 U5308 (.ZN(n4616), 
	.B2(n16893), 
	.B1(n4969), 
	.A2(n16895), 
	.A1(n5284));
   AOI221_X1 U5311 (.ZN(n4612), 
	.C2(vis_r12_o[31]), 
	.C1(n16886), 
	.B2(vis_r9_o[31]), 
	.B1(n16891), 
	.A(n4617));
   OAI22_X1 U5312 (.ZN(n4617), 
	.B2(n16882), 
	.B1(n5392), 
	.A2(n16885), 
	.A1(n4981));
   AOI221_X1 U5315 (.ZN(n4611), 
	.C2(vis_r3_o[31]), 
	.C1(n16877), 
	.B2(vis_r0_o[31]), 
	.B1(n4224), 
	.A(n4619));
   OAI22_X1 U5316 (.ZN(n4619), 
	.B2(n16873), 
	.B1(n5305), 
	.A2(n16875), 
	.A1(n4962));
   OAI22_X1 U5319 (.ZN(U180_Z_0), 
	.B2(n2083), 
	.B1(n2462), 
	.A2(n4620), 
	.A1(n2461));
   INV_X1 U5320 (.ZN(n4620), 
	.A(n2083));
   NAND4_X2 U5321 (.ZN(n2083), 
	.A4(n4624), 
	.A3(n4623), 
	.A2(n4622), 
	.A1(n4621));
   AOI221_X1 U5322 (.ZN(n4624), 
	.C2(vis_r5_o[30]), 
	.C1(n16913), 
	.B2(vis_r4_o[30]), 
	.B1(n16916), 
	.A(n4625));
   OAI222_X1 U5323 (.ZN(n4625), 
	.C2(n16905), 
	.C1(n5455), 
	.B2(n16908), 
	.B1(n5174), 
	.A2(n16910), 
	.A1(n4955));
   AOI221_X1 U5326 (.ZN(n4623), 
	.C2(vis_r10_o[30]), 
	.C1(n16897), 
	.B2(vis_psp_o[28]), 
	.B1(n16902), 
	.A(n4626));
   OAI22_X1 U5327 (.ZN(n4626), 
	.B2(n16893), 
	.B1(n5642), 
	.A2(n16895), 
	.A1(n5641));
   AOI221_X1 U5330 (.ZN(n4622), 
	.C2(vis_r12_o[30]), 
	.C1(n16886), 
	.B2(vis_r9_o[30]), 
	.B1(n16891), 
	.A(n4627));
   OAI22_X1 U5331 (.ZN(n4627), 
	.B2(n16882), 
	.B1(n5397), 
	.A2(n16885), 
	.A1(n5080));
   AOI221_X1 U5334 (.ZN(n4621), 
	.C2(vis_r3_o[30]), 
	.C1(n16877), 
	.B2(vis_r0_o[30]), 
	.B1(n4224), 
	.A(n4629));
   OAI22_X1 U5335 (.ZN(n4629), 
	.B2(n16873), 
	.B1(n5310), 
	.A2(n16875), 
	.A1(n5082));
   OAI22_X1 U5338 (.ZN(U175_Z_0), 
	.B2(n2427), 
	.B1(n2462), 
	.A2(n4630), 
	.A1(n2461));
   INV_X1 U5339 (.ZN(n4630), 
	.A(n2427));
   NAND4_X1 U5340 (.ZN(n2427), 
	.A4(n4634), 
	.A3(n4633), 
	.A2(n4632), 
	.A1(n4631));
   AOI221_X1 U5341 (.ZN(n4634), 
	.C2(vis_r5_o[27]), 
	.C1(n16913), 
	.B2(vis_r4_o[27]), 
	.B1(n16916), 
	.A(n4635));
   OAI222_X1 U5342 (.ZN(n4635), 
	.C2(n16905), 
	.C1(n5457), 
	.B2(n16908), 
	.B1(n5176), 
	.A2(n16910), 
	.A1(n4761));
   AOI221_X1 U5345 (.ZN(n4633), 
	.C2(vis_r10_o[27]), 
	.C1(n16897), 
	.B2(vis_psp_o[25]), 
	.B1(n16902), 
	.A(n4636));
   OAI22_X1 U5346 (.ZN(n4636), 
	.B2(n16893), 
	.B1(n5629), 
	.A2(n16895), 
	.A1(n5628));
   AOI221_X1 U5349 (.ZN(n4632), 
	.C2(vis_r12_o[27]), 
	.C1(n16886), 
	.B2(vis_r9_o[27]), 
	.B1(n16891), 
	.A(n4637));
   OAI22_X1 U5350 (.ZN(n4637), 
	.B2(n16882), 
	.B1(n5399), 
	.A2(n16885), 
	.A1(n5111));
   AOI221_X1 U5353 (.ZN(n4631), 
	.C2(vis_r3_o[27]), 
	.C1(n16877), 
	.B2(vis_r0_o[27]), 
	.B1(n4224), 
	.A(n4639));
   OAI22_X1 U5354 (.ZN(n4639), 
	.B2(n16873), 
	.B1(n5312), 
	.A2(n16875), 
	.A1(n5113));
   OAI22_X1 U5357 (.ZN(U163_Z_0), 
	.B2(n2496), 
	.B1(n2462), 
	.A2(n4640), 
	.A1(n2461));
   INV_X1 U5358 (.ZN(n4640), 
	.A(n2496));
   NAND4_X1 U5359 (.ZN(n2496), 
	.A4(n4644), 
	.A3(n4643), 
	.A2(n4642), 
	.A1(n4641));
   AOI221_X1 U5360 (.ZN(n4644), 
	.C2(vis_r5_o[24]), 
	.C1(n16913), 
	.B2(vis_r4_o[24]), 
	.B1(n16916), 
	.A(n4645));
   OAI222_X1 U5361 (.ZN(n4645), 
	.C2(n16905), 
	.C1(n5460), 
	.B2(n16908), 
	.B1(n5179), 
	.A2(n16910), 
	.A1(n4971));
   AOI221_X1 U5364 (.ZN(n4643), 
	.C2(vis_r10_o[24]), 
	.C1(n16897), 
	.B2(vis_psp_o[22]), 
	.B1(n16902), 
	.A(n4646));
   OAI22_X1 U5365 (.ZN(n4646), 
	.B2(n16893), 
	.B1(n5646), 
	.A2(n16895), 
	.A1(n5645));
   AOI221_X1 U5368 (.ZN(n4642), 
	.C2(vis_r12_o[24]), 
	.C1(n16886), 
	.B2(vis_r9_o[24]), 
	.B1(n16891), 
	.A(n4647));
   OAI22_X1 U5369 (.ZN(n4647), 
	.B2(n16882), 
	.B1(n5402), 
	.A2(n16885), 
	.A1(n4982));
   AOI221_X1 U5372 (.ZN(n4641), 
	.C2(vis_r3_o[24]), 
	.C1(n16877), 
	.B2(vis_r0_o[24]), 
	.B1(n4224), 
	.A(n4649));
   OAI22_X1 U5373 (.ZN(n4649), 
	.B2(n16873), 
	.B1(n5315), 
	.A2(n16875), 
	.A1(n4972));
   OAI22_X1 U5376 (.ZN(U158_Z_0), 
	.B2(n4650), 
	.B1(n2461), 
	.A2(n1755), 
	.A1(n2462));
   INV_X1 U5377 (.ZN(n4650), 
	.A(n1755));
   INV_X1 U5378 (.ZN(n2461), 
	.A(n2492));
   OAI21_X1 U5379 (.ZN(n2492), 
	.B2(FE_OFN559_n3180), 
	.B1(n16991), 
	.A(n4651));
   NAND4_X2 U5381 (.ZN(n1755), 
	.A4(n4655), 
	.A3(n4654), 
	.A2(n4653), 
	.A1(n4652));
   AOI221_X1 U5382 (.ZN(n4655), 
	.C2(vis_r5_o[29]), 
	.C1(n16913), 
	.B2(vis_r4_o[29]), 
	.B1(n16916), 
	.A(n4656));
   OAI222_X1 U5383 (.ZN(n4656), 
	.C2(n16905), 
	.C1(n5456), 
	.B2(n16908), 
	.B1(n5175), 
	.A2(n16910), 
	.A1(n4773));
   NAND2_X1 U5386 (.ZN(n4211), 
	.A2(n4661), 
	.A1(n4660));
   AOI221_X1 U5391 (.ZN(n4654), 
	.C2(vis_r10_o[29]), 
	.C1(n16897), 
	.B2(vis_psp_o[27]), 
	.B1(n16902), 
	.A(n4664));
   OAI22_X1 U5392 (.ZN(n4664), 
	.B2(n16893), 
	.B1(n5078), 
	.A2(n16895), 
	.A1(n5289));
   NOR2_X1 U5397 (.ZN(n4658), 
	.A2(n5545), 
	.A1(n3489));
   AOI221_X1 U5401 (.ZN(n4653), 
	.C2(vis_r12_o[29]), 
	.C1(n16886), 
	.B2(vis_r9_o[29]), 
	.B1(n16891), 
	.A(n4666));
   OAI22_X1 U5402 (.ZN(n4666), 
	.B2(n16882), 
	.B1(n5398), 
	.A2(n16885), 
	.A1(n5075));
   NOR2_X1 U5407 (.ZN(n4660), 
	.A2(n5259), 
	.A1(n5544));
   NOR2_X1 U5410 (.ZN(n4662), 
	.A2(n5004), 
	.A1(n1353));
   AOI221_X1 U5411 (.ZN(n4652), 
	.C2(vis_r3_o[29]), 
	.C1(n16877), 
	.B2(vis_r0_o[29]), 
	.B1(n4224), 
	.A(n4668));
   OAI22_X1 U5412 (.ZN(n4668), 
	.B2(n16873), 
	.B1(n5311), 
	.A2(n16875), 
	.A1(n5077));
   NOR2_X1 U5414 (.ZN(n4665), 
	.A2(n5544), 
	.A1(n3493));
   NOR2_X2 U5416 (.ZN(n4659), 
	.A2(n5259), 
	.A1(n3496));
   NOR2_X1 U5419 (.ZN(n4661), 
	.A2(n5545), 
	.A1(n5004));
   INV_X4 U5421 (.ZN(n4224), 
	.A(n4427));
   NOR2_X1 U5423 (.ZN(n4657), 
	.A2(n3496), 
	.A1(n3493));
   NOR2_X2 U5426 (.ZN(n4663), 
	.A2(n3489), 
	.A1(n1353));
   INV_X1 U5429 (.ZN(n2462), 
	.A(n2493));
   OAI21_X1 U5430 (.ZN(n2493), 
	.B2(n16990), 
	.B1(n4669), 
	.A(n4651));
   AOI21_X1 U5431 (.ZN(n4651), 
	.B2(n4669), 
	.B1(n16990), 
	.A(n4670));
   NOR3_X1 U5432 (.ZN(n4670), 
	.A3(n16990), 
	.A2(n16988), 
	.A1(n4669));
   OAI21_X1 U5434 (.ZN(n3180), 
	.B2(n4672), 
	.B1(n4671), 
	.A(FE_OFN10_n1697));
   OAI222_X1 U5435 (.ZN(n4672), 
	.C2(n758), 
	.C1(n16833), 
	.B2(n4673), 
	.B1(n16851), 
	.A2(n673), 
	.A1(n1784));
   INV_X1 U5436 (.ZN(n758), 
	.A(n515));
   NOR2_X1 U5437 (.ZN(n515), 
	.A2(n16825), 
	.A1(FE_OFN17_n16805));
   NOR4_X1 U5438 (.ZN(n4673), 
	.A4(n4674), 
	.A3(n529), 
	.A2(n2042), 
	.A1(n3506));
   NOR3_X1 U5439 (.ZN(n4674), 
	.A3(FE_OFN85_n16839), 
	.A2(n16828), 
	.A1(n617));
   INV_X1 U5441 (.ZN(n2042), 
	.A(n666));
   NAND2_X1 U5442 (.ZN(n666), 
	.A2(n16831), 
	.A1(n16855));
   INV_X1 U5443 (.ZN(n3506), 
	.A(n1103));
   NAND2_X1 U5444 (.ZN(n1103), 
	.A2(n16831), 
	.A1(n16826));
   OAI221_X1 U5446 (.ZN(n4671), 
	.C2(n16867), 
	.C1(n16824), 
	.B2(n1278), 
	.B1(n617), 
	.A(n4675));
   NAND3_X1 U5447 (.ZN(n4675), 
	.A3(n1042), 
	.A2(n991), 
	.A1(n1805));
   INV_X1 U5448 (.ZN(n1042), 
	.A(n641));
   NAND2_X1 U5449 (.ZN(n641), 
	.A2(FE_OFN90_n16849), 
	.A1(FE_OFN81_n16856));
   INV_X4 U5452 (.ZN(n1805), 
	.A(n1579));
   NAND2_X1 U5453 (.ZN(n1579), 
	.A2(n16860), 
	.A1(n16837));
   NAND2_X2 U5454 (.ZN(n1278), 
	.A2(n16831), 
	.A1(n565));
   OAI211_X1 U5456 (.ZN(n4676), 
	.C2(n890), 
	.C1(n16859), 
	.B(n4678), 
	.A(n4677));
   AOI21_X1 U5457 (.ZN(n4678), 
	.B2(n1564), 
	.B1(n667), 
	.A(n4679));
   OAI33_X1 U5458 (.ZN(n4679), 
	.B3(n4680), 
	.B2(n16824), 
	.B1(FE_OFN72_n16867), 
	.A3(FE_OFN70_n16867), 
	.A2(FE_OFN633_n16868), 
	.A1(n1518));
   AOI21_X1 U5459 (.ZN(n4680), 
	.B2(n16842), 
	.B1(n16862), 
	.A(n501));
   INV_X4 U5460 (.ZN(n501), 
	.A(n617));
   NAND2_X1 U5462 (.ZN(n1518), 
	.A2(n16860), 
	.A1(n2646));
   INV_X1 U5463 (.ZN(n2646), 
	.A(n1233));
   NAND2_X1 U5464 (.ZN(n1233), 
	.A2(FE_OFN85_n16839), 
	.A1(n16842));
   INV_X4 U5465 (.ZN(n1564), 
	.A(n1580));
   NAND2_X2 U5466 (.ZN(n1580), 
	.A2(n16843), 
	.A1(n16851));
   INV_X1 U5467 (.ZN(n667), 
	.A(n1706));
   NAND2_X1 U5468 (.ZN(n1706), 
	.A2(FE_OFN85_n16839), 
	.A1(n16828));
   INV_X1 U5469 (.ZN(n4677), 
	.A(n1705));
   OAI222_X1 U5470 (.ZN(n1705), 
	.C2(n1517), 
	.C1(FE_OFN633_n16868), 
	.B2(n568), 
	.B1(n745), 
	.A2(n849), 
	.A1(n1104));
   NAND2_X2 U5471 (.ZN(n568), 
	.A2(n16690), 
	.A1(n16837));
   NAND2_X2 U5472 (.ZN(n849), 
	.A2(FE_OFN85_n16839), 
	.A1(FE_OFN70_n16867));
   NAND2_X1 U5473 (.ZN(n890), 
	.A2(n17096), 
	.A1(n565));
   OR2_X1 U5475 (.ZN(n4669), 
	.A2(n2716), 
	.A1(n2732));
   NOR2_X1 U5476 (.ZN(n2716), 
	.A2(n5254), 
	.A1(n2543));
   NAND4_X1 U5477 (.ZN(n2543), 
	.A4(FE_OFN10_n1697), 
	.A3(n16826), 
	.A2(FE_OFN628_n16833), 
	.A1(n3430));
   INV_X4 U5478 (.ZN(n3430), 
	.A(n1104));
   NAND2_X1 U5481 (.ZN(n2719), 
	.A2(n1723), 
	.A1(n3164));
   INV_X1 U5482 (.ZN(n3164), 
	.A(n3186));
   NAND3_X1 U5483 (.ZN(n3186), 
	.A3(n483), 
	.A2(FE_OFN10_n1697), 
	.A1(n1095));
   INV_X4 U5485 (.ZN(n1095), 
	.A(n1784));
   NAND2_X2 U5486 (.ZN(n1784), 
	.A2(n16843), 
	.A1(n16854));
   OAI22_X1 U5487 (.ZN(U144_Z_0), 
	.B2(n4683), 
	.B1(n4682), 
	.A2(n4681), 
	.A1(n4959));
   AOI21_X1 U5488 (.ZN(n4682), 
	.B2(n16798), 
	.B1(n4684), 
	.A(n4685));
   OAI21_X1 U5489 (.ZN(n4684), 
	.B2(n4686), 
	.B1(n16816), 
	.A(n782));
   OAI22_X1 U5490 (.ZN(U134_Z_0), 
	.B2(n4683), 
	.B1(n4687), 
	.A2(n4681), 
	.A1(n4978));
   AOI211_X1 U5491 (.ZN(n4687), 
	.C2(n451), 
	.C1(n4688), 
	.B(n4685), 
	.A(n4689));
   OAI22_X1 U5492 (.ZN(n4689), 
	.B2(n4691), 
	.B1(n17099), 
	.A2(n4690), 
	.A1(n16794));
   OAI22_X1 U5493 (.ZN(U122_Z_0), 
	.B2(n1715), 
	.B1(n4692), 
	.A2(n1713), 
	.A1(FE_PHN3764_n5004));
   AOI211_X1 U5494 (.ZN(n4692), 
	.C2(n486), 
	.C1(n597), 
	.B(n4694), 
	.A(n4693));
   OAI22_X1 U5495 (.ZN(n4694), 
	.B2(n1719), 
	.B1(n4967), 
	.A2(n1307), 
	.A1(n4695));
   NAND2_X1 U5496 (.ZN(n1719), 
	.A2(n16816), 
	.A1(n473));
   AOI221_X1 U5497 (.ZN(n4695), 
	.C2(n664), 
	.C1(n4697), 
	.B2(n1286), 
	.B1(n4696), 
	.A(n4698));
   OAI22_X1 U5498 (.ZN(n4698), 
	.B2(n437), 
	.B1(n4699), 
	.A2(n486), 
	.A1(n5003));
   NAND2_X1 U5499 (.ZN(n664), 
	.A2(n4697), 
	.A1(n5258));
   INV_X1 U5500 (.ZN(n4697), 
	.A(n1294));
   OAI221_X1 U5501 (.ZN(n4693), 
	.C2(n819), 
	.C1(n16801), 
	.B2(n1721), 
	.B1(n16794), 
	.A(n1720));
   NOR3_X1 U5502 (.ZN(n1720), 
	.A3(n896), 
	.A2(n1478), 
	.A1(n483));
   INV_X1 U5503 (.ZN(n896), 
	.A(n1170));
   NOR2_X1 U5504 (.ZN(n1170), 
	.A2(n493), 
	.A1(n784));
   NOR2_X1 U5505 (.ZN(n493), 
	.A2(n16845), 
	.A1(n640));
   INV_X1 U5506 (.ZN(n784), 
	.A(n4318));
   NAND2_X1 U5507 (.ZN(n4318), 
	.A2(n16843), 
	.A1(n608));
   INV_X1 U5508 (.ZN(n608), 
	.A(n745));
   OAI21_X1 U5510 (.ZN(n1721), 
	.B2(n16817), 
	.B1(n822), 
	.A(n1728));
   NAND2_X1 U5511 (.ZN(n1728), 
	.A2(n1198), 
	.A1(n1594));
   INV_X1 U5514 (.ZN(n1713), 
	.A(n1715));
   NAND2_X1 U5515 (.ZN(n1715), 
	.A2(n4700), 
	.A1(n17124));
   NAND4_X1 U5516 (.ZN(n4700), 
	.A4(n4704), 
	.A3(n4703), 
	.A2(n4702), 
	.A1(n4701));
   NOR4_X1 U5517 (.ZN(n4704), 
	.A4(n4705), 
	.A3(n1302), 
	.A2(n495), 
	.A1(n741));
   NOR4_X1 U5518 (.ZN(n4705), 
	.A4(n1307), 
	.A3(n918), 
	.A2(n16821), 
	.A1(n16828));
   INV_X4 U5519 (.ZN(n1307), 
	.A(n614));
   NOR2_X1 U5520 (.ZN(n614), 
	.A2(n16826), 
	.A1(n4590));
   NAND2_X1 U5521 (.ZN(n4590), 
	.A2(n16851), 
	.A1(n16870));
   NOR2_X1 U5523 (.ZN(n1302), 
	.A2(n1467), 
	.A1(n3528));
   INV_X1 U5524 (.ZN(n1467), 
	.A(n911));
   NAND3_X1 U5525 (.ZN(n911), 
	.A3(n5230), 
	.A2(vis_pc_o[2]), 
	.A1(n3313));
   NOR4_X1 U5528 (.ZN(n495), 
	.A4(n16854), 
	.A3(n16826), 
	.A2(n640), 
	.A1(n610));
   AOI222_X1 U5530 (.ZN(n4708), 
	.C2(n1723), 
	.C1(n437), 
	.B2(FE_OFN15_n16671), 
	.B1(n776), 
	.A2(FE_OFN549_n2774), 
	.A1(n486));
   AOI22_X1 U5535 (.ZN(n4707), 
	.B2(n2865), 
	.B1(n768), 
	.A2(n2731), 
	.A1(n455));
   AOI22_X1 U5538 (.ZN(n4706), 
	.B2(n2827), 
	.B1(n1286), 
	.A2(n2819), 
	.A1(n1294));
   NAND2_X1 U5541 (.ZN(n1294), 
	.A2(n1976), 
	.A1(n5257));
   INV_X1 U5542 (.ZN(n1976), 
	.A(n1286));
   NAND2_X1 U5543 (.ZN(n1286), 
	.A2(n4696), 
	.A1(FE_PHN1586_n5256));
   INV_X1 U5544 (.ZN(n4696), 
	.A(n768));
   NAND2_X1 U5545 (.ZN(n768), 
	.A2(n16810), 
	.A1(n4699));
   INV_X1 U5546 (.ZN(n4699), 
	.A(n776));
   NAND2_X1 U5547 (.ZN(n776), 
	.A2(n1974), 
	.A1(n5254));
   INV_X1 U5548 (.ZN(n1974), 
	.A(n437));
   NAND2_X1 U5549 (.ZN(n437), 
	.A2(n1975), 
	.A1(n5253));
   INV_X1 U5550 (.ZN(n1975), 
	.A(n455));
   NAND2_X1 U5551 (.ZN(n455), 
	.A2(n5162), 
	.A1(n5003));
   INV_X1 U5552 (.ZN(n741), 
	.A(n619));
   NAND2_X1 U5553 (.ZN(n619), 
	.A2(FE_OFN90_n16849), 
	.A1(n1478));
   INV_X1 U5554 (.ZN(n1478), 
	.A(n694));
   NAND2_X1 U5555 (.ZN(n694), 
	.A2(n16860), 
	.A1(n527));
   AOI222_X1 U5556 (.ZN(n4703), 
	.C2(n589), 
	.C1(n4712), 
	.B2(n1265), 
	.B1(n4711), 
	.A2(n4710), 
	.A1(n4709));
   NOR2_X1 U5557 (.ZN(n4712), 
	.A2(FE_OFN87_n16848), 
	.A1(n16837));
   INV_X1 U5558 (.ZN(n1265), 
	.A(n1908));
   NAND3_X1 U5559 (.ZN(n1908), 
	.A3(n732), 
	.A2(n16820), 
	.A1(n16811));
   INV_X1 U5560 (.ZN(n732), 
	.A(n819));
   AOI21_X1 U5562 (.ZN(n4711), 
	.B2(n1562), 
	.B1(n16803), 
	.A(FE_OFN21_n503));
   NAND2_X1 U5563 (.ZN(n1562), 
	.A2(n16733), 
	.A1(n16816));
   NAND2_X1 U5564 (.ZN(n4710), 
	.A2(n1303), 
	.A1(n1517));
   NAND2_X1 U5565 (.ZN(n1303), 
	.A2(n16867), 
	.A1(n526));
   NAND2_X1 U5566 (.ZN(n1517), 
	.A2(n16838), 
	.A1(FE_OFN70_n16867));
   INV_X1 U5567 (.ZN(n4709), 
	.A(n514));
   NAND2_X2 U5568 (.ZN(n514), 
	.A2(n16870), 
	.A1(n592));
   AOI222_X1 U5569 (.ZN(n4702), 
	.C2(n16821), 
	.C1(n4715), 
	.B2(n4714), 
	.B1(n16814), 
	.A2(n4713), 
	.A1(n333));
   INV_X1 U5570 (.ZN(n4715), 
	.A(n3528));
   NAND2_X1 U5571 (.ZN(n3528), 
	.A2(n527), 
	.A1(n195));
   OAI33_X1 U5576 (.ZN(n4714), 
	.B3(n1928), 
	.B2(FE_OFN426_n659), 
	.B1(n4717), 
	.A3(n583), 
	.A2(n1920), 
	.A1(n4716));
   NAND2_X1 U5577 (.ZN(n1928), 
	.A2(n16686), 
	.A1(n16725));
   NAND3_X1 U5579 (.ZN(n4717), 
	.A3(n721), 
	.A2(n505), 
	.A1(n440));
   INV_X1 U5580 (.ZN(n505), 
	.A(n469));
   INV_X1 U5581 (.ZN(n440), 
	.A(n892));
   NAND3_X1 U5582 (.ZN(n892), 
	.A3(n821), 
	.A2(n16820), 
	.A1(n708));
   INV_X1 U5583 (.ZN(n821), 
	.A(n1552));
   NAND2_X1 U5584 (.ZN(n583), 
	.A2(n17099), 
	.A1(n504));
   NOR2_X1 U5585 (.ZN(n504), 
	.A2(n5244), 
	.A1(n669));
   NAND2_X1 U5586 (.ZN(n669), 
	.A2(n16674), 
	.A1(n16800));
   NAND2_X1 U5588 (.ZN(n4716), 
	.A2(n731), 
	.A1(n476));
   INV_X1 U5589 (.ZN(n476), 
	.A(n443));
   NAND2_X1 U5592 (.ZN(n579), 
	.A2(n16820), 
	.A1(n16804));
   NAND2_X1 U5594 (.ZN(n1198), 
	.A2(n16683), 
	.A1(n16871));
   INV_X1 U5595 (.ZN(n4713), 
	.A(n479));
   NAND2_X1 U5596 (.ZN(n479), 
	.A2(n16820), 
	.A1(n1492));
   INV_X1 U5597 (.ZN(n1492), 
	.A(n725));
   NAND2_X1 U5598 (.ZN(n725), 
	.A2(n16802), 
	.A1(n475));
   INV_X1 U5599 (.ZN(n333), 
	.A(n932));
   NAND2_X1 U5600 (.ZN(n932), 
	.A2(n791), 
	.A1(n16812));
   INV_X1 U5601 (.ZN(n791), 
	.A(n1261));
   AOI221_X1 U5602 (.ZN(n4701), 
	.C2(n526), 
	.C1(n506), 
	.B2(n16734), 
	.B1(n1263), 
	.A(n1883));
   OAI21_X1 U5603 (.ZN(n1883), 
	.B2(n4718), 
	.B1(n650), 
	.A(n1957));
   NAND2_X1 U5604 (.ZN(n1957), 
	.A2(n16843), 
	.A1(n17096));
   NAND2_X1 U5605 (.ZN(n4718), 
	.A2(n16831), 
	.A1(n997));
   INV_X4 U5606 (.ZN(n997), 
	.A(n653));
   NAND2_X1 U5611 (.ZN(n1882), 
	.A2(n16843), 
	.A1(FE_OFN626_n16820));
   INV_X2 U5616 (.ZN(n506), 
	.A(n1465));
   NAND2_X1 U5617 (.ZN(n1465), 
	.A2(n16831), 
	.A1(n589));
   INV_X4 U5618 (.ZN(n589), 
	.A(n696));
   NOR3_X1 U5619 (.ZN(n1263), 
	.A3(n594), 
	.A2(n16839), 
	.A1(n851));
   NAND4_X1 U5620 (.ZN(n594), 
	.A4(FE_OFN631_n16851), 
	.A3(n16803), 
	.A2(n1468), 
	.A1(n483));
   NAND2_X1 U5622 (.ZN(n945), 
	.A2(n16826), 
	.A1(n16870));
   OAI22_X1 U5625 (.ZN(U121_Z_0), 
	.B2(n4683), 
	.B1(n4719), 
	.A2(n4681), 
	.A1(n5036));
   AOI211_X1 U5626 (.ZN(n4719), 
	.C2(n461), 
	.C1(n4688), 
	.B(n4721), 
	.A(n4720));
   OAI221_X1 U5627 (.ZN(n4720), 
	.C2(n4690), 
	.C1(n5243), 
	.B2(n4691), 
	.B1(n16796), 
	.A(n4722));
   NAND4_X1 U5628 (.ZN(n4722), 
	.A4(n16683), 
	.A3(n592), 
	.A2(n1468), 
	.A1(n16814));
   OAI22_X1 U5629 (.ZN(U105_Z_0), 
	.B2(n4683), 
	.B1(n4723), 
	.A2(n4681), 
	.A1(n5252));
   AOI211_X1 U5630 (.ZN(n4723), 
	.C2(n454), 
	.C1(n4688), 
	.B(n4685), 
	.A(n4724));
   NAND4_X1 U5631 (.ZN(n4685), 
	.A4(n4727), 
	.A3(n4726), 
	.A2(n755), 
	.A1(n4725));
   AOI21_X1 U5632 (.ZN(n4727), 
	.B2(n16683), 
	.B1(n1468), 
	.A(n4721));
   OAI221_X1 U5633 (.ZN(n4721), 
	.C2(n1920), 
	.C1(n4729), 
	.B2(n4686), 
	.B1(n4728), 
	.A(n4730));
   OR4_X1 U5634 (.ZN(n4730), 
	.A4(n16794), 
	.A3(n782), 
	.A2(n461), 
	.A1(n451));
   AOI21_X1 U5637 (.ZN(n4728), 
	.B2(n16686), 
	.B1(n731), 
	.A(n16813));
   NOR2_X1 U5638 (.ZN(n1468), 
	.A2(n16811), 
	.A1(n16725));
   OAI21_X1 U5639 (.ZN(n4726), 
	.B2(n16734), 
	.B1(FE_OFN631_n16851), 
	.A(FE_OFN17_n16805));
   OAI21_X1 U5640 (.ZN(n4725), 
	.B2(n16807), 
	.B1(n16796), 
	.A(n630));
   OAI22_X1 U5641 (.ZN(n4724), 
	.B2(n4691), 
	.B1(n16816), 
	.A2(n4690), 
	.A1(n5244));
   OAI221_X1 U5642 (.ZN(n4691), 
	.C2(n16802), 
	.C1(n16811), 
	.B2(n16659), 
	.B1(n1547), 
	.A(n592));
   NOR2_X1 U5643 (.ZN(n1547), 
	.A2(n16807), 
	.A1(n16802));
   OAI21_X1 U5644 (.ZN(n4690), 
	.B2(n4732), 
	.B1(n4731), 
	.A(n592));
   OAI33_X1 U5645 (.ZN(n4732), 
	.B3(n16659), 
	.B2(n16795), 
	.B1(n16683), 
	.A3(n16725), 
	.A2(n16802), 
	.A1(n16683));
   NAND2_X1 U5646 (.ZN(n4731), 
	.A2(n1552), 
	.A1(n4733));
   NAND2_X1 U5647 (.ZN(n1552), 
	.A2(n16683), 
	.A1(n16802));
   NAND3_X1 U5648 (.ZN(n4733), 
	.A3(n630), 
	.A2(n16683), 
	.A1(n16657));
   INV_X1 U5649 (.ZN(n630), 
	.A(n1920));
   NAND2_X1 U5650 (.ZN(n1920), 
	.A2(n16725), 
	.A1(n16659));
   OAI21_X1 U5653 (.ZN(n4688), 
	.B2(n16734), 
	.B1(n782), 
	.A(n4686));
   NAND4_X1 U5654 (.ZN(n4686), 
	.A4(n16795), 
	.A3(n2672), 
	.A2(n16811), 
	.A1(n16807));
   INV_X1 U5655 (.ZN(n2672), 
	.A(n4729));
   NAND2_X1 U5656 (.ZN(n4729), 
	.A2(n16802), 
	.A1(n592));
   NAND2_X1 U5661 (.ZN(n782), 
	.A2(FE_OFN17_n16805), 
	.A1(FE_OFN90_n16849));
   INV_X1 U5663 (.ZN(n4681), 
	.A(n4683));
   OAI21_X1 U5664 (.ZN(n4683), 
	.B2(n4735), 
	.B1(n4734), 
	.A(n17124));
   OAI221_X1 U5665 (.ZN(n4735), 
	.C2(n696), 
	.C1(n1519), 
	.B2(n692), 
	.B1(FE_OFN72_n16867), 
	.A(n488));
   INV_X1 U5666 (.ZN(n488), 
	.A(n4736));
   OAI211_X1 U5667 (.ZN(n4736), 
	.C2(n1267), 
	.C1(n1261), 
	.B(n4737), 
	.A(n1953));
   NOR2_X1 U5668 (.ZN(n4737), 
	.A2(n4738), 
	.A1(n1220));
   NOR4_X1 U5669 (.ZN(n4738), 
	.A4(n469), 
	.A3(n1297), 
	.A2(n17098), 
	.A1(n721));
   NAND2_X1 U5670 (.ZN(n469), 
	.A2(n16657), 
	.A1(n16816));
   INV_X1 U5671 (.ZN(n721), 
	.A(n1021));
   NAND2_X1 U5672 (.ZN(n1021), 
	.A2(n16798), 
	.A1(n16801));
   NOR2_X1 U5674 (.ZN(n1220), 
	.A2(n16811), 
	.A1(n478));
   AOI21_X1 U5676 (.ZN(n1953), 
	.B2(n730), 
	.B1(n550), 
	.A(n1471));
   INV_X1 U5677 (.ZN(n1471), 
	.A(n738));
   NAND2_X1 U5678 (.ZN(n738), 
	.A2(n753), 
	.A1(n799));
   NAND4_X1 U5679 (.ZN(n753), 
	.A4(n4739), 
	.A3(n2599), 
	.A2(vis_pc_o[30]), 
	.A1(vis_pc_o[28]));
   NOR3_X1 U5680 (.ZN(n4739), 
	.A3(n4822), 
	.A2(n4817), 
	.A1(n4843));
   NAND4_X1 U5681 (.ZN(n2599), 
	.A4(n170), 
	.A3(n4348), 
	.A2(n191), 
	.A1(n4382));
   NOR2_X1 U5683 (.ZN(n4348), 
	.A2(vis_ipsr_o[4]), 
	.A1(vis_ipsr_o[5]));
   NOR2_X1 U5685 (.ZN(n4382), 
	.A2(vis_ipsr_o[0]), 
	.A1(vis_ipsr_o[2]));
   INV_X2 U5688 (.ZN(n799), 
	.A(n755));
   NAND2_X1 U5689 (.ZN(n755), 
	.A2(n16821), 
	.A1(n17097));
   INV_X1 U5691 (.ZN(n730), 
	.A(n1297));
   NAND2_X1 U5692 (.ZN(n1297), 
	.A2(n16804), 
	.A1(n708));
   INV_X1 U5693 (.ZN(n550), 
	.A(n582));
   NAND2_X1 U5694 (.ZN(n582), 
	.A2(n16817), 
	.A1(n16796));
   NAND2_X1 U5695 (.ZN(n1267), 
	.A2(n16804), 
	.A1(n4974));
   NAND2_X2 U5698 (.ZN(n692), 
	.A2(FE_OFN17_n16805), 
	.A1(n16828));
   INV_X4 U5699 (.ZN(n797), 
	.A(FE_OFN73_n16806));
   OAI221_X1 U5702 (.ZN(n4734), 
	.C2(n941), 
	.C1(n16811), 
	.B2(FE_OFN21_n503), 
	.B1(n4740), 
	.A(n4741));
   AOI22_X1 U5703 (.ZN(n4741), 
	.B2(n16816), 
	.B1(n4743), 
	.A2(n475), 
	.A1(n4742));
   INV_X1 U5704 (.ZN(n4743), 
	.A(n497));
   NAND2_X1 U5705 (.ZN(n497), 
	.A2(n1540), 
	.A1(n16797));
   INV_X1 U5706 (.ZN(n1540), 
	.A(n580));
   NAND2_X1 U5707 (.ZN(n580), 
	.A2(n16812), 
	.A1(n708));
   NAND2_X1 U5709 (.ZN(n1228), 
	.A2(n16659), 
	.A1(n16871));
   AOI21_X1 U5712 (.ZN(n4742), 
	.B2(n16799), 
	.B1(n729), 
	.A(n16870));
   INV_X1 U5713 (.ZN(n729), 
	.A(n625));
   NAND2_X1 U5714 (.ZN(n625), 
	.A2(n16807), 
	.A1(n16812));
   NOR3_X1 U5716 (.ZN(n4740), 
	.A3(n4745), 
	.A2(n629), 
	.A1(n4744));
   NOR3_X1 U5717 (.ZN(n4745), 
	.A3(n16813), 
	.A2(n16803), 
	.A1(n329));
   NAND2_X1 U5719 (.ZN(n329), 
	.A2(n16725), 
	.A1(n16871));
   INV_X1 U5721 (.ZN(n629), 
	.A(n1486));
   NAND2_X1 U5722 (.ZN(n1486), 
	.A2(n16803), 
	.A1(n822));
   OAI22_X1 U5723 (.ZN(n4744), 
	.B2(n17098), 
	.B1(n941), 
	.A2(n1261), 
	.A1(n731));
   NAND2_X1 U5725 (.ZN(n941), 
	.A2(n822), 
	.A1(n16812));
   INV_X1 U5726 (.ZN(n822), 
	.A(n1594));
   NAND2_X1 U5727 (.ZN(n1594), 
	.A2(n16871), 
	.A1(n16795));
   NAND2_X1 U5728 (.ZN(n1261), 
	.A2(n16871), 
	.A1(n16807));
   NAND2_X1 U5731 (.ZN(n1963), 
	.A2(n16817), 
	.A1(n16657));
   DFFR_X1 Nbm2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n5034), 
	.Q(n194), 
	.D(FE_PHN1682_n16735), 
	.CK(HCLK__L5_N5));
   DFFR_X2 Ypi3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4746), 
	.Q(sys_reset_req_o), 
	.D(FE_PHN1457_n5654), 
	.CK(HCLK__L5_N2));
   DFFS_X1 F2o2z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n260), 
	.Q(sub_2068_A_0_), 
	.D(FE_PHN3217_n5736), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Z8b3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n300), 
	.Q(sub_2068_A_6_), 
	.D(FE_PHN1396_n5730), 
	.CK(HCLK__L5_N2));
   DFFS_X1 W0b3z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n306), 
	.Q(sub_2068_A_3_), 
	.D(FE_PHN3654_n5733), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Qxa3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n302), 
	.Q(sub_2068_A_5_), 
	.D(FE_PHN1136_n5731), 
	.CK(HCLK__L5_N2));
   DFFS_X1 M2b3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n308), 
	.Q(sub_2068_A_2_), 
	.D(FE_PHN3585_n5734), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Gza3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n304), 
	.Q(sub_2068_A_4_), 
	.D(FE_PHN1137_n5732), 
	.CK(HCLK__L5_N2));
   DFFS_X1 C4b3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n310), 
	.Q(sub_2068_A_1_), 
	.D(FE_PHN3639_n5735), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Dhb3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n298), 
	.Q(sub_2068_A_7_), 
	.D(FE_PHN3078_n5729), 
	.CK(HCLK__L5_N13));
   DFFS_X1 M5f3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n296), 
	.Q(sub_2068_A_8_), 
	.D(FE_PHN3547_n5728), 
	.CK(HCLK__L5_N13));
   DFFS_X1 Aze3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n294), 
	.Q(sub_2068_A_9_), 
	.D(FE_PHN1398_n5727), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Zva3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n292), 
	.Q(sub_2068_A_10_), 
	.D(FE_PHN1130_n5726), 
	.CK(HCLK__L5_N13));
   DFFS_X1 Jca3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n262), 
	.D(FE_PHN5066_n5653), 
	.CK(HCLK__L5_N2));
   DFFS_X1 She3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n290), 
	.Q(sub_2068_A_11_), 
	.D(FE_PHN1397_n5725), 
	.CK(HCLK__L5_N13));
   DFFS_X1 Iua3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n288), 
	.Q(sub_2068_A_12_), 
	.D(FE_PHN1393_n5724), 
	.CK(HCLK__L5_N13));
   DFFS_X1 K7g3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n286), 
	.Q(sub_2068_A_13_), 
	.D(FE_PHN1399_n5723), 
	.CK(HCLK__L5_N13));
   DFFS_X1 Rsa3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n284), 
	.Q(sub_2068_A_14_), 
	.D(FE_PHN1135_n5722), 
	.CK(HCLK__L5_N13));
   DFFS_X1 Ara3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n282), 
	.Q(sub_2068_A_15_), 
	.D(FE_PHN1394_n5721), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Xeo2z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n280), 
	.Q(sub_2068_A_16_), 
	.D(FE_PHN1085_n5720), 
	.CK(HCLK__L5_N13));
   DFFS_X1 S3i3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n278), 
	.Q(sub_2068_A_17_), 
	.D(FE_PHN1395_n5719), 
	.CK(HCLK__L5_N5));
   DFFS_X1 O0o2z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n276), 
	.Q(sub_2068_A_18_), 
	.D(FE_PHN1131_n5718), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Jpa3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n274), 
	.Q(sub_2068_A_19_), 
	.D(FE_PHN3071_n5717), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Z2h3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n272), 
	.Q(sub_2068_A_20_), 
	.D(FE_PHN3544_n5716), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Ogo2z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n270), 
	.Q(sub_2068_A_21_), 
	.D(FE_PHN1138_n5715), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Ddi3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n268), 
	.Q(sub_2068_A_22_), 
	.D(FE_PHN1129_n5714), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Uei3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n264), 
	.Q(sub_2068_A_23_), 
	.D(FE_PHN3050_n5713), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Ufy2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n370), 
	.D(FE_PHN3133_n14432), 
	.CK(HCLK__L5_N5));
   DFFS_X1 T1y2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n1319), 
	.D(n14934), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Fey2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n335), 
	.D(FE_PHN972_n5755), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Y7y2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n6), 
	.D(FE_PHN2981_n5760), 
	.CK(HCLK__L5_N5));
   DFFS_X1 I3y2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n9), 
	.D(FE_PHN3200_n5763), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Bdm2z4_reg (.SN(FE_OFN174_HRESETn), 
	.QN(n2), 
	.D(FE_PHN3199_n5756), 
	.CK(HCLK__L5_N5));
   DFFS_X1 K6y2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n7), 
	.D(FE_PHN3094_n5761), 
	.CK(HCLK__L5_N5));
   DFFS_X1 W4y2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n8), 
	.D(FE_PHN3134_n5762), 
	.CK(HCLK__L5_N4));
   DFFS_X1 M9y2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n5), 
	.D(FE_PHN2972_n5759), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Bby2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4), 
	.D(FE_PHN801_n5758), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Qcy2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n3), 
	.D(FE_PHN2974_n5757), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Owq2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n164), 
	.Q(n4806), 
	.D(FE_PHN3142_n5765), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Lbn2z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n175), 
	.Q(n4804), 
	.D(FE_PHN3198_n5767), 
	.CK(HCLK__L5_N5));
   DFFS_X1 G0w2z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n191), 
	.Q(vis_ipsr_o[1]), 
	.D(FE_PHN731_n5691), 
	.CK(hclk));
   DFFS_X1 R1w2z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n186), 
	.Q(vis_ipsr_o[0]), 
	.D(FE_PHN4639_n5692), 
	.CK(hclk));
   DFFR_X1 I6w2z4_reg (.RN(FE_OFN175_HRESETn), 
	.QN(n184), 
	.D(FE_PHN1615_n5827), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Uic3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n3010), 
	.Q(n4799), 
	.D(FE_PHN2046_n5699), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Pab3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n1885), 
	.Q(n4753), 
	.D(FE_PHN4595_U791_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Fed3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n1896), 
	.Q(n4752), 
	.D(FE_PHN4580_U763_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 W5c3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n1411), 
	.D(FE_PHN1600_n13907), 
	.CK(HCLK__L5_N39));
   DFFR_X1 E9c3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n1447), 
	.D(FE_PHN1601_n13758), 
	.CK(HCLK__L5_N39));
   DFFR_X1 Zqb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n1310), 
	.D(FE_PHN1673_n14956), 
	.CK(HCLK__L5_N27));
   DFFR_X1 D4g3z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n244), 
	.D(FE_PHN2903_n5707), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Thm2z4_reg (.RN(FE_OFN159_HRESETn), 
	.QN(n1045), 
	.Q(vis_primask_o), 
	.D(FE_PHN1433_n5824), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Jje3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n4338), 
	.Q(n4755), 
	.D(n13846), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Wuq2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n3775), 
	.Q(n4751), 
	.D(n4897), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Uaj2z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n176), 
	.Q(vis_ipsr_o[2]), 
	.D(FE_PHN3474_n5689), 
	.CK(hclk));
   DFFR_X1 Cam2z4_reg (.RN(FE_OFN152_HRESETn), 
	.QN(n170), 
	.Q(vis_ipsr_o[3]), 
	.D(FE_PHN712_n5687), 
	.CK(hclk));
   DFFR_X1 Tdp2z4_reg (.RN(FE_OFN152_HRESETn), 
	.QN(n159), 
	.Q(vis_ipsr_o[5]), 
	.D(FE_PHN2926_n5683), 
	.CK(hclk));
   DFFR_X1 Trq2z4_reg (.RN(FE_OFN152_HRESETn), 
	.QN(n165), 
	.Q(vis_ipsr_o[4]), 
	.D(FE_PHN3282_n5685), 
	.CK(hclk));
   DFFR_X1 Idk2z4_reg (.RN(FE_OFN159_HRESETn), 
	.QN(n83), 
	.Q(vis_apsr_o[0]), 
	.D(FE_PHN3153_n5668), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Jcw2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n4847), 
	.D(FE_PHN1624_n4881), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Ydw2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4777), 
	.Q(n367), 
	.D(FE_PHN762_n4906), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Xuw2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4788), 
	.Q(n345), 
	.D(FE_PHN847_n4917), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Urw2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4786), 
	.Q(n349), 
	.D(FE_PHN2939_n4915), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Sow2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n4784), 
	.Q(n353), 
	.D(FE_PHN825_n4913), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Qzw2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n4791), 
	.Q(n339), 
	.D(FE_PHN851_n4920), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Qlw2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4782), 
	.Q(n357), 
	.D(FE_PHN821_n4911), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Oiw2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4780), 
	.Q(n361), 
	.D(FE_PHN2944_n4909), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Mww2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n4789), 
	.Q(n343), 
	.D(FE_PHN849_n4918), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Mfw2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4778), 
	.Q(n365), 
	.D(FE_PHN793_n4907), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Itw2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n4787), 
	.Q(n347), 
	.D(FE_PHN820_n4916), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Gqw2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n4785), 
	.Q(n351), 
	.D(FE_PHN823_n4914), 
	.CK(HCLK__L5_N4));
   DFFS_X1 F1x2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n4792), 
	.Q(n372), 
	.D(FE_PHN826_n4921), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Enw2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n4783), 
	.Q(n355), 
	.D(FE_PHN2943_n4912), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Ckw2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4781), 
	.Q(n359), 
	.D(FE_PHN822_n4910), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Byw2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4790), 
	.Q(n369), 
	.D(FE_PHN845_n4919), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Ahw2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n4779), 
	.Q(n363), 
	.D(FE_PHN824_n4908), 
	.CK(HCLK__L5_N5));
   DFFS_X1 M1j2z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n4968), 
	.Q(n3436), 
	.D(FE_PHN1488_U691_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 B2i3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n5639), 
	.D(FE_PHN4552_n4885), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Ieh3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n5625), 
	.D(FE_PHN4602_n4890), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Xyn2z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n5067), 
	.Q(n3250), 
	.D(n4888), 
	.CK(HCLK__L5_N5));
   DFFS_X1 I1h3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n5618), 
	.D(FE_PHN4383_n4891), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Mka3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n5514), 
	.Q(n3012), 
	.D(n4871), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Gdo2z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n5074), 
	.Q(n3381), 
	.D(n4892), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Gha3z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n5512), 
	.Q(n3227), 
	.D(FE_PHN4472_n4869), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Qfa3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n5511), 
	.Q(n3311), 
	.D(n4868), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Taa3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n5509), 
	.Q(n3056), 
	.D(n4867), 
	.CK(HCLK__L5_N2));
   DFFS_X1 L8m2z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n5033), 
	.Q(n3126), 
	.D(n4887), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Aea3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n5510), 
	.D(n4861), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Wia3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n5513), 
	.Q(n3104), 
	.D(FE_PHN4407_n4870), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Nfb3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n5520), 
	.D(FE_PHN4561_n4857), 
	.CK(HCLK__L5_N2));
   DFFS_X1 J7b3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n5517), 
	.Q(n2946), 
	.D(n4859), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Cma3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n5515), 
	.Q(n2881), 
	.D(n4855), 
	.CK(HCLK__L5_N13));
   DFFS_X1 Wzy2z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5252), 
	.Q(n3492), 
	.D(FE_PHN4324_U105_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Rni2z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n4959), 
	.Q(n3495), 
	.D(FE_PHN4571_U144_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Kxe3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n5579), 
	.Q(n3326), 
	.D(n4889), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Bge3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n5571), 
	.Q(n3111), 
	.D(FE_PHN4358_n4872), 
	.CK(HCLK__L5_N2));
   DFFS_X1 C9a3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n5508), 
	.Q(n3268), 
	.D(n4866), 
	.CK(HCLK__L5_N2));
   DFFS_X1 W3f3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n5581), 
	.D(FE_PHN4488_n4884), 
	.CK(HCLK__L5_N2));
   DFFS_X1 T5g3z4_reg (.SN(FE_OFN30_HRESETn), 
	.QN(n5600), 
	.Q(n2986), 
	.D(n4873), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Hxx2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n4845), 
	.Q(n1008), 
	.D(FE_PHN3070_n4879), 
	.CK(HCLK__L5_N3));
   DFFS_X1 D4a3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n5505), 
	.D(FE_PHN4550_n4856), 
	.CK(HCLK__L5_N2));
   DFFS_X1 U5a3z4_reg (.SN(FE_OFN28_HRESETn), 
	.QN(n5506), 
	.Q(n2917), 
	.D(n4858), 
	.CK(HCLK__L5_N2));
   DFFS_X1 L7a3z4_reg (.SN(FE_OFN55_HRESETn), 
	.QN(n5507), 
	.D(FE_PHN4431_n4865), 
	.CK(HCLK__L5_N2));
   DFFS_X1 Tyx2z4_reg (.SN(FE_OFN192_HRESETn), 
	.Q(n1009), 
	.D(FE_PHN1379_n5798), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Wai2z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n4947), 
	.Q(n1759), 
	.D(FE_PHN1906_n5800), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Yaz2z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5259), 
	.Q(n3493), 
	.D(FE_PHN3606_U98_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Svk2z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5004), 
	.Q(n3489), 
	.D(FE_PHN1967_U122_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 T1d3z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5544), 
	.Q(n3496), 
	.D(FE_PHN3576_U97_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 H3d3z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5545), 
	.Q(n1353), 
	.D(FE_PHN1970_U754_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 W7z2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n5257), 
	.Q(n2827), 
	.D(FE_PHN3755_n8706), 
	.CK(HCLK__L5_N3));
   DFFS_X1 K9z2z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n5258), 
	.Q(n2819), 
	.D(FE_PHN3690_n8698), 
	.CK(HCLK__L5_N9));
   DFFS_X1 I6z2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n5256), 
	.Q(n2865), 
	.D(FE_PHN1657_n5779), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Qzq2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n5120), 
	.Q(n2172), 
	.D(FE_PHN1648_U811_Z_0), 
	.CK(HCLK__L5_N3));
   DFFS_X1 I2t2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n5162), 
	.Q(n486), 
	.D(FE_PHN1571_n5771), 
	.CK(HCLK__L5_N3));
   DFFS_X1 C3z2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n5254), 
	.Q(n1723), 
	.D(FE_PHN4544_n5770), 
	.CK(HCLK__L5_N3));
   DFFS_X1 K1z2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n5253), 
	.Q(n2731), 
	.D(FE_PHN4541_n5772), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Auk2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n5003), 
	.Q(n2774), 
	.D(n5773), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Fzl2z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n5027), 
	.Q(n2231), 
	.D(FE_PHN3506_U795_Z_0), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Uup2z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n5100), 
	.Q(n795), 
	.D(FE_PHN3502_U755_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Iwp2z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5101), 
	.Q(n2188), 
	.D(FE_PHN3880_n5738), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Jw93z4_reg (.SN(FE_OFN152_HRESETn), 
	.QN(n5500), 
	.Q(n2620), 
	.D(FE_PHN1627_n5786), 
	.CK(hclk));
   DFFS_X1 U4z2z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n5255), 
	.Q(n2635), 
	.D(FE_PHN4126_n5776), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Xx93z4_reg (.SN(FE_OFN152_HRESETn), 
	.QN(n5501), 
	.Q(n2593), 
	.D(FE_PHN1629_n5784), 
	.CK(hclk));
   DFFS_X1 Ovc3z4_reg (.SN(FE_OFN152_HRESETn), 
	.QN(n4853), 
	.Q(n2570), 
	.D(FE_PHN1461_n4944), 
	.CK(hclk));
   DFFS_X1 Qdj2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n4974), 
	.Q(n503), 
	.D(FE_PHN4804_n14928), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Dvy2z4_reg (.SN(FE_OFN42_HRESETn), 
	.QN(n16818), 
	.Q(n16687), 
	.D(FE_PHN2918_n5742), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Rxl2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n5026), 
	.Q(n461), 
	.D(FE_PHN3090_n5751), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Viy2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n5241), 
	.Q(n454), 
	.D(FE_PHN2965_n5750), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Efp2z4_reg (.SN(FE_OFN152_HRESETn), 
	.QN(n4852), 
	.Q(n2539), 
	.D(FE_PHN1631_n4943), 
	.CK(hclk));
   DFFS_X1 U593z4_reg (.SN(FE_OFN195_HRESETn), 
	.Q(n1152), 
	.D(n4927), 
	.CK(hclk));
   DFFS_X1 I793z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n4828), 
	.Q(n2221), 
	.D(FE_PHN1983_n4923), 
	.CK(hclk));
   DFFS_X1 Szr2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4851), 
	.Q(n1161), 
	.D(n4940), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Rkd3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4771), 
	.Q(n3142), 
	.D(FE_PHN3277_n4939), 
	.CK(HCLK__L5_N25));
   DFFS_X1 G1s2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5140), 
	.Q(n869), 
	.D(FE_PHN3437_n5783), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Dkr2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4830), 
	.Q(n3028), 
	.D(FE_PHN3521_n4937), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Wce3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4831), 
	.Q(n3049), 
	.D(FE_PHN3536_n4938), 
	.CK(HCLK__L5_N26));
   DFFS_X1 G9w2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n5230), 
	.Q(n651), 
	.D(FE_PHN1905_n5828), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Slr2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n4832), 
	.Q(n2970), 
	.D(FE_PHN3518_n4936), 
	.CK(HCLK__L5_N25));
   DFFS_X1 J7q2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4850), 
	.Q(n2961), 
	.D(FE_PHN3519_n4935), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Y8q2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4827), 
	.Q(n1163), 
	.D(n4941), 
	.CK(HCLK__L5_N26));
   DFFS_X1 H4p2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4769), 
	.Q(n2817), 
	.D(FE_PHN3274_n4933), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Ym93z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4770), 
	.Q(n2841), 
	.D(FE_PHN3278_n4934), 
	.CK(HCLK__L5_N26));
   DFFS_X1 F0y2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n5240), 
	.Q(n403), 
	.D(FE_PHN1005_n5764), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Kyi2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n4966), 
	.Q(n413), 
	.D(FE_PHN3057_n5769), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Gtp2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n5099), 
	.Q(n415), 
	.D(FE_PHN2966_n5766), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Dwl2z4_reg (.SN(FE_OFN43_HRESETn), 
	.QN(n5025), 
	.D(FE_PHN3091_n5768), 
	.CK(HCLK__L5_N5));
   DFFS_X1 W5p2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4768), 
	.Q(n2795), 
	.D(FE_PHN1392_n4932), 
	.CK(HCLK__L5_N1));
   DFFS_X1 L7p2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4767), 
	.Q(n2772), 
	.D(FE_PHN3190_n4931), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Llq2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4765), 
	.Q(n2714), 
	.D(FE_PHN1177_n4929), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Tzg3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4766), 
	.Q(n2746), 
	.D(FE_PHN3276_n4930), 
	.CK(HCLK__L5_N1));
   DFFS_X1 G6d3z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n5546), 
	.D(FE_PHN4601_U317_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Zfh3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n4764), 
	.Q(n2713), 
	.D(FE_PHN3275_n4928), 
	.CK(HCLK__L5_N26));
   DFFS_X1 B6j2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n4772), 
	.Q(n2515), 
	.D(FE_PHN3516_n4942), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Q7j2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4971), 
	.Q(n2481), 
	.D(FE_PHN4584_n5737), 
	.CK(HCLK__L5_N25));
   DFFS_X1 S8k2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4762), 
	.Q(n2441), 
	.D(FE_PHN3520_n4925), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Lgi3z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4763), 
	.Q(n2460), 
	.D(FE_PHN3517_n4926), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Ohh3z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5626), 
	.Q(n2279), 
	.D(FE_PHN1490_n5787), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Hak2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4761), 
	.Q(n2280), 
	.D(FE_PHN3534_n4924), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Cqo2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4773), 
	.Q(n881), 
	.D(FE_PHN3072_n5788), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Rhi2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4955), 
	.Q(n874), 
	.D(FE_PHN1500_n5785), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Rbi3z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n4846), 
	.D(FE_PHN1429_n4945), 
	.CK(HCLK__L5_N3));
   DFFS_X1 V1l2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4774), 
	.Q(n867), 
	.D(FE_PHN3073_n5782), 
	.CK(HCLK__L5_N8));
   DFFR_X1 Nen2z4_reg (.RN(FE_OFN192_HRESETn), 
	.QN(n5055), 
	.Q(vis_control_o), 
	.D(FE_PHN1126_U692_Z_0), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Zei2z4_reg (.RN(FE_OFN159_HRESETn), 
	.QN(n4953), 
	.Q(vis_apsr_o[1]), 
	.D(FE_PHN1237_U809_Z_0), 
	.CK(HCLK__L5_N3));
   DFFR_X1 S4w2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n5228), 
	.Q(n596), 
	.D(n4880), 
	.CK(HCLK__L5_N3));
   DFFR_X1 J6i2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4905), 
	.Q(n251), 
	.D(FE_PHN3482_n5711), 
	.CK(hclk));
   DFFR_X1 Ffs2z4_reg (.RN(FE_OFN152_HRESETn), 
	.QN(n5149), 
	.Q(n1110), 
	.D(FE_PHN4829_n5791), 
	.CK(hclk));
   DFFR_X1 Lz93z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5502), 
	.Q(n4073), 
	.D(FE_PHN3477_n5790), 
	.CK(hclk));
   DFFS_X1 Zjq2z4_reg (.SN(FE_OFN194_HRESETn), 
	.QN(n5114), 
	.Q(vis_pc_o[18]), 
	.D(FE_PHN1463_n5665), 
	.CK(HCLK__L5_N1));
   DFFS_X1 Plx2z4_reg (.SN(FE_OFN29_HRESETn), 
	.QN(n5236), 
	.Q(vis_pc_o[16]), 
	.D(FE_PHN1195_n5663), 
	.CK(HCLK__L5_N1));
   DFFS_X1 Foe3z4_reg (.SN(FE_OFN194_HRESETn), 
	.QN(n5573), 
	.Q(vis_pc_o[20]), 
	.D(FE_PHN1462_n5660), 
	.CK(HCLK__L5_N1));
   DFFS_X1 Dkx2z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n5235), 
	.Q(vis_pc_o[15]), 
	.D(FE_PHN1196_n5664), 
	.CK(HCLK__L5_N1));
   DFFS_X1 Bnx2z4_reg (.SN(FE_OFN194_HRESETn), 
	.QN(n5237), 
	.Q(vis_pc_o[17]), 
	.D(FE_PHN1468_n5662), 
	.CK(HCLK__L5_N1));
   DFFS_X1 B9g3z4_reg (.SN(FE_OFN194_HRESETn), 
	.QN(n5601), 
	.Q(vis_pc_o[19]), 
	.D(FE_PHN1183_n5659), 
	.CK(HCLK__L5_N1));
   DFFS_X1 Rix2z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n4813), 
	.Q(vis_pc_o[13]), 
	.D(FE_PHN3405_n5677), 
	.CK(hclk));
   DFFS_X1 Gmd3z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n4815), 
	.Q(vis_pc_o[10]), 
	.D(FE_PHN3353_n5675), 
	.CK(hclk));
   DFFS_X1 Fhx2z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n4812), 
	.Q(vis_pc_o[11]), 
	.D(FE_PHN839_n5678), 
	.CK(hclk));
   DFFS_X1 V4d3z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n4814), 
	.Q(vis_pc_o[8]), 
	.D(FE_PHN3375_n5676), 
	.CK(hclk));
   DFFS_X1 Ycx2z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n4825), 
	.Q(vis_pc_o[6]), 
	.D(FE_PHN2976_n5656), 
	.CK(hclk));
   DFFS_X1 Nbx2z4_reg (.SN(FE_OFN152_HRESETn), 
	.Q(vis_pc_o[5]), 
	.D(FE_PHN741_n5681), 
	.CK(hclk));
   DFFS_X1 J4x2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n5233), 
	.Q(vis_pc_o[1]), 
	.D(n5688), 
	.CK(hclk));
   DFFS_X1 G7x2z4_reg (.SN(FE_OFN152_HRESETn), 
	.Q(vis_pc_o[2]), 
	.D(n5686), 
	.CK(hclk));
   DFFS_X1 Cax2z4_reg (.SN(FE_OFN152_HRESETn), 
	.Q(vis_pc_o[4]), 
	.D(FE_PHN3377_n5682), 
	.CK(hclk));
   DFFS_X1 R8x2z4_reg (.SN(FE_OFN152_HRESETn), 
	.Q(vis_pc_o[3]), 
	.D(FE_PHN3421_n5684), 
	.CK(hclk));
   DFFS_X1 Zjg3z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5608), 
	.Q(vis_r10_o[20]), 
	.D(U474_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Z523z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5325), 
	.Q(vis_r11_o[16]), 
	.D(FE_PHN3769_U407_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Y6o2z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5070), 
	.Q(vis_r5_o[16]), 
	.D(U409_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Wu53z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5410), 
	.Q(vis_r8_o[18]), 
	.D(U438_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Wrg3z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5613), 
	.Q(vis_r7_o[20]), 
	.D(FE_PHN2866_U479_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Vgg3z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5606), 
	.Q(vis_r8_o[20]), 
	.D(U472_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 V223z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5323), 
	.Q(vis_r11_o[18]), 
	.D(FE_PHN5039_U441_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Tvn2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5065), 
	.Q(vis_msp_o[16]), 
	.D(FE_PHN2851_U448_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Sog3z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5611), 
	.Q(vis_r5_o[20]), 
	.D(U477_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Skv2z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5218), 
	.Q(vis_r4_o[16]), 
	.D(U408_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Sg83z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5470), 
	.Q(vis_r2_o[16]), 
	.D(U402_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ro43z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5383), 
	.Q(vis_r9_o[16]), 
	.D(U405_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Rdg3z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5604), 
	.Q(vis_r2_o[20]), 
	.D(U470_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Rbo2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5073), 
	.Q(vis_psp_o[14]), 
	.D(U415_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Pwg3z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5616), 
	.Q(vis_msp_o[18]), 
	.D(U482_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Psn2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5063), 
	.Q(vis_r5_o[18]), 
	.D(U443_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Olg3z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5609), 
	.Q(vis_r11_o[20]), 
	.D(FE_PHN2847_U475_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Ohv2z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5216), 
	.Q(vis_r4_o[18]), 
	.D(U442_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Od83z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5468), 
	.Q(vis_r2_o[18]), 
	.D(U436_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 O403z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5278), 
	.Q(vis_r12_o[16]), 
	.D(U412_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Nl43z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5381), 
	.Q(vis_r9_o[18]), 
	.D(U439_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Nag3z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5602), 
	.Q(vis_r0_o[20]), 
	.D(U468_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 N8o2z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5071), 
	.Q(vis_r7_o[16]), 
	.D(FE_PHN2848_U411_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ltg3z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5614), 
	.Q(vis_r12_o[20]), 
	.D(U480_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Kig3z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5607), 
	.Q(vis_r9_o[20]), 
	.D(U473_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 K103z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5276), 
	.Q(vis_r12_o[18]), 
	.D(U446_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Jl93z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5494), 
	.Q(vis_r0_o[16]), 
	.D(U400_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Jbu2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5189), 
	.Q(vis_r6_o[16]), 
	.D(U410_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 J773z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5441), 
	.Q(vis_r3_o[16]), 
	.D(U403_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 J5o2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5069), 
	.Q(vis_r1_o[16]), 
	.D(U401_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Ixn2z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5066), 
	.Q(vis_psp_o[16]), 
	.D(U449_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 If33z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5354), 
	.Q(vis_r10_o[16]), 
	.D(U406_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 I113z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5299), 
	.Q(vis_r14_o[16]), 
	.D(U413_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Hqg3z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5612), 
	.Q(vis_r6_o[20]), 
	.D(U478_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Gfg3z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5605), 
	.Q(vis_r3_o[20]), 
	.D(FE_PHN2819_U471_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Fi93z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5492), 
	.Q(vis_r0_o[18]), 
	.D(U434_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 F473z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5439), 
	.Q(vis_r3_o[18]), 
	.D(U437_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 F8u2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5187), 
	.Q(vis_r6_o[18]), 
	.D(U444_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Eyg3z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5617), 
	.Q(vis_psp_o[18]), 
	.D(U483_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Ey03z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5297), 
	.Q(vis_r14_o[18]), 
	.D(U447_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Eun2z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5064), 
	.Q(vis_r7_o[18]), 
	.D(FE_PHN2809_U445_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ec33z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5352), 
	.Q(vis_r10_o[18]), 
	.D(U440_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Dng3z4_reg (.SN(FE_OFN164_HRESETn), 
	.QN(n5610), 
	.Q(vis_r4_o[20]), 
	.D(U476_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Ccg3z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5603), 
	.Q(vis_r1_o[20]), 
	.D(U469_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Cao2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5072), 
	.Q(vis_msp_o[14]), 
	.D(U414_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Ay53z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5412), 
	.Q(vis_r8_o[16]), 
	.D(U404_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Avg3z4_reg (.SN(FE_OFN166_HRESETn), 
	.QN(n5615), 
	.Q(vis_r14_o[20]), 
	.D(FE_PHN2795_U481_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Arn2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5062), 
	.Q(vis_r1_o[18]), 
	.D(U435_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Zxo2z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5084), 
	.Q(vis_r5_o[17]), 
	.D(U427_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Zfv2z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5215), 
	.Q(vis_r4_o[19]), 
	.D(U460_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Zb83z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5467), 
	.Q(vis_r2_o[19]), 
	.D(FE_PHN2805_U454_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Z203z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5277), 
	.Q(vis_r12_o[17]), 
	.D(U430_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Yj43z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5380), 
	.Q(vis_r9_o[19]), 
	.D(U457_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Xyh3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5637), 
	.Q(vis_msp_o[17]), 
	.D(FE_PHN2835_U466_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Uj93z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5493), 
	.Q(vis_r0_o[17]), 
	.D(U418_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 U573z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5440), 
	.Q(vis_r3_o[17]), 
	.D(U421_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 U9u2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5188), 
	.Q(vis_r6_o[17]), 
	.D(FE_PHN2824_U428_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Tz03z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5298), 
	.Q(vis_r14_o[17]), 
	.D(U431_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Tvh3z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5635), 
	.Q(vis_r12_o[19]), 
	.D(U464_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Td33z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5353), 
	.Q(vis_r10_o[17]), 
	.D(U424_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 S2p2z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5087), 
	.Q(vis_psp_o[15]), 
	.D(U433_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Qg93z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5491), 
	.Q(vis_r0_o[19]), 
	.D(U452_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Q273z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5438), 
	.Q(vis_r3_o[19]), 
	.D(U455_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Q6u2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5186), 
	.Q(vis_r6_o[19]), 
	.D(U462_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Pap2z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5089), 
	.Q(vis_r5_o[19]), 
	.D(U461_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Pa33z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5351), 
	.Q(vis_r10_o[19]), 
	.D(U458_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Ozo2z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5085), 
	.Q(vis_r7_o[17]), 
	.D(FE_PHN2864_U429_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 M0i3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5638), 
	.Q(vis_psp_o[17]), 
	.D(U467_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Lw53z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5411), 
	.Q(vis_r8_o[17]), 
	.D(U422_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Kwo2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5083), 
	.Q(vis_r1_o[17]), 
	.D(U419_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 K423z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5324), 
	.Q(vis_r11_o[17]), 
	.D(FE_PHN3814_U425_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Ixh3z4_reg (.SN(FE_OFN165_HRESETn), 
	.QN(n5636), 
	.Q(vis_r14_o[19]), 
	.D(U465_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Ht53z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5409), 
	.Q(vis_r8_o[19]), 
	.D(U456_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 G123z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5322), 
	.Q(vis_r11_o[19]), 
	.D(FE_PHN2873_U459_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Ecp2z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5090), 
	.Q(vis_r7_o[19]), 
	.D(FE_PHN3733_U463_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Djv2z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5217), 
	.Q(vis_r4_o[17]), 
	.D(U426_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Df83z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5469), 
	.Q(vis_r2_o[17]), 
	.D(U420_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 D1p2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5086), 
	.Q(vis_msp_o[15]), 
	.D(U432_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Cn43z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5382), 
	.Q(vis_r9_o[17]), 
	.D(U423_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 A9p2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5088), 
	.Q(vis_r1_o[19]), 
	.D(FE_PHN3582_U453_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Nox2z4_reg (.SN(FE_OFN194_HRESETn), 
	.QN(n5238), 
	.Q(vis_pc_o[21]), 
	.D(FE_PHN1086_n5661), 
	.CK(HCLK__L5_N1));
   DFFS_X1 Tch3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5624), 
	.Q(vis_psp_o[19]), 
	.D(U501_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Sr53z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5408), 
	.Q(vis_r8_o[21]), 
	.D(FE_PHN2815_U490_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Rz13z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5321), 
	.Q(vis_r11_o[21]), 
	.D(FE_PHN3647_U493_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Poq2z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5116), 
	.Q(vis_r5_o[21]), 
	.D(U495_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 P9h3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5622), 
	.Q(vis_r14_o[21]), 
	.D(U499_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Kev2z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5214), 
	.Q(vis_r4_o[21]), 
	.D(U494_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Ka83z4_reg (.SN(FE_OFN163_HRESETn), 
	.QN(n5466), 
	.Q(vis_r2_o[21]), 
	.D(U488_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Ji43z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5379), 
	.Q(vis_r9_o[21]), 
	.D(U491_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Eqq2z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5117), 
	.Q(vis_r7_o[21]), 
	.D(FE_PHN3730_U497_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ebh3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5623), 
	.Q(vis_msp_o[19]), 
	.D(FE_PHN2794_U500_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Bf93z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5490), 
	.Q(vis_r0_o[21]), 
	.D(U486_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 B173z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5437), 
	.Q(vis_r3_o[21]), 
	.D(U489_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 B5u2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5185), 
	.Q(vis_r6_o[21]), 
	.D(FE_PHN2802_U496_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Anq2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5115), 
	.Q(vis_r1_o[21]), 
	.D(U487_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 A933z4_reg (.SN(FE_OFN167_HRESETn), 
	.QN(n5350), 
	.Q(vis_r10_o[21]), 
	.D(U492_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 A8h3z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5621), 
	.Q(vis_r12_o[21]), 
	.D(U498_Z_0), 
	.CK(HCLK__L5_N22));
   DFFS_X1 Kaf3z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n4824), 
	.Q(vis_pc_o[22]), 
	.D(FE_PHN749_n5657), 
	.CK(hclk));
   DFFS_X1 Tme3z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n4816), 
	.Q(vis_pc_o[12]), 
	.D(FE_PHN941_n5674), 
	.CK(hclk));
   DFFS_X1 Ufx2z4_reg (.SN(FE_OFN195_HRESETn), 
	.QN(n4811), 
	.Q(vis_pc_o[9]), 
	.D(FE_PHN3414_n5679), 
	.CK(hclk));
   DFFS_X1 Jwf3z4_reg (.SN(FE_OFN195_HRESETn), 
	.Q(vis_pc_o[14]), 
	.D(FE_PHN3084_n5658), 
	.CK(HCLK__L5_N1));
   DFFS_X1 Jex2z4_reg (.SN(FE_OFN195_HRESETn), 
	.Q(vis_pc_o[7]), 
	.D(FE_PHN939_n5680), 
	.CK(hclk));
   DFFS_X1 W5s2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5143), 
	.Q(vis_r7_o[9]), 
	.D(FE_PHN2829_U295_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Uku2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5195), 
	.Q(vis_r6_o[9]), 
	.D(U294_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ug73z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5447), 
	.Q(vis_r3_o[9]), 
	.D(U287_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 U2s2z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5141), 
	.Q(vis_r1_o[9]), 
	.D(U285_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Tse3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5576), 
	.Q(vis_msp_o[7]), 
	.D(U298_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 To33z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5360), 
	.Q(vis_r10_o[9]), 
	.D(U290_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Rpe3z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5574), 
	.Q(vis_r12_o[9]), 
	.D(U296_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 L763z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5418), 
	.Q(vis_r8_o[9]), 
	.D(U288_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Kf23z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5331), 
	.Q(vis_r11_o[9]), 
	.D(FE_PHN2843_U291_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 I4s2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5142), 
	.Q(vis_r5_o[9]), 
	.D(U293_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Hue3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5577), 
	.Q(vis_psp_o[7]), 
	.D(U299_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Fre3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5575), 
	.Q(vis_r14_o[9]), 
	.D(U297_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Duv2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5224), 
	.Q(vis_r4_o[9]), 
	.D(U292_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Dq83z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5476), 
	.Q(vis_r2_o[9]), 
	.D(U286_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Cy43z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5389), 
	.Q(vis_r9_o[9]), 
	.D(U289_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Cxc3z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5541), 
	.Q(vis_r0_o[9]), 
	.D(U284_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Zgr2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5130), 
	.Q(vis_msp_o[10]), 
	.D(U366_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Vdr2z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5128), 
	.Q(vis_r5_o[12]), 
	.D(U361_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 T263z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5415), 
	.Q(vis_r8_o[12]), 
	.D(U356_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Sa23z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5328), 
	.Q(vis_r11_o[12]), 
	.D(FE_PHN2858_U359_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 S703z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5280), 
	.Q(vis_r12_o[12]), 
	.D(U364_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Rr93z4_reg (.SN(FE_OFN177_HRESETn), 
	.QN(n5497), 
	.Q(vis_r0_o[12]), 
	.D(U352_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Oir2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5131), 
	.Q(vis_psp_o[10]), 
	.D(U367_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 M413z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5301), 
	.Q(vis_r14_o[12]), 
	.D(U365_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Lpv2z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5221), 
	.Q(vis_r4_o[12]), 
	.D(U360_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ll83z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5473), 
	.Q(vis_r2_o[12]), 
	.D(U354_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Kt43z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5386), 
	.Q(vis_r9_o[12]), 
	.D(U357_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Kfr2z4_reg (.SN(FE_OFN177_HRESETn), 
	.QN(n5129), 
	.Q(vis_r7_o[12]), 
	.D(FE_PHN5026_U363_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Gcr2z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5127), 
	.Q(vis_r1_o[12]), 
	.D(FE_PHN3878_U353_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Cgu2z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5192), 
	.Q(vis_r6_o[12]), 
	.D(U362_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Cc73z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5444), 
	.Q(vis_r3_o[12]), 
	.D(U355_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Bk33z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5357), 
	.Q(vis_r10_o[12]), 
	.D(U358_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Y1n2z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5049), 
	.Q(vis_r5_o[22]), 
	.D(U511_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Vzz2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5275), 
	.Q(vis_r12_o[22]), 
	.D(U514_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Vcv2z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5213), 
	.Q(vis_r4_o[22]), 
	.D(U510_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 V883z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5465), 
	.Q(vis_r2_o[22]), 
	.D(FE_PHN2822_U504_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ug43z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5378), 
	.Q(vis_r9_o[22]), 
	.D(U507_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 R6n2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5052), 
	.Q(vis_psp_o[20]), 
	.D(U517_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Pw03z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5296), 
	.Q(vis_r14_o[22]), 
	.D(U515_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 N3n2z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5050), 
	.Q(vis_r7_o[22]), 
	.D(FE_PHN4897_U513_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Mz63z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5436), 
	.Q(vis_r3_o[22]), 
	.D(U505_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Md93z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5489), 
	.Q(vis_r0_o[22]), 
	.D(U502_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 M3u2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5184), 
	.Q(vis_r6_o[22]), 
	.D(U512_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 L733z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5349), 
	.Q(vis_r10_o[22]), 
	.D(U508_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 J0n2z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5048), 
	.Q(vis_r1_o[22]), 
	.D(FE_PHN2827_U503_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Dq53z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5407), 
	.Q(vis_r8_o[22]), 
	.D(FE_PHN2853_U506_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Cy13z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5320), 
	.Q(vis_r11_o[22]), 
	.D(FE_PHN2854_U509_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 C5n2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5051), 
	.Q(vis_msp_o[20]), 
	.D(U516_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Z853z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5396), 
	.Q(vis_r8_o[0]), 
	.D(U738_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Yg13z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5309), 
	.Q(vis_r11_o[0]), 
	.D(U723_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Unm2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5040), 
	.Q(vis_r0_o[0]), 
	.D(U803_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Skm2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5038), 
	.Q(vis_r7_o[0]), 
	.D(FE_PHN2799_U708_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Rvu2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5202), 
	.Q(vis_r4_o[0]), 
	.D(U693_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Rr73z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5454), 
	.Q(vis_r2_o[0]), 
	.D(FE_PHN2798_U748_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Qz33z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5367), 
	.Q(vis_r9_o[0]), 
	.D(U733_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Knz2z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5267), 
	.Q(vis_r12_o[0]), 
	.D(U713_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Imt2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5173), 
	.Q(vis_r6_o[0]), 
	.D(U703_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Ii63z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5425), 
	.Q(vis_r3_o[0]), 
	.D(FE_PHN2804_U743_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Hq23z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5338), 
	.Q(vis_r10_o[0]), 
	.D(FE_PHN2811_U728_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Gmm2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5039), 
	.Q(vis_r1_o[0]), 
	.D(U797_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Ek03z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5288), 
	.Q(vis_r14_o[0]), 
	.D(U718_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Ejm2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5037), 
	.Q(vis_r5_o[0]), 
	.D(U698_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Yfn2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5056), 
	.Q(vis_r1_o[2]), 
	.D(FE_PHN2141_U301_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 X563z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5417), 
	.Q(vis_r8_o[2]), 
	.D(FE_PHN2061_U304_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Wd23z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5330), 
	.Q(vis_r11_o[2]), 
	.D(FE_PHN2090_U307_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Wa03z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5282), 
	.Q(vis_r12_o[2]), 
	.D(FE_PHN2078_U312_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Vu93z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5499), 
	.Q(vis_r0_o[2]), 
	.D(FE_PHN2107_U300_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Q713z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5303), 
	.Q(vis_r14_o[2]), 
	.D(FE_PHN1743_U313_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Psv2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5223), 
	.Q(vis_r4_o[2]), 
	.D(FE_PHN2064_U308_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Po83z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5475), 
	.Q(vis_r2_o[2]), 
	.D(FE_PHN2154_U302_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Ow43z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5388), 
	.Q(vis_r9_o[2]), 
	.D(FE_PHN3527_U305_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Okn2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5059), 
	.Q(vis_msp_o[0]), 
	.D(FE_PHN2103_U314_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Mhn2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5057), 
	.Q(vis_r5_o[2]), 
	.D(FE_PHN3529_U309_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Gju2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5194), 
	.Q(vis_r6_o[2]), 
	.D(FE_PHN2150_U310_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Gf73z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5446), 
	.Q(vis_r3_o[2]), 
	.D(FE_PHN2145_U303_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Fn33z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5359), 
	.Q(vis_r10_o[2]), 
	.D(FE_PHN2094_U306_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Cmn2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5060), 
	.Q(vis_psp_o[0]), 
	.D(FE_PHN2053_U315_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Ajn2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5058), 
	.Q(vis_r7_o[2]), 
	.D(FE_PHN2156_U311_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Z7i2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n4922), 
	.Q(vis_tbit_o), 
	.D(FE_PHN774_n14825), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Yx63z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5435), 
	.Q(vis_r3_o[3]), 
	.D(U522_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Yb93z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5488), 
	.Q(vis_r0_o[3]), 
	.D(FE_PHN3541_U519_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Y1u2z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5183), 
	.Q(vis_r6_o[3]), 
	.D(U529_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 X533z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5348), 
	.Q(vis_r10_o[3]), 
	.D(U525_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 X6m2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5032), 
	.Q(vis_psp_o[1]), 
	.D(FE_PHN2092_U534_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 V3m2z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5030), 
	.Q(vis_r7_o[3]), 
	.D(U530_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 T0m2z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5028), 
	.Q(vis_r1_o[3]), 
	.D(U520_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Po53z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5406), 
	.Q(vis_r8_o[3]), 
	.D(FE_PHN2079_U523_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Ow13z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5319), 
	.Q(vis_r11_o[3]), 
	.D(U526_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 J5m2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5031), 
	.Q(vis_msp_o[1]), 
	.D(FE_PHN2054_U533_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Hyz2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5274), 
	.Q(vis_r12_o[3]), 
	.D(FE_PHN1744_U531_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Hbv2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5212), 
	.Q(vis_r4_o[3]), 
	.D(U527_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 H783z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5464), 
	.Q(vis_r2_o[3]), 
	.D(U521_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 H2m2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5029), 
	.Q(vis_r5_o[3]), 
	.D(FE_PHN3532_U528_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Gf43z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5377), 
	.Q(vis_r9_o[3]), 
	.D(FE_PHN2104_U524_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Bv03z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5295), 
	.Q(vis_r14_o[3]), 
	.D(FE_PHN2082_U532_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Zr03z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5293), 
	.Q(vis_r14_o[5]), 
	.D(FE_PHN2076_U564_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Wyt2z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5181), 
	.Q(vis_r6_o[5]), 
	.D(U561_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Wu63z4_reg (.SN(FE_OFN180_HRESETn), 
	.QN(n5433), 
	.Q(vis_r3_o[5]), 
	.D(U554_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Wmp2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5095), 
	.Q(vis_psp_o[3]), 
	.D(FE_PHN3526_U566_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 W893z4_reg (.SN(FE_OFN178_HRESETn), 
	.QN(n5486), 
	.Q(vis_r0_o[5]), 
	.D(U551_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 V233z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5346), 
	.Q(vis_r10_o[5]), 
	.D(FE_PHN3528_U557_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Ujp2z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5093), 
	.Q(vis_r7_o[5]), 
	.D(U562_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Sgp2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5091), 
	.Q(vis_r1_o[5]), 
	.D(U552_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Nl53z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5404), 
	.Q(vis_r8_o[5]), 
	.D(FE_PHN2077_U555_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Mt13z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5317), 
	.Q(vis_r11_o[5]), 
	.D(U558_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Ilp2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5094), 
	.Q(vis_msp_o[3]), 
	.D(FE_PHN2089_U565_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Gip2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5092), 
	.Q(vis_r5_o[5]), 
	.D(U560_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Fvz2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5272), 
	.Q(vis_r12_o[5]), 
	.D(FE_PHN3524_U563_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 F483z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5462), 
	.Q(vis_r2_o[5]), 
	.D(U553_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 F8v2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5210), 
	.Q(vis_r4_o[5]), 
	.D(U559_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Ec43z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5375), 
	.Q(vis_r9_o[5]), 
	.D(FE_PHN2065_U556_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 U5r2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5124), 
	.Q(vis_msp_o[2]), 
	.D(U549_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Twz2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5273), 
	.Q(vis_r12_o[4]), 
	.D(U547_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 T583z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5463), 
	.Q(vis_r2_o[4]), 
	.D(U537_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 T9v2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5211), 
	.Q(vis_r4_o[4]), 
	.D(U543_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Sd43z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5376), 
	.Q(vis_r9_o[4]), 
	.D(U540_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 S2r2z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5122), 
	.Q(vis_r5_o[4]), 
	.D(U544_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Nt03z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5294), 
	.Q(vis_r14_o[4]), 
	.D(U548_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Kw63z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5434), 
	.Q(vis_r3_o[4]), 
	.D(U538_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Ka93z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5487), 
	.Q(vis_r0_o[4]), 
	.D(U535_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 K0u2z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5182), 
	.Q(vis_r6_o[4]), 
	.D(U545_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 J433z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5347), 
	.Q(vis_r10_o[4]), 
	.D(U541_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 I7r2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5125), 
	.Q(vis_psp_o[2]), 
	.D(U550_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 G4r2z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5123), 
	.Q(vis_r7_o[4]), 
	.D(U546_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 E1r2z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5121), 
	.Q(vis_r1_o[4]), 
	.D(U536_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Bn53z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5405), 
	.Q(vis_r8_o[4]), 
	.D(U539_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Av13z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5318), 
	.Q(vis_r11_o[4]), 
	.D(U542_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Zu43z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5387), 
	.Q(vis_r9_o[10]), 
	.D(FE_PHN3522_U323_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Z8s2z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5145), 
	.Q(vis_r5_o[10]), 
	.D(FE_PHN2083_U327_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Rhu2z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5193), 
	.Q(vis_r6_o[10]), 
	.D(FE_PHN2157_U328_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Rds2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5148), 
	.Q(vis_psp_o[8]), 
	.D(FE_PHN2075_U333_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Rd73z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5445), 
	.Q(vis_r3_o[10]), 
	.D(FE_PHN3539_U321_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ql33z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5358), 
	.Q(vis_r10_o[10]), 
	.D(FE_PHN3525_U324_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Oas2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5146), 
	.Q(vis_r7_o[10]), 
	.D(FE_PHN2286_U329_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 K7s2z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5144), 
	.Q(vis_r1_o[10]), 
	.D(FE_PHN3546_U319_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 I463z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5416), 
	.Q(vis_r8_o[10]), 
	.D(FE_PHN2120_U322_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Hc23z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5329), 
	.Q(vis_r11_o[10]), 
	.D(FE_PHN2294_U325_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 H903z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5281), 
	.Q(vis_r12_o[10]), 
	.D(FE_PHN2068_U330_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Gt93z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5498), 
	.Q(vis_r0_o[10]), 
	.D(FE_PHN3523_U318_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Dcs2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5147), 
	.Q(vis_msp_o[8]), 
	.D(FE_PHN2163_U332_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 B613z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5302), 
	.Q(vis_r14_o[10]), 
	.D(FE_PHN2102_U331_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Arv2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5222), 
	.Q(vis_r4_o[10]), 
	.D(FE_PHN2096_U326_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 An83z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5474), 
	.Q(vis_r2_o[10]), 
	.D(FE_PHN3573_U320_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Xyk2z4_reg (.SN(FE_OFN152_HRESETn), 
	.Q(vis_pc_o[23]), 
	.D(n5672), 
	.CK(hclk));
   DFFS_X1 Wnu2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5197), 
	.Q(vis_r6_o[15]), 
	.D(U260_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Wj73z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5449), 
	.Q(vis_r3_o[15]), 
	.D(U253_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Vr33z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5362), 
	.Q(vis_r10_o[15]), 
	.D(U256_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Rdq2z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5110), 
	.Q(vis_r7_o[15]), 
	.D(FE_PHN2872_U261_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Psh3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5633), 
	.Q(vis_msp_o[13]), 
	.D(U264_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 Naq2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5108), 
	.Q(vis_r1_o[15]), 
	.D(U251_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Na63z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5420), 
	.Q(vis_r8_o[15]), 
	.D(U254_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Mi23z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5333), 
	.Q(vis_r11_o[15]), 
	.D(FE_PHN2836_U257_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Lph3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5631), 
	.Q(vis_r12_o[15]), 
	.D(U262_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Fxv2z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5226), 
	.Q(vis_r4_o[15]), 
	.D(U258_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ft83z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5478), 
	.Q(vis_r2_o[15]), 
	.D(U252_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Euh3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5634), 
	.Q(vis_psp_o[13]), 
	.D(U265_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 E153z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5391), 
	.Q(vis_r9_o[15]), 
	.D(U255_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 E0d3z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5543), 
	.Q(vis_r0_o[15]), 
	.D(U250_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ccq2z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5109), 
	.Q(vis_r5_o[15]), 
	.D(U259_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Arh3z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5632), 
	.Q(vis_r14_o[15]), 
	.D(FE_PHN2823_U263_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Z863z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5419), 
	.Q(vis_r8_o[8]), 
	.D(U272_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Yg23z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5332), 
	.Q(vis_r11_o[8]), 
	.D(FE_PHN2861_U275_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Rvv2z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5225), 
	.Q(vis_r4_o[8]), 
	.D(U276_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Rr83z4_reg (.SN(FE_OFN68_HRESETn), 
	.QN(n5477), 
	.Q(vis_r2_o[8]), 
	.D(U270_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Qz43z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5390), 
	.Q(vis_r9_o[8]), 
	.D(U273_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Qyc3z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5542), 
	.Q(vis_r0_o[8]), 
	.D(U268_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Qwr2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5138), 
	.Q(vis_msp_o[6]), 
	.D(U282_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Otr2z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5136), 
	.Q(vis_r5_o[8]), 
	.D(U277_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Kc03z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5283), 
	.Q(vis_r12_o[8]), 
	.D(U280_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Imu2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5196), 
	.Q(vis_r6_o[8]), 
	.D(U278_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Ii73z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5448), 
	.Q(vis_r3_o[8]), 
	.D(U271_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Hq33z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5361), 
	.Q(vis_r10_o[8]), 
	.D(U274_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Eyr2z4_reg (.SN(FE_OFN48_HRESETn), 
	.QN(n5139), 
	.Q(vis_psp_o[6]), 
	.D(U283_Z_0), 
	.CK(HCLK__L5_N26));
   DFFS_X1 E913z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5304), 
	.Q(vis_r14_o[8]), 
	.D(U281_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Cvr2z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5137), 
	.Q(vis_r7_o[8]), 
	.D(FE_PHN2869_U279_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Asr2z4_reg (.SN(FE_OFN49_HRESETn), 
	.QN(n5135), 
	.Q(vis_r1_o[8]), 
	.D(U269_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Fcj2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n4973), 
	.Q(vis_pc_o[0]), 
	.D(FE_PHN1024_n5690), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Zj53z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5403), 
	.Q(vis_r8_o[6]), 
	.D(U571_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Ytm2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5044), 
	.Q(vis_msp_o[4]), 
	.D(U581_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Yr13z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5316), 
	.Q(vis_r11_o[6]), 
	.D(U574_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Wqm2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5042), 
	.Q(vis_r5_o[6]), 
	.D(U576_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Rtz2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5271), 
	.Q(vis_r12_o[6]), 
	.D(U579_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 R283z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5461), 
	.Q(vis_r2_o[6]), 
	.D(U569_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 R6v2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5209), 
	.Q(vis_r4_o[6]), 
	.D(U575_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Qa43z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5374), 
	.Q(vis_r9_o[6]), 
	.D(U572_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Mvm2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5045), 
	.Q(vis_psp_o[4]), 
	.D(U582_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Lq03z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5292), 
	.Q(vis_r14_o[6]), 
	.D(U580_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Ksm2z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5043), 
	.Q(vis_r7_o[6]), 
	.D(U578_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Ixt2z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5180), 
	.Q(vis_r6_o[6]), 
	.D(U577_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 It63z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5432), 
	.Q(vis_r3_o[6]), 
	.D(U570_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Ipm2z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5041), 
	.Q(vis_r1_o[6]), 
	.D(U568_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 H133z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5345), 
	.Q(vis_r10_o[6]), 
	.D(U573_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 G493z4_reg (.SN(FE_OFN179_HRESETn), 
	.QN(n5485), 
	.Q(vis_r0_o[6]), 
	.D(U567_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 X553z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5394), 
	.Q(vis_r8_o[7]), 
	.D(U740_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Wd13z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5307), 
	.Q(vis_r11_o[7]), 
	.D(U725_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Spl2z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5021), 
	.Q(vis_r1_o[7]), 
	.D(U799_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Qml2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5019), 
	.Q(vis_r5_o[7]), 
	.D(U700_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Psu2z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5200), 
	.Q(vis_r4_o[7]), 
	.D(U695_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Po73z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5452), 
	.Q(vis_r2_o[7]), 
	.D(U750_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Ow33z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5365), 
	.Q(vis_r9_o[7]), 
	.D(U735_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Mcz2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5260), 
	.Q(vis_psp_o[5]), 
	.D(U687_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Ikz2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5265), 
	.Q(vis_r12_o[7]), 
	.D(U715_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Grl2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5022), 
	.Q(vis_r0_o[7]), 
	.D(U804_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Gjt2z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n5171), 
	.Q(vis_r6_o[7]), 
	.D(U705_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Gf63z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5423), 
	.Q(vis_r3_o[7]), 
	.D(FE_PHN2807_U745_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Fn23z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5336), 
	.Q(vis_r10_o[7]), 
	.D(U730_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Eol2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5020), 
	.Q(vis_r7_o[7]), 
	.D(U710_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Cll2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5018), 
	.Q(vis_msp_o[5]), 
	.D(U684_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Ch03z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5286), 
	.Q(vis_r14_o[7]), 
	.D(U720_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Ycu2z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5190), 
	.Q(vis_r6_o[14]), 
	.D(U394_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Y873z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5442), 
	.Q(vis_r3_o[14]), 
	.D(U387_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Xg33z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5355), 
	.Q(vis_r10_o[14]), 
	.D(U390_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 X213z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5300), 
	.Q(vis_r14_o[14]), 
	.D(U397_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 U5q2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5107), 
	.Q(vis_psp_o[12]), 
	.D(U399_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Q2q2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5105), 
	.Q(vis_r7_o[14]), 
	.D(FE_PHN2856_U395_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Pz53z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5413), 
	.Q(vis_r8_o[14]), 
	.D(U388_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 O723z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5326), 
	.Q(vis_r11_o[14]), 
	.D(FE_PHN2813_U391_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 No93z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5495), 
	.Q(vis_r0_o[14]), 
	.D(U384_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Mzp2z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5103), 
	.Q(vis_r1_o[14]), 
	.D(U385_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Hmv2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5219), 
	.Q(vis_r4_o[14]), 
	.D(U392_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Hi83z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5471), 
	.Q(vis_r2_o[14]), 
	.D(FE_PHN2828_U386_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Gq43z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5384), 
	.Q(vis_r9_o[14]), 
	.D(U389_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 F4q2z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5106), 
	.Q(vis_msp_o[12]), 
	.D(U398_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 D603z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5279), 
	.Q(vis_r12_o[14]), 
	.D(U396_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 B1q2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5104), 
	.Q(vis_r5_o[14]), 
	.D(U393_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Wlz2z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5266), 
	.Q(vis_r12_o[1]), 
	.D(U714_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Ukt2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5172), 
	.Q(vis_r6_o[1]), 
	.D(U704_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Ug63z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5424), 
	.Q(vis_r3_o[1]), 
	.D(U744_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Txj2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n4987), 
	.Q(vis_r0_o[1]), 
	.D(U810_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 To23z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5337), 
	.Q(vis_r10_o[1]), 
	.D(U729_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Ruj2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n4985), 
	.Q(vis_r7_o[1]), 
	.D(U709_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Qi03z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5287), 
	.Q(vis_r14_o[1]), 
	.D(U719_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 L753z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5395), 
	.Q(vis_r8_o[1]), 
	.D(U739_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Kf13z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5308), 
	.Q(vis_r11_o[1]), 
	.D(U724_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Fwj2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n4986), 
	.Q(vis_r1_o[1]), 
	.D(U798_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Duu2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5201), 
	.Q(vis_r4_o[1]), 
	.D(U694_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Dtj2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n4984), 
	.Q(vis_r5_o[1]), 
	.D(U699_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Dq73z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5453), 
	.Q(vis_r2_o[1]), 
	.D(U749_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Cy33z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5366), 
	.Q(vis_r9_o[1]), 
	.D(U734_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Xmf3z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5590), 
	.Q(vis_r4_o[23]), 
	.D(FE_PHN2073_U240_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Wbf3z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5583), 
	.Q(vis_r0_o[23]), 
	.D(FE_PHN2091_U232_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Uuf3z4_reg (.SN(FE_OFN184_HRESETn), 
	.QN(n5595), 
	.Q(vis_psp_o[21]), 
	.D(FE_PHN3535_U247_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Tjf3z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5588), 
	.Q(vis_r10_o[23]), 
	.D(FE_PHN2084_U238_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Qrf3z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5593), 
	.Q(vis_r12_o[23]), 
	.D(FE_PHN2052_U244_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Mof3z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5591), 
	.Q(vis_r5_o[23]), 
	.D(FE_PHN2055_U241_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Eif3z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5587), 
	.Q(vis_r9_o[23]), 
	.D(FE_PHN2071_U237_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Orj2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n4983), 
	.Q(vis_r1_o[23]), 
	.D(FE_PHN2212_U233_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Ftf3z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5594), 
	.Q(vis_r14_o[23]), 
	.D(FE_PHN2196_U245_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Pgf3z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5586), 
	.Q(vis_r8_o[23]), 
	.D(FE_PHN2125_U236_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 M4j2z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n4970), 
	.Q(vis_msp_o[21]), 
	.D(FE_PHN3552_U246_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Ilf3z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5589), 
	.Q(vis_r11_o[23]), 
	.D(FE_PHN2300_U239_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Aff3z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5585), 
	.Q(vis_r3_o[23]), 
	.D(FE_PHN3540_U235_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Bqf3z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5592), 
	.Q(vis_r6_o[23]), 
	.D(FE_PHN2215_U242_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Ldf3z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5584), 
	.Q(vis_r2_o[23]), 
	.D(FE_PHN2241_U234_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Fpi2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n4960), 
	.Q(vis_r7_o[23]), 
	.D(FE_PHN2346_U243_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Zpx2z4_reg (.SN(FE_OFN152_HRESETn), 
	.QN(n4819), 
	.Q(vis_pc_o[24]), 
	.D(FE_PHN963_n5671), 
	.CK(hclk));
   DFFS_X1 X1e3z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5563), 
	.Q(vis_r5_o[11]), 
	.D(U343_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Wqd3z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5556), 
	.Q(vis_r2_o[11]), 
	.D(U336_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 U9e3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5568), 
	.Q(vis_msp_o[9]), 
	.D(U348_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Tyd3z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5561), 
	.Q(vis_r11_o[11]), 
	.D(FE_PHN3636_U341_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Snd3z4_reg (.SN(FE_OFN177_HRESETn), 
	.QN(n5554), 
	.Q(vis_r0_o[11]), 
	.D(U334_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Q6e3z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5566), 
	.Q(vis_r12_o[11]), 
	.D(U346_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Pvd3z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5559), 
	.Q(vis_r9_o[11]), 
	.D(U339_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 M3e3z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5564), 
	.Q(vis_r6_o[11]), 
	.D(U344_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Lsd3z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5557), 
	.Q(vis_r3_o[11]), 
	.D(U337_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Ibe3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5569), 
	.Q(vis_psp_o[9]), 
	.D(U349_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 I0e3z4_reg (.SN(FE_OFN135_HRESETn), 
	.QN(n5562), 
	.Q(vis_r4_o[11]), 
	.D(U342_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 Hpd3z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5555), 
	.Q(vis_r1_o[11]), 
	.D(FE_PHN3799_U335_Z_0), 
	.CK(HCLK__L5_N20));
   DFFS_X1 F8e3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5567), 
	.Q(vis_r14_o[11]), 
	.D(U347_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Exd3z4_reg (.SN(FE_OFN190_HRESETn), 
	.QN(n5560), 
	.Q(vis_r10_o[11]), 
	.D(U340_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 B5e3z4_reg (.SN(FE_OFN177_HRESETn), 
	.QN(n5565), 
	.Q(vis_r7_o[11]), 
	.D(FE_PHN3865_U345_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Aud3z4_reg (.SN(FE_OFN60_HRESETn), 
	.QN(n5558), 
	.Q(vis_r8_o[11]), 
	.D(U338_Z_0), 
	.CK(HCLK__L5_N24));
   DFFS_X1 Z0g3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5598), 
	.Q(vis_msp_o[11]), 
	.D(U382_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Wor2z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5133), 
	.Q(vis_r5_o[13]), 
	.D(U377_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Wnv2z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5220), 
	.Q(vis_r4_o[13]), 
	.D(U376_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Wj83z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5472), 
	.Q(vis_r2_o[13]), 
	.D(U370_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Vxf3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5596), 
	.Q(vis_r12_o[13]), 
	.D(U380_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Vr43z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5385), 
	.Q(vis_r9_o[13]), 
	.D(U373_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 O2g3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5599), 
	.Q(vis_psp_o[11]), 
	.D(U383_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Neu2z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5191), 
	.Q(vis_r6_o[13]), 
	.D(U378_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Na73z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5443), 
	.Q(vis_r3_o[13]), 
	.D(U371_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Mi33z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5356), 
	.Q(vis_r10_o[13]), 
	.D(U374_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Lqr2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5134), 
	.Q(vis_r7_o[13]), 
	.D(U379_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Kzf3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5597), 
	.Q(vis_r14_o[13]), 
	.D(U381_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Hnr2z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5132), 
	.Q(vis_r1_o[13]), 
	.D(U369_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 E163z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5414), 
	.Q(vis_r8_o[13]), 
	.D(U372_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 D923z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5327), 
	.Q(vis_r11_o[13]), 
	.D(U375_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Cq93z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5496), 
	.Q(vis_r0_o[13]), 
	.D(U368_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 Zpj2z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n4982), 
	.Q(vis_r1_o[24]), 
	.D(FE_PHN2181_U584_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Vmj2z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n4980), 
	.Q(vis_r5_o[24]), 
	.D(FE_PHN2100_U592_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Umi3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5646), 
	.Q(vis_msp_o[22]), 
	.D(FE_PHN3542_U597_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Tvt2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5179), 
	.Q(vis_r6_o[24]), 
	.D(FE_PHN2200_U593_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Tr63z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5431), 
	.Q(vis_r3_o[24]), 
	.D(FE_PHN3545_U586_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Sz23z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5344), 
	.Q(vis_r10_o[24]), 
	.D(FE_PHN3530_U589_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 R293z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n5484), 
	.Q(vis_r0_o[24]), 
	.D(FE_PHN3533_U583_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Qji3z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5644), 
	.Q(vis_r12_o[24]), 
	.D(FE_PHN3531_U595_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Ki53z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5402), 
	.Q(vis_r8_o[24]), 
	.D(FE_PHN2098_U587_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Jq13z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5315), 
	.Q(vis_r11_o[24]), 
	.D(FE_PHN1846_U590_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Joi3z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5647), 
	.Q(vis_psp_o[22]), 
	.D(FE_PHN2063_U598_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 Fli3z4_reg (.SN(FE_OFN33_HRESETn), 
	.QN(n5645), 
	.Q(vis_r14_o[24]), 
	.D(FE_PHN2166_U596_Z_0), 
	.CK(HCLK__L5_N25));
   DFFS_X1 F9j2z4_reg (.SN(FE_OFN41_HRESETn), 
	.QN(n4972), 
	.Q(vis_r7_o[24]), 
	.D(FE_PHN3725_U594_Z_0), 
	.CK(HCLK__L5_N19));
   DFFS_X1 C183z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5460), 
	.Q(vis_r2_o[24]), 
	.D(FE_PHN2219_U585_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 C5v2z4_reg (.SN(FE_OFN145_HRESETn), 
	.QN(n5208), 
	.Q(vis_r4_o[24]), 
	.D(FE_PHN3537_U591_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 B943z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5373), 
	.Q(vis_r9_o[24]), 
	.D(FE_PHN2067_U588_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Lrx2z4_reg (.SN(FE_OFN152_HRESETn), 
	.QN(n4820), 
	.Q(vis_pc_o[25]), 
	.D(FE_PHN813_n5670), 
	.CK(hclk));
   DFFS_X1 Xhl2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5016), 
	.Q(vis_psp_o[23]), 
	.D(U614_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Wo03z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5291), 
	.Q(vis_r14_o[25]), 
	.D(FE_PHN2814_U612_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Vg53z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5401), 
	.Q(vis_r8_o[25]), 
	.D(U603_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Uo13z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5314), 
	.Q(vis_r11_o[25]), 
	.D(FE_PHN2863_U606_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Tel2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5014), 
	.Q(vis_r7_o[25]), 
	.D(FE_PHN3744_U610_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Pbl2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5012), 
	.Q(vis_r1_o[25]), 
	.D(U600_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Nz73z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5459), 
	.Q(vis_r2_o[25]), 
	.D(U601_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 N3v2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5207), 
	.Q(vis_r4_o[25]), 
	.D(U607_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 M743z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5372), 
	.Q(vis_r9_o[25]), 
	.D(U604_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Igl2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5015), 
	.Q(vis_msp_o[23]), 
	.D(U613_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Eut2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5178), 
	.Q(vis_r6_o[25]), 
	.D(U609_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Eq63z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5430), 
	.Q(vis_r3_o[25]), 
	.D(U602_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Edl2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5013), 
	.Q(vis_r5_o[25]), 
	.D(U608_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Dy23z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5343), 
	.Q(vis_r10_o[25]), 
	.D(U605_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Csz2z4_reg (.SN(FE_OFN185_HRESETn), 
	.QN(n5270), 
	.Q(vis_r12_o[25]), 
	.D(U611_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 C193z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5483), 
	.Q(vis_r0_o[25]), 
	.D(U599_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Xsx2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n4821), 
	.Q(vis_pc_o[26]), 
	.D(FE_PHN779_n5669), 
	.CK(hclk));
   DFFS_X1 Z3k2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n4991), 
	.Q(vis_r7_o[26]), 
	.D(FE_PHN2224_U628_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Yx73z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5458), 
	.Q(vis_r2_o[26]), 
	.D(FE_PHN2225_U619_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Y1v2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5206), 
	.Q(vis_r4_o[26]), 
	.D(FE_PHN2070_U625_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 X543z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5371), 
	.Q(vis_r9_o[26]), 
	.D(FE_PHN2080_U622_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 V0k2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n4989), 
	.Q(vis_r1_o[26]), 
	.D(FE_PHN2187_U618_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Pst2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5177), 
	.Q(vis_r6_o[26]), 
	.D(FE_PHN3548_U627_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Po63z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5429), 
	.Q(vis_r3_o[26]), 
	.D(FE_PHN2189_U620_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Ow23z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5342), 
	.Q(vis_r10_o[26]), 
	.D(FE_PHN2081_U623_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 O5k2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4992), 
	.Q(vis_msp_o[24]), 
	.D(FE_PHN2143_U631_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Nz83z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5482), 
	.Q(vis_r0_o[26]), 
	.D(FE_PHN2087_U617_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Nqz2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5269), 
	.Q(vis_r12_o[26]), 
	.D(FE_PHN2095_U629_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 K2k2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n4990), 
	.Q(vis_r5_o[26]), 
	.D(FE_PHN2097_U626_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Hn03z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5290), 
	.Q(vis_r14_o[26]), 
	.D(FE_PHN3561_U630_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Gf53z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5400), 
	.Q(vis_r8_o[26]), 
	.D(FE_PHN2149_U621_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Fn13z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5313), 
	.Q(vis_r11_o[26]), 
	.D(FE_PHN2233_U624_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 D7k2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4993), 
	.Q(vis_psp_o[24]), 
	.D(FE_PHN3538_U632_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Jux2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n4822), 
	.Q(vis_pc_o[27]), 
	.D(FE_PHN1063_n5667), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Aez2z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5261), 
	.Q(vis_psp_o[26]), 
	.D(U686_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Zu33z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5364), 
	.Q(vis_r9_o[28]), 
	.D(U736_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Zkk2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n4998), 
	.Q(vis_r0_o[28]), 
	.D(U806_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Tiz2z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5264), 
	.Q(vis_r12_o[28]), 
	.D(U716_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Ql23z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5335), 
	.Q(vis_r10_o[28]), 
	.D(U731_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Ggk2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n4995), 
	.Q(vis_r5_o[28]), 
	.D(U701_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Aru2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5199), 
	.Q(vis_r4_o[28]), 
	.D(U696_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Nf03z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5285), 
	.Q(vis_r14_o[28]), 
	.D(FE_PHN3597_U721_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Kjk2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n4997), 
	.Q(vis_r1_o[28]), 
	.D(FE_PHN4986_U800_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Rek2z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n4994), 
	.Q(vis_msp_o[26]), 
	.D(FE_PHN2812_U683_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Rd63z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5422), 
	.Q(vis_r3_o[28]), 
	.D(U746_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 I453z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5393), 
	.Q(vis_r8_o[28]), 
	.D(U741_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Hc13z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5306), 
	.Q(vis_r11_o[28]), 
	.D(FE_PHN2859_U726_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Rht2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5170), 
	.Q(vis_r6_o[28]), 
	.D(U706_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 An73z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5451), 
	.Q(vis_r2_o[28]), 
	.D(U751_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Vhk2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n4996), 
	.Q(vis_r7_o[28]), 
	.D(FE_PHN2830_U711_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Zu23z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5341), 
	.Q(vis_r10_o[27]), 
	.D(U639_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Yx83z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5481), 
	.Q(vis_r0_o[27]), 
	.D(U633_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Wnh3z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5630), 
	.Q(vis_psp_o[25]), 
	.D(U648_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Vgq2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5112), 
	.Q(vis_r5_o[27]), 
	.D(U642_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Skh3z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5628), 
	.Q(vis_r14_o[27]), 
	.D(FE_PHN2820_U646_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Rd53z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5399), 
	.Q(vis_r8_o[27]), 
	.D(U637_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Ql13z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5312), 
	.Q(vis_r11_o[27]), 
	.D(U640_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Kiq2z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5113), 
	.Q(vis_r7_o[27]), 
	.D(FE_PHN2831_U644_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Jw73z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5457), 
	.Q(vis_r2_o[27]), 
	.D(U635_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 J0v2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5205), 
	.Q(vis_r4_o[27]), 
	.D(U641_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 I443z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5370), 
	.Q(vis_r9_o[27]), 
	.D(U638_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Hmh3z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5629), 
	.Q(vis_msp_o[25]), 
	.D(U647_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Gfq2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5111), 
	.Q(vis_r1_o[27]), 
	.D(FE_PHN2792_U634_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Djh3z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5627), 
	.Q(vis_r12_o[27]), 
	.D(U645_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Art2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5176), 
	.Q(vis_r6_o[27]), 
	.D(U643_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 An63z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5428), 
	.Q(vis_r3_o[27]), 
	.D(U636_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Vvx2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n5239), 
	.Q(vis_pc_o[28]), 
	.D(FE_PHN760_n5666), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Omk2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n4817), 
	.Q(vis_pc_o[29]), 
	.D(FE_PHN3391_n5673), 
	.CK(HCLK__L5_N3));
   DFFS_X1 J0l2z4_reg (.SN(FE_OFN192_HRESETn), 
	.QN(n5006), 
	.Q(vis_pc_o[30]), 
	.D(FE_PHN3387_n5655), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Y6i3z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5641), 
	.Q(vis_r14_o[30]), 
	.D(U679_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Wnt2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5174), 
	.Q(vis_r6_o[30]), 
	.D(U676_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Wj63z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5426), 
	.Q(vis_r3_o[30]), 
	.D(U669_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Vuo2z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5082), 
	.Q(vis_r7_o[30]), 
	.D(FE_PHN2821_U677_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Vr23z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5339), 
	.Q(vis_r10_o[30]), 
	.D(U672_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Uu83z4_reg (.SN(FE_OFN139_HRESETn), 
	.QN(n5479), 
	.Q(vis_r0_o[30]), 
	.D(U666_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Rro2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5080), 
	.Q(vis_r1_o[30]), 
	.D(FE_PHN4857_U667_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Na53z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5397), 
	.Q(vis_r8_o[30]), 
	.D(U670_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 N8i3z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5642), 
	.Q(vis_msp_o[28]), 
	.D(FE_PHN2806_U680_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Mi13z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5310), 
	.Q(vis_r11_o[30]), 
	.D(FE_PHN2845_U673_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 J5i3z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5640), 
	.Q(vis_r12_o[30]), 
	.D(U678_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Gto2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5081), 
	.Q(vis_r5_o[30]), 
	.D(U675_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Fxu2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5203), 
	.Q(vis_r4_o[30]), 
	.D(U674_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Ft73z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5455), 
	.Q(vis_r2_o[30]), 
	.D(U668_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 E143z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5368), 
	.Q(vis_r9_o[30]), 
	.D(U671_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Cai3z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5643), 
	.Q(vis_psp_o[28]), 
	.D(U681_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Yoz2z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5268), 
	.Q(vis_r12_o[29]), 
	.D(U661_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Ymo2z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5078), 
	.Q(vis_msp_o[27]), 
	.D(FE_PHN2810_U663_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Uyu2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5204), 
	.Q(vis_r4_o[29]), 
	.D(U657_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Uu73z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5456), 
	.Q(vis_r2_o[29]), 
	.D(FE_PHN2808_U651_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Ujo2z4_reg (.SN(FE_OFN182_HRESETn), 
	.QN(n5076), 
	.Q(vis_r5_o[29]), 
	.D(U658_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 T243z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5369), 
	.Q(vis_r9_o[29]), 
	.D(U654_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Sl03z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5289), 
	.Q(vis_r14_o[29]), 
	.D(U662_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Noo2z4_reg (.SN(FE_OFN61_HRESETn), 
	.QN(n5079), 
	.Q(vis_psp_o[27]), 
	.D(U664_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Lpt2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5175), 
	.Q(vis_r6_o[29]), 
	.D(U659_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Ll63z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5427), 
	.Q(vis_r3_o[29]), 
	.D(U652_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Kt23z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5340), 
	.Q(vis_r10_o[29]), 
	.D(U655_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Jw83z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5480), 
	.Q(vis_r0_o[29]), 
	.D(U649_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Jlo2z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5077), 
	.Q(vis_r7_o[29]), 
	.D(FE_PHN2852_U660_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Fio2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5075), 
	.Q(vis_r1_o[29]), 
	.D(U650_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Cc53z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5398), 
	.Q(vis_r8_o[29]), 
	.D(U653_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Bk13z4_reg (.SN(FE_OFN181_HRESETn), 
	.QN(n5311), 
	.Q(vis_r11_o[29]), 
	.D(FE_PHN2793_U656_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Yd03z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5284), 
	.Q(vis_r14_o[31]), 
	.D(U722_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Xti2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n4963), 
	.Q(vis_r0_o[31]), 
	.D(U805_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 X2j2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n4969), 
	.Q(vis_msp_o[29]), 
	.D(U682_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 T253z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5392), 
	.Q(vis_r8_o[31]), 
	.D(U742_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Sa13z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5305), 
	.Q(vis_r11_o[31]), 
	.D(FE_PHN2833_U727_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Pfz2z4_reg (.SN(FE_OFN38_HRESETn), 
	.QN(n5262), 
	.Q(vis_psp_o[29]), 
	.D(U685_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Lpu2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n5198), 
	.Q(vis_r4_o[31]), 
	.D(U697_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Ll73z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5450), 
	.Q(vis_r2_o[31]), 
	.D(U752_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Kt33z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5363), 
	.Q(vis_r9_o[31]), 
	.D(U737_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Koj2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n4981), 
	.Q(vis_r1_o[31]), 
	.D(FE_PHN2839_U801_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Isi2z4_reg (.SN(FE_OFN138_HRESETn), 
	.QN(n4962), 
	.Q(vis_r7_o[31]), 
	.D(FE_PHN2834_U712_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Glj2z4_reg (.SN(FE_OFN65_HRESETn), 
	.QN(n4979), 
	.Q(vis_r5_o[31]), 
	.D(U702_Z_0), 
	.CK(HCLK__L5_N7));
   DFFS_X1 Ehz2z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5263), 
	.Q(vis_r12_o[31]), 
	.D(U717_Z_0), 
	.CK(HCLK__L5_N23));
   DFFS_X1 Cgt2z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5169), 
	.Q(vis_r6_o[31]), 
	.D(U707_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Cc63z4_reg (.SN(FE_OFN66_HRESETn), 
	.QN(n5421), 
	.Q(vis_r3_o[31]), 
	.D(U747_Z_0), 
	.CK(HCLK__L5_N21));
   DFFS_X1 Bk23z4_reg (.SN(FE_OFN40_HRESETn), 
	.QN(n5334), 
	.Q(vis_r10_o[31]), 
	.D(U732_Z_0), 
	.CK(HCLK__L5_N8));
   DFFS_X1 Gci2z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n4948), 
	.Q(vis_apsr_o[3]), 
	.D(FE_PHN1241_U229_Z_0), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Igi2z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n4954), 
	.Q(vis_apsr_o[2]), 
	.D(FE_PHN1614_U665_Z_0), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Pet2z4_reg (.RN(FE_OFN192_HRESETn), 
	.QN(n4843), 
	.Q(n2029), 
	.D(FE_PHN1636_n4878), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Y6t2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n5165), 
	.Q(n808), 
	.D(FE_PHN1390_n4876), 
	.CK(HCLK__L5_N4));
   DFFR_X1 V3o2z4_reg (.RN(FE_OFN30_HRESETn), 
	.QN(n5068), 
	.D(FE_PHN3206_n5712), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Y9t2z4_reg (.RN(FE_OFN175_HRESETn), 
	.QN(n5167), 
	.Q(n1063), 
	.D(FE_PHN1610_n4886), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Mbt2z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n4829), 
	.Q(n3229), 
	.D(FE_PHN1625_n4864), 
	.CK(HCLK__L5_N2));
   DFFR_X1 S5b3z4_reg (.RN(FE_OFN192_HRESETn), 
	.QN(n4833), 
	.D(FE_PHN1809_n4874), 
	.CK(HCLK__L5_N2));
   DFFR_X1 R0t2z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n4848), 
	.Q(n3313), 
	.D(FE_PHN2086_n4882), 
	.CK(hclk));
   DFFR_X1 Adt2z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n5168), 
	.Q(n3059), 
	.D(FE_PHN2164_n4863), 
	.CK(hclk));
   DFFR_X1 Tna3z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n5516), 
	.D(FE_PHN1655_n4860), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Bec3z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n4801), 
	.Q(n217), 
	.D(n5696), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Zad3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5549), 
	.Q(n3847), 
	.D(FE_PHN4303_U766_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Bmb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5523), 
	.D(FE_PHN4394_U774_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Kkb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5522), 
	.Q(n3812), 
	.D(FE_PHN2886_U782_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Tib3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5521), 
	.Q(n3784), 
	.D(U790_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Mcc3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5535), 
	.Q(n214), 
	.D(n5695), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Fhc3z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n4800), 
	.Q(n223), 
	.D(n5698), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Ztc3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5540), 
	.D(FE_PHN4611_n5710), 
	.CK(HCLK__L5_N27));
   DFFR_X1 U5x2z4_reg (.RN(FE_OFN175_HRESETn), 
	.QN(n5234), 
	.D(FE_PHN1172_n5826), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Qfc3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5536), 
	.Q(n220), 
	.D(n5697), 
	.CK(HCLK__L5_N2));
   DFFR_X1 X9n2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4826), 
	.Q(n2889), 
	.D(FE_PHN2865_n4854), 
	.CK(hclk));
   DFFR_X1 Ylc3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4797), 
	.Q(n231), 
	.D(n5701), 
	.CK(HCLK__L5_N2));
   DFFR_X1 J9d3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5548), 
	.Q(n2951), 
	.D(U767_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Xdb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5519), 
	.Q(n2952), 
	.D(FE_PHN2882_U775_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Gcb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5518), 
	.D(FE_PHN2885_U783_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 G8n2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5053), 
	.Q(n4367), 
	.D(FE_PHN2887_U771_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Bus2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5158), 
	.Q(n2888), 
	.D(FE_PHN2817_U779_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Dks2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5152), 
	.Q(n2890), 
	.D(FE_PHN2878_U787_Z_0), 
	.CK(hclk));
   DFFR_X1 Jkc3z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n4798), 
	.Q(n228), 
	.D(n5700), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Uqi2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4961), 
	.Q(n3731), 
	.D(FE_PHN2420_n5652), 
	.CK(hclk));
   DFFR_X1 Aqp2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5097), 
	.Q(n2929), 
	.D(n4883), 
	.CK(hclk));
   DFFR_X1 B1a3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5503), 
	.D(FE_PHN2889_n4862), 
	.CK(hclk));
   DFFR_X1 Vfd3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5551), 
	.Q(n3834), 
	.D(FE_PHN2896_U762_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Z4l2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5008), 
	.Q(n3863), 
	.D(FE_PHN2875_U770_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Svs2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5159), 
	.Q(n3793), 
	.D(U778_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Uls2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5153), 
	.Q(n3790), 
	.D(FE_PHN2877_U786_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Lns2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5154), 
	.Q(n2927), 
	.D(FE_PHN2837_U785_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Lhd3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5552), 
	.Q(n2933), 
	.D(FE_PHN2849_U761_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Q6l2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5009), 
	.Q(n2931), 
	.D(FE_PHN2803_U769_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Jxs2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5160), 
	.Q(n2932), 
	.D(FE_PHN2841_U777_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Wbk2z4_reg (.RN(FE_OFN152_HRESETn), 
	.QN(n4802), 
	.Q(n209), 
	.D(FE_PHN2050_n5694), 
	.CK(hclk));
   DFFR_X1 Yvb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5527), 
	.D(FE_PHN1674_n13951), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Qsb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5525), 
	.D(FE_PHN1672_n13963), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Vve3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5578), 
	.D(FE_PHN2902_n5703), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Rnb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5524), 
	.D(FE_PHN1669_n13894), 
	.CK(HCLK__L5_N39));
   DFFR_X1 T7d3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5547), 
	.Q(n3719), 
	.D(FE_PHN4441_U764_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Usl2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5023), 
	.Q(n3720), 
	.D(FE_PHN2884_U772_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Tqs2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5156), 
	.Q(n3813), 
	.D(FE_PHN2870_U780_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Vgs2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5150), 
	.Q(n4356), 
	.D(FE_PHN2881_U788_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Pcd3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5550), 
	.Q(n2901), 
	.D(U765_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Axm2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5046), 
	.Q(n2902), 
	.D(U773_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Kss2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5157), 
	.D(FE_PHN2894_U781_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Mis2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5151), 
	.D(FE_PHN2893_U789_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Lee3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5570), 
	.D(FE_PHN2888_n5705), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Gzb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5529), 
	.D(FE_PHN1670_n13932), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Hzj2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4988), 
	.Q(n203), 
	.D(n5693), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Aok2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16844), 
	.Q(n16846), 
	.D(n10055), 
	.CK(HCLK__L5_N9));
   DFFR_X1 Nnc3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5537), 
	.D(FE_PHN2892_n5704), 
	.CK(HCLK__L5_N2));
   DFFR_X1 H2f3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n4796), 
	.D(FE_PHN4562_n5702), 
	.CK(HCLK__L5_N27));
   DFFR_X1 N7c3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5533), 
	.Q(n3861), 
	.D(n11945), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Pxb3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5528), 
	.Q(n3238), 
	.D(n4894), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Jsc3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5539), 
	.Q(n3785), 
	.D(n5709), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Vac3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5534), 
	.D(n11939), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Tqc3z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n5538), 
	.Q(n2916), 
	.D(n5708), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Dpc3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n4795), 
	.D(FE_PHN4585_n5706), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Gxk2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5005), 
	.D(n11929), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Hub3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5526), 
	.Q(n3107), 
	.D(n4893), 
	.CK(HCLK__L5_N27));
   DFFR_X1 O2c3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5531), 
	.D(FE_PHN1666_n13919), 
	.CK(HCLK__L5_N39));
   DFFR_X1 Ipb3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n4750), 
	.Q(n3060), 
	.D(n4901), 
	.CK(HCLK__L5_N27));
   DFFR_X1 X0c3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5530), 
	.D(n4899), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Q0f3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5580), 
	.Q(n1129), 
	.D(n4904), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Qnn2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5061), 
	.D(FE_PHN1602_n13835), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Etq2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5118), 
	.D(FE_PHN1667_n13989), 
	.CK(HCLK__L5_N27));
   DFFR_X1 C7f3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5582), 
	.D(FE_PHN1603_n13813), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Fij2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16850), 
	.Q(n16852), 
	.D(FE_PHN1612_n5781), 
	.CK(HCLK__L5_N9));
   DFFR_X1 W8r2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5126), 
	.Q(n4333), 
	.D(FE_PHN1606_n13795), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Uyv2z4_reg (.RN(FE_OFN152_HRESETn), 
	.Q(n1053), 
	.D(n5825), 
	.CK(hclk));
   DFFR_X1 F4c3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5532), 
	.Q(n2953), 
	.D(n4898), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Qrp2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5098), 
	.Q(n3740), 
	.D(FE_PHN2891_n5651), 
	.CK(hclk));
   DFFR_X1 Cps2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5155), 
	.Q(n3791), 
	.D(FE_PHN2832_U784_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Bjd3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5553), 
	.Q(n3833), 
	.D(U760_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 H8l2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5010), 
	.Q(n3862), 
	.D(U768_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 Azs2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5161), 
	.Q(n3792), 
	.D(U776_Z_0), 
	.CK(HCLK__L5_N1));
   DFFR_X1 P2a3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5504), 
	.Q(n3732), 
	.D(FE_PHN2818_n5650), 
	.CK(hclk));
   DFFR_X1 Nsk2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16827), 
	.Q(n16690), 
	.D(n9796), 
	.CK(HCLK__L5_N9));
   DFFR_X1 Npk2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16840), 
	.Q(n16728), 
	.D(n9972), 
	.CK(HCLK__L5_N9));
   DFFR_X1 Oar2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4749), 
	.Q(n3089), 
	.D(n4900), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Y9l2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5011), 
	.D(n11957), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Ble3z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5572), 
	.D(n11971), 
	.CK(HCLK__L5_N27));
   DFFR_X1 I6h3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5620), 
	.Q(n1379), 
	.D(FE_PHN1425_n14001), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Mvi2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4964), 
	.D(FE_PHN1671_n13870), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Ipn2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4748), 
	.D(FE_PHN1902_n4903), 
	.CK(HCLK__L5_N27));
   DFFR_X1 T8f3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n4747), 
	.D(FE_PHN1901_n4902), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Lul2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5024), 
	.Q(n3786), 
	.D(FE_PHN3001_n4895), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Rym2z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5047), 
	.Q(n2914), 
	.D(FE_PHN1364_n4896), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Ywi2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n4965), 
	.Q(n1066), 
	.D(FE_PHN3048_n11928), 
	.CK(HCLK__L5_N2));
   DFFR_X1 Q4h3z4_reg (.RN(FE_OFN34_HRESETn), 
	.QN(n5619), 
	.D(FE_PHN1664_n13747), 
	.CK(HCLK__L5_N27));
   DFFR_X1 Ark2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16834), 
	.Q(n16835), 
	.D(FE_PHN1613_n5777), 
	.CK(HCLK__L5_N9));
   DFFR_X1 U7w2z4_reg (.RN(FE_OFN152_HRESETn), 
	.QN(n5229), 
	.Q(n3066), 
	.D(FE_PHN4316_n5799), 
	.CK(hclk));
   DFFR_X1 Ffj2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16861), 
	.Q(n16863), 
	.D(FE_PHN1428_n5789), 
	.CK(HCLK__L5_N9));
   DFFR_X1 Sgj2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16857), 
	.Q(n16694), 
	.D(n5774), 
	.CK(HCLK__L5_N9));
   DFFR_X1 C3w2z4_reg (.RN(FE_OFN192_HRESETn), 
	.QN(n5227), 
	.Q(n3222), 
	.D(FE_PHN1653_U802_Z_0), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Vaw2z4_reg (.RN(FE_OFN175_HRESETn), 
	.QN(n5231), 
	.Q(n375), 
	.D(FE_PHN1903_n5795), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Wxp2z4_reg (.RN(FE_OFN192_HRESETn), 
	.QN(n5102), 
	.Q(n3223), 
	.D(FE_PHN1646_U518_Z_0), 
	.CK(HCLK__L5_N3));
   DFFR_X1 Gji2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n4956), 
	.Q(n1096), 
	.D(FE_PHN1426_U227_Z_0), 
	.CK(HCLK__L5_N4));
   DFFR_X1 L8t2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16822), 
	.Q(n16681), 
	.D(FE_PHN1157_n5823), 
	.CK(HCLK__L5_N4));
   DFFR_X1 Aii3z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n4834), 
	.D(FE_PHN1469_n4875), 
	.CK(HCLK__L5_N4));
   DFFR_X1 Jhy2z4_reg (.RN(FE_OFN175_HRESETn), 
	.Q(n1002), 
	.D(n5796), 
	.CK(HCLK__L5_N5));
   DFFR_X1 Kop2z4_reg (.RN(FE_OFN152_HRESETn), 
	.QN(n5096), 
	.Q(n3874), 
	.D(FE_PHN3497_n5792), 
	.CK(hclk));
   DFFR_X1 Mjl2z4_reg (.RN(FE_OFN56_HRESETn), 
	.QN(n5017), 
	.Q(n3875), 
	.D(FE_PHN3478_n5793), 
	.CK(hclk));
   DFFR_X1 Tki2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16872), 
	.Q(n16689), 
	.D(FE_PHN1431_n5775), 
	.CK(HCLK__L5_N4));
   DFFS_X1 O5t2z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n16806), 
	.Q(n16805), 
	.D(n5778), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Sjj2z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n4978), 
	.Q(n3488), 
	.D(FE_PHN1652_U134_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Fgm2z4_reg (.SN(FE_OFN144_HRESETn), 
	.QN(n5036), 
	.Q(n3480), 
	.D(FE_PHN1651_U121_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Cyq2z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n16810), 
	.Q(n16671), 
	.D(n5780), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Zcn2z4_reg (.SN(FE_OFN159_HRESETn), 
	.QN(n16809), 
	.Q(n16656), 
	.D(U756_Z_0), 
	.CK(HCLK__L5_N9));
   DFFS_X1 Yzi2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n4967), 
	.Q(n451), 
	.D(FE_PHN2948_n5752), 
	.CK(HCLK__L5_N3));
   DFFS_X1 Xly2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n5243), 
	.Q(n781), 
	.D(FE_PHN3056_n5748), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Lny2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n5244), 
	.Q(n659), 
	.D(FE_PHN2922_n5747), 
	.CK(HCLK__L5_N5));
   DFFS_X1 Bsy2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n16797), 
	.Q(n16686), 
	.D(FE_PHN3088_n5744), 
	.CK(HCLK__L5_N4));
   DFFS_X1 Pdi2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n4950), 
	.Q(n1697), 
	.D(n11746), 
	.CK(HCLK__L5_N9));
   DFFS_X2 Pty2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n16796), 
	.Q(n16657), 
	.D(FE_PHN2920_n5743), 
	.CK(HCLK__L5_N5));
   DFFS_X2 Qem2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n16807), 
	.Q(n16683), 
	.D(FE_PHN2954_n5753), 
	.CK(HCLK__L5_N5));
   DFFS_X2 U2x2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n16811), 
	.Q(n16659), 
	.D(FE_PHN3089_n5754), 
	.CK(HCLK__L5_N4));
   DFFS_X2 Zoy2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n16801), 
	.Q(n16674), 
	.D(FE_PHN729_n5746), 
	.CK(HCLK__L5_N5));
   DFFR_X2 K3l2z4_reg (.RN(FE_OFN55_HRESETn), 
	.QN(n5007), 
	.Q(n253), 
	.D(U792_Z_0), 
	.CK(HCLK__L5_N2));
   DFFS_X2 Jky2z4_reg (.SN(FE_OFN175_HRESETn), 
	.QN(n16794), 
	.Q(n16734), 
	.D(FE_PHN2921_n5749), 
	.CK(HCLK__L5_N3));
   DFFS_X2 Hyy2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n16795), 
	.Q(n16725), 
	.D(FE_PHN2952_n5740), 
	.CK(HCLK__L5_N4));
   DFFS_X2 Swy2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n16814), 
	.Q(n16733), 
	.D(FE_PHN2955_n5741), 
	.CK(HCLK__L5_N5));
   DFFR_X2 A4t2z4_reg (.RN(FE_OFN159_HRESETn), 
	.QN(n16680), 
	.Q(n16808), 
	.D(n5794), 
	.CK(HCLK__L5_N3));
   DFFS_X2 Nqy2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n16800), 
	.Q(n16798), 
	.D(FE_PHN2935_n5745), 
	.CK(HCLK__L5_N4));
   DFFR_X2 Emi2z4_reg (.RN(FE_OFN52_HRESETn), 
	.QN(n16865), 
	.Q(n16867), 
	.D(FE_PHN1508_n10553), 
	.CK(HCLK__L5_N9));
   DFFS_X2 H9i2z4_reg (.SN(FE_OFN52_HRESETn), 
	.QN(n16803), 
	.Q(n16802), 
	.D(FE_PHN2953_n5739), 
	.CK(HCLK__L5_N4));
   OR2_X4 U108 (.ZN(n16644), 
	.A2(n187), 
	.A1(n42));
   NOR2_X2 U112 (.ZN(n16645), 
	.A2(n16788), 
	.A1(n2998));
   NOR3_X2 U124 (.ZN(n16646), 
	.A3(n377), 
	.A2(n374), 
	.A1(n376));
   OR3_X4 U135 (.ZN(n16647), 
	.A3(n314), 
	.A2(n258), 
	.A1(n17108));
   AND2_X4 U137 (.ZN(n16648), 
	.A2(n4663), 
	.A1(n4665));
   AND2_X4 U141 (.ZN(n16649), 
	.A2(n4659), 
	.A1(n4661));
   AND2_X4 U144 (.ZN(n16650), 
	.A2(n4661), 
	.A1(n4665));
   AND3_X4 U145 (.ZN(n16651), 
	.A3(n4968), 
	.A2(n4662), 
	.A1(n4660));
   AND2_X4 U159 (.ZN(n16652), 
	.A2(n4658), 
	.A1(n4660));
   XOR2_X2 U190 (.Z(n16653), 
	.B(n16714), 
	.A(add_2073_A_13_));
   AND2_X4 U191 (.ZN(n16654), 
	.A2(n16661), 
	.A1(add_2073_A_30_));
   NAND2_X2 U197 (.ZN(n2169), 
	.A2(n4676), 
	.A1(FE_OFN10_n1697));
   XOR2_X2 U200 (.Z(n16655), 
	.B(n16665), 
	.A(add_2073_A_26_));
   XOR2_X2 U213 (.Z(n16658), 
	.B(n16707), 
	.A(add_2073_A_15_));
   OAI22_X2 U224 (.ZN(n247), 
	.B2(n2254), 
	.B1(n4239), 
	.A2(n2196), 
	.A1(n4401));
   AND2_X4 U227 (.ZN(n16660), 
	.A2(n16654), 
	.A1(add_2073_A_31_));
   AND2_X4 U236 (.ZN(n16661), 
	.A2(n16692), 
	.A1(add_2073_A_29_));
   AND2_X4 U239 (.ZN(n16662), 
	.A2(n16697), 
	.A1(add_2073_A_27_));
   XOR2_X2 U242 (.Z(n16663), 
	.B(n16697), 
	.A(add_2073_A_27_));
   AND2_X4 U250 (.ZN(n16664), 
	.A2(n16700), 
	.A1(add_2073_A_23_));
   AND2_X4 U251 (.ZN(n16665), 
	.A2(n16696), 
	.A1(add_2073_A_25_));
   AND2_X4 U253 (.ZN(n16666), 
	.A2(n16708), 
	.A1(add_2073_A_17_));
   AND2_X4 U254 (.ZN(n16667), 
	.A2(n16704), 
	.A1(add_2073_A_20_));
   XOR2_X2 U260 (.Z(n16668), 
	.B(n16699), 
	.A(add_2073_A_22_));
   AND2_X4 U267 (.ZN(n16669), 
	.A2(n16707), 
	.A1(add_2073_A_15_));
   AND2_X4 U270 (.ZN(n16670), 
	.A2(n16714), 
	.A1(add_2073_A_13_));
   XOR2_X2 U273 (.Z(n16672), 
	.B(n16703), 
	.A(add_2073_A_19_));
   AND2_X4 U276 (.ZN(n16673), 
	.A2(n16718), 
	.A1(add_2073_A_9_));
   XOR2_X2 U279 (.Z(n16675), 
	.B(add_2082_A_1_), 
	.A(add_2082_B_1_));
   AND2_X4 U282 (.ZN(n16676), 
	.A2(n16717), 
	.A1(add_2073_A_5_));
   AND2_X4 U285 (.ZN(n16677), 
	.A2(n16676), 
	.A1(add_2073_A_6_));
   AND2_X4 U288 (.ZN(n16678), 
	.A2(n16721), 
	.A1(add_2073_A_3_));
   XOR2_X2 U291 (.Z(n16679), 
	.B(n16670), 
	.A(add_2073_A_14_));
   XOR2_X2 U294 (.Z(n16682), 
	.B(n16678), 
	.A(add_2073_A_4_));
   XOR2_X2 U297 (.Z(n16684), 
	.B(n4168), 
	.A(n4068));
   OR3_X4 U300 (.ZN(n16685), 
	.A3(n261), 
	.A2(n4905), 
	.A1(n2926));
   XOR2_X2 U303 (.Z(n16688), 
	.B(n16660), 
	.A(add_2073_A_32_));
   AND2_X2 U306 (.ZN(n16691), 
	.A2(add_2082_A_1_), 
	.A1(add_2082_B_1_));
   AND2_X4 U309 (.ZN(n16692), 
	.A2(n16662), 
	.A1(add_2073_A_28_));
   XOR2_X1 U312 (.Z(n16693), 
	.B(n16661), 
	.A(add_2073_A_30_));
   XOR2_X2 U313 (.Z(n16695), 
	.B(n16692), 
	.A(add_2073_A_29_));
   AND2_X4 U315 (.ZN(n16696), 
	.A2(n16664), 
	.A1(add_2073_A_24_));
   AND2_X4 U316 (.ZN(n16697), 
	.A2(n16665), 
	.A1(add_2073_A_26_));
   XOR2_X2 U319 (.Z(n16698), 
	.B(n16662), 
	.A(add_2073_A_28_));
   AND2_X4 U353 (.ZN(n16699), 
	.A2(n16667), 
	.A1(add_2073_A_21_));
   AND2_X4 U359 (.ZN(n16700), 
	.A2(n16699), 
	.A1(add_2073_A_22_));
   XOR2_X2 U468 (.Z(n16701), 
	.B(n16696), 
	.A(add_2073_A_25_));
   XOR2_X2 U512 (.Z(n16702), 
	.B(n16700), 
	.A(add_2073_A_23_));
   AND2_X4 U582 (.ZN(n16703), 
	.A2(n16666), 
	.A1(add_2073_A_18_));
   AND2_X4 U648 (.ZN(n16704), 
	.A2(n16703), 
	.A1(add_2073_A_19_));
   XOR2_X2 U711 (.Z(n16705), 
	.B(n16664), 
	.A(add_2073_A_24_));
   XOR2_X2 U742 (.Z(n16706), 
	.B(n16667), 
	.A(add_2073_A_21_));
   AND2_X4 U751 (.ZN(n16707), 
	.A2(n16670), 
	.A1(add_2073_A_14_));
   AND2_X4 U752 (.ZN(n16708), 
	.A2(n16669), 
	.A1(add_2073_A_16_));
   XOR2_X2 U753 (.Z(n16709), 
	.B(n16704), 
	.A(add_2073_A_20_));
   XOR2_X2 U754 (.Z(n16710), 
	.B(n16666), 
	.A(add_2073_A_18_));
   XOR2_X2 U756 (.Z(n16711), 
	.B(n16708), 
	.A(add_2073_A_17_));
   AND2_X4 U757 (.ZN(n16712), 
	.A2(n16673), 
	.A1(add_2073_A_10_));
   AND2_X4 U758 (.ZN(n16713), 
	.A2(n16712), 
	.A1(add_2073_A_11_));
   AND2_X4 U759 (.ZN(n16714), 
	.A2(n16713), 
	.A1(add_2073_A_12_));
   XOR2_X2 U785 (.Z(n16715), 
	.B(n16669), 
	.A(add_2073_A_16_));
   AND2_X4 U812 (.ZN(n16716), 
	.A2(n16677), 
	.A1(add_2073_A_7_));
   AND2_X4 U820 (.ZN(n16717), 
	.A2(n16678), 
	.A1(add_2073_A_4_));
   AND2_X4 U837 (.ZN(n16718), 
	.A2(n16716), 
	.A1(add_2073_A_8_));
   XOR2_X2 U840 (.Z(n16719), 
	.B(n16713), 
	.A(add_2073_A_12_));
   AND2_X4 U841 (.ZN(n16720), 
	.A2(n16675), 
	.A1(add_2073_B_1_));
   AND2_X4 U845 (.ZN(n16721), 
	.A2(n16720), 
	.A1(add_2073_A_2_));
   XOR2_X2 U850 (.Z(n16722), 
	.B(n16718), 
	.A(add_2073_A_9_));
   XOR2_X2 U851 (.Z(n16723), 
	.B(n16712), 
	.A(add_2073_A_11_));
   OR2_X4 U852 (.ZN(haddr_o[15]), 
	.A2(n16737), 
	.A1(n16736));
   NAND3_X2 U856 (.ZN(n381), 
	.A3(n400), 
	.A2(n379), 
	.A1(n373));
   XOR2_X2 U857 (.Z(n16726), 
	.B(n16716), 
	.A(add_2073_A_8_));
   XOR2_X2 U858 (.Z(n16727), 
	.B(n16673), 
	.A(add_2073_A_10_));
   NOR2_X2 U879 (.ZN(n3118), 
	.A2(n4130), 
	.A1(n4131));
   XOR2_X2 U880 (.Z(n16729), 
	.B(n16721), 
	.A(add_2073_A_3_));
   XOR2_X2 U996 (.Z(n16730), 
	.B(n16717), 
	.A(add_2073_A_5_));
   XOR2_X2 U997 (.Z(n16731), 
	.B(n16676), 
	.A(add_2073_A_6_));
   NOR2_X2 U1000 (.ZN(n3275), 
	.A2(n4131), 
	.A1(n4142));
   XOR2_X2 U1006 (.Z(n16732), 
	.B(n16720), 
	.A(add_2073_A_2_));
   NAND4_X2 U1013 (.ZN(n979), 
	.A4(n2677), 
	.A3(n2676), 
	.A2(n2675), 
	.A1(n2674));
   OAI22_X2 U1022 (.ZN(n245), 
	.B2(n2253), 
	.B1(n4239), 
	.A2(n2250), 
	.A1(n4401));
   NAND2_X1 U1024 (.ZN(n16735), 
	.A2(n422), 
	.A1(n5649));
   OAI21_X2 U1027 (.ZN(n1632), 
	.B2(n2644), 
	.B1(n2643), 
	.A(n979));
   OAI221_X2 U1031 (.ZN(n2644), 
	.C2(FE_OFN103_n715), 
	.C1(n16862), 
	.B2(FE_OFN100_n1086), 
	.B1(n16845), 
	.A(n2645));
   NOR2_X1 U1051 (.ZN(n16736), 
	.A2(n1622), 
	.A1(n1661));
   INV_X1 U1054 (.ZN(n16737), 
	.A(n1662));
   OAI21_X2 U1112 (.ZN(n1622), 
	.B2(n2627), 
	.B1(n2626), 
	.A(n979));
   INV_X4 U1259 (.ZN(haddr_o[2]), 
	.A(n876));
   AOI221_X2 U1260 (.ZN(n876), 
	.C2(n1628), 
	.C1(n1640), 
	.B2(n17088), 
	.B1(n16729), 
	.A(n1641));
   OAI221_X2 U1264 (.ZN(haddr_o[19]), 
	.C2(n1632), 
	.C1(n1655), 
	.B2(n1622), 
	.B1(n1654), 
	.A(n1656));
   NAND4_X2 U1265 (.ZN(n1612), 
	.A4(n4590), 
	.A3(n4589), 
	.A2(n4588), 
	.A1(n1603));
   XOR2_X2 U1266 (.Z(n5818), 
	.B(n3407), 
	.A(n16990));
   NOR2_X2 U1267 (.ZN(n4240), 
	.A2(n5167), 
	.A1(n1614));
   INV_X4 U1270 (.ZN(haddr_o[5]), 
	.A(n968));
   AOI221_X2 U1271 (.ZN(n968), 
	.C2(n17088), 
	.C1(n16731), 
	.B2(n1628), 
	.B1(n1634), 
	.A(n1635));
   OAI21_X2 U1273 (.ZN(haddr_o[11]), 
	.B2(n1622), 
	.B1(n1695), 
	.A(n1731));
   XOR2_X2 U1275 (.Z(n5815), 
	.B(n2730), 
	.A(n16990));
   INV_X4 U1278 (.ZN(hwdata_o[31]), 
	.A(n4260));
   INV_X4 U1280 (.ZN(hwdata_o[26]), 
	.A(n24));
   INV_X4 U1281 (.ZN(haddr_o[4]), 
	.A(n967));
   AOI221_X2 U1283 (.ZN(n967), 
	.C2(n17088), 
	.C1(n16730), 
	.B2(n1628), 
	.B1(n1636), 
	.A(n1637));
   OAI22_X2 U1284 (.ZN(htrans_o[1]), 
	.B2(n999), 
	.B1(n1609), 
	.A2(n1608), 
	.A1(n1607));
   NOR3_X2 U1286 (.ZN(hsize_o[0]), 
	.A3(n1613), 
	.A2(n17090), 
	.A1(n1614));
   OAI221_X2 U1288 (.ZN(haddr_o[6]), 
	.C2(FE_OFN493_n1632), 
	.C1(n16782), 
	.B2(FE_OFN490_n1622), 
	.B1(n1630), 
	.A(n1633));
   XOR2_X2 U1289 (.Z(n5807), 
	.B(n3035), 
	.A(n2169));
   INV_X4 U1294 (.ZN(haddr_o[26]), 
	.A(n1149));
   AOI221_X2 U1296 (.ZN(n1149), 
	.C2(n17088), 
	.C1(n16663), 
	.B2(n1628), 
	.B1(n1645), 
	.A(n1646));
   INV_X4 U1297 (.ZN(haddr_o[17]), 
	.A(n1158));
   AOI221_X2 U1299 (.ZN(n1158), 
	.C2(n17088), 
	.C1(n16710), 
	.B2(n1628), 
	.B1(n1658), 
	.A(n1659));
   INV_X4 U1301 (.ZN(hwdata_o[27]), 
	.A(n208));
   INV_X4 U1303 (.ZN(haddr_o[20]), 
	.A(n1155));
   OAI21_X2 U1305 (.ZN(n2004), 
	.B2(n3213), 
	.B1(n3218), 
	.A(n2756));
   INV_X4 U1307 (.ZN(hwdata_o[29]), 
	.A(n4272));
   INV_X4 U1308 (.ZN(haddr_o[10]), 
	.A(n948));
   AOI221_X2 U1310 (.ZN(n948), 
	.C2(n17088), 
	.C1(n16723), 
	.B2(n1628), 
	.B1(n1667), 
	.A(n1668));
   NAND2_X2 U1312 (.ZN(FE_OFN113_HADDR_29_), 
	.A2(n1869), 
	.A1(n1620));
   OAI21_X2 U1313 (.ZN(haddr_o[9]), 
	.B2(n1622), 
	.B1(n1621), 
	.A(n1623));
   OAI22_X2 U1315 (.ZN(U186_Z_0), 
	.B2(n3534), 
	.B1(n2462), 
	.A2(n4610), 
	.A1(n2461));
   XOR2_X2 U1317 (.Z(n5819), 
	.B(n3356), 
	.A(n16990));
   INV_X4 U1318 (.ZN(hwdata_o[21]), 
	.A(n1116));
   AOI22_X2 U1320 (.ZN(n1116), 
	.B2(n4203), 
	.B1(n21), 
	.A2(n2556), 
	.A1(n4202));
   INV_X4 U1322 (.ZN(haddr_o[27]), 
	.A(n1148));
   INV_X4 U1324 (.ZN(haddr_o[18]), 
	.A(n1157));
   INV_X4 U1326 (.ZN(hwdata_o[28]), 
	.A(n205));
   INV_X4 U1328 (.ZN(hwdata_o[17]), 
	.A(n1112));
   AOI22_X2 U1329 (.ZN(n1112), 
	.B2(n4203), 
	.B1(n2258), 
	.A2(FE_OFN510_n2028), 
	.A1(n4202));
   INV_X4 U1331 (.ZN(hwdata_o[24]), 
	.A(n25));
   INV_X4 U1332 (.ZN(haddr_o[21]), 
	.A(n1154));
   AOI221_X2 U1334 (.ZN(n1154), 
	.C2(n17088), 
	.C1(n16668), 
	.B2(n1628), 
	.B1(n1651), 
	.A(n1652));
   OAI21_X2 U1367 (.ZN(n866), 
	.B2(n1169), 
	.B1(n1168), 
	.A(n17122));
   OAI211_X2 U1396 (.ZN(n1169), 
	.C2(n912), 
	.C1(FE_OFN425_n650), 
	.B(n1171), 
	.A(n1170));
   NAND4_X2 U1402 (.ZN(hwrite_o), 
	.A4(n1878), 
	.A3(n1877), 
	.A2(n1876), 
	.A1(n1875));
   OAI21_X2 U1465 (.ZN(n2871), 
	.B2(n3213), 
	.B1(n3427), 
	.A(n2756));
   NOR3_X2 U1466 (.ZN(haddr_o[1]), 
	.A3(n1613), 
	.A2(n683), 
	.A1(n1612));
   AOI222_X1 U1500 (.ZN(n683), 
	.C2(n1628), 
	.C1(n2232), 
	.B2(n17088), 
	.B1(n16732), 
	.A2(n2625), 
	.A1(n17090));
   OAI211_X2 U1501 (.ZN(n2011), 
	.C2(n3243), 
	.C1(n3242), 
	.B(n3245), 
	.A(n3244));
   INV_X4 U1509 (.ZN(hwdata_o[30]), 
	.A(n1077));
   AOI222_X1 U1512 (.ZN(n1077), 
	.C2(n4203), 
	.C1(n2083), 
	.B2(n4240), 
	.B1(n2253), 
	.A2(n4239), 
	.A1(n2250));
   OAI21_X2 U1519 (.ZN(hprot_o[3]), 
	.B2(n1617), 
	.B1(n1616), 
	.A(hprot_o[2]));
   OAI21_X2 U1521 (.ZN(haddr_o[3]), 
	.B2(FE_OFN490_n1622), 
	.B1(n1638), 
	.A(n1639));
   NOR2_X2 U1524 (.ZN(n2895), 
	.A2(n2926), 
	.A1(n3962));
   NAND2_X2 U1529 (.ZN(n2926), 
	.A2(n4172), 
	.A1(n1759));
   INV_X4 U1531 (.ZN(hwdata_o[23]), 
	.A(n4261));
   AOI22_X2 U1533 (.ZN(n4261), 
	.B2(FE_OFN516_n2196), 
	.B1(n4202), 
	.A2(n4203), 
	.A1(n3450));
   INV_X4 U1546 (.ZN(hwdata_o[18]), 
	.A(n1115));
   AOI22_X2 U1551 (.ZN(n1115), 
	.B2(n4203), 
	.B1(n2249), 
	.A2(n3177), 
	.A1(n4202));
   INV_X4 U1561 (.ZN(hsize_o[1]), 
	.A(n955));
   AOI21_X2 U1571 (.ZN(n955), 
	.B2(n979), 
	.B1(n1612), 
	.A(n1613));
   INV_X4 U1581 (.ZN(hwdata_o[20]), 
	.A(n1117));
   AOI22_X2 U1598 (.ZN(n1117), 
	.B2(n4203), 
	.B1(n20), 
	.A2(n2578), 
	.A1(n4202));
   INV_X4 U1604 (.ZN(hwdata_o[16]), 
	.A(n1118));
   AOI22_X2 U1607 (.ZN(n1118), 
	.B2(n4203), 
	.B1(n17), 
	.A2(n1354), 
	.A1(n4202));
   INV_X4 U1761 (.ZN(haddr_o[23]), 
	.A(n973));
   INV_X4 U1767 (.ZN(haddr_o[12]), 
	.A(n952));
   AOI221_X2 U1775 (.ZN(n952), 
	.C2(n17088), 
	.C1(n16653), 
	.B2(n1628), 
	.B1(n1665), 
	.A(n1666));
   INV_X4 U1776 (.ZN(haddr_o[24]), 
	.A(n317));
   INV_X4 U1807 (.ZN(haddr_o[14]), 
	.A(n956));
   INV_X4 U1813 (.ZN(haddr_o[13]), 
	.A(n957));
   INV_X4 U1818 (.ZN(hwdata_o[12]), 
	.A(n240));
   AOI22_X2 U1835 (.ZN(n240), 
	.B2(n2247), 
	.B1(n4401), 
	.A2(n4239), 
	.A1(n2578));
   INV_X4 U1900 (.ZN(lockup_o), 
	.A(n185));
   NOR2_X2 U1948 (.ZN(n185), 
	.A2(n1862), 
	.A1(n1861));
   INV_X4 U1950 (.ZN(hwdata_o[19]), 
	.A(n1114));
   AOI22_X2 U1951 (.ZN(n1114), 
	.B2(n4203), 
	.B1(n22), 
	.A2(n2257), 
	.A1(n4202));
   INV_X4 U1953 (.ZN(haddr_o[25]), 
	.A(n1150));
   INV_X4 U1962 (.ZN(haddr_o[16]), 
	.A(n1159));
   INV_X4 U1964 (.ZN(hwdata_o[25]), 
	.A(n201));
   INV_X4 U1965 (.ZN(haddr_o[22]), 
	.A(n1153));
   OR2_X4 U1967 (.ZN(hprot_o[2]), 
	.A2(haddr_o[30]), 
	.A1(SPCPT1_HADDR_29_));
   OAI221_X2 U2016 (.ZN(FE_OFN110_HADDR_30_), 
	.C2(n1632), 
	.C1(n16783), 
	.B2(n1622), 
	.B1(n1677), 
	.A(n1874));
   AOI22_X2 U2019 (.ZN(n4952), 
	.B2(n2463), 
	.B1(n2462), 
	.A2(n2461), 
	.A1(n2260));
   NOR2_X2 U2026 (.ZN(sleeping_o), 
	.A2(n16821), 
	.A1(n4834));
   INV_X4 U2028 (.ZN(hwdata_o[4]), 
	.A(n221));
   NAND2_X2 U2029 (.ZN(n221), 
	.A2(FE_OFN19_n1063), 
	.A1(n2578));
   OAI221_X2 U2031 (.ZN(n2909), 
	.C2(n3762), 
	.C1(n3761), 
	.B2(n3760), 
	.B1(n3754), 
	.A(n3763));
   INV_X4 U2033 (.ZN(hwdata_o[7]), 
	.A(n229));
   INV_X4 U2034 (.ZN(hwdata_o[5]), 
	.A(n224));
   NAND2_X2 U2056 (.ZN(n224), 
	.A2(FE_OFN19_n1063), 
	.A1(n2556));
   INV_X4 U2066 (.ZN(hwdata_o[3]), 
	.A(n218));
   NAND2_X2 U2068 (.ZN(n218), 
	.A2(FE_OFN19_n1063), 
	.A1(n2257));
   INV_X4 U2069 (.ZN(hwdata_o[6]), 
	.A(n226));
   INV_X4 U2071 (.ZN(hwdata_o[1]), 
	.A(n210));
   NAND2_X2 U2073 (.ZN(n210), 
	.A2(FE_OFN19_n1063), 
	.A1(n2028));
   INV_X4 U2091 (.ZN(hwdata_o[0]), 
	.A(n249));
   NAND2_X2 U2099 (.ZN(n249), 
	.A2(FE_OFN19_n1063), 
	.A1(n1354));
   INV_X4 U2101 (.ZN(haddr_o[28]), 
	.A(n878));
   AOI221_X2 U2102 (.ZN(n878), 
	.C2(n17088), 
	.C1(n16695), 
	.B2(n1628), 
	.B1(n1832), 
	.A(n1833));
   INV_X4 U2104 (.ZN(hwdata_o[10]), 
	.A(n236));
   AOI22_X2 U2106 (.ZN(n236), 
	.B2(n3145), 
	.B1(n4401), 
	.A2(n4239), 
	.A1(n3177));
   INV_X4 U2107 (.ZN(hwdata_o[13]), 
	.A(n242));
   AOI22_X2 U2128 (.ZN(n242), 
	.B2(n2259), 
	.B1(n4401), 
	.A2(n4239), 
	.A1(FE_OFN541_n2556));
   INV_X4 U2137 (.ZN(hwdata_o[8]), 
	.A(n232));
   AOI22_X2 U2139 (.ZN(n232), 
	.B2(n2261), 
	.B1(FE_OFN568_n4401), 
	.A2(n4239), 
	.A1(FE_OFN484_n1354));
   OAI211_X2 U2140 (.ZN(n2008), 
	.C2(n3217), 
	.C1(n3215), 
	.B(n3285), 
	.A(n3284));
   NAND2_X2 U2142 (.ZN(n3217), 
	.A2(n3867), 
	.A1(n1777));
   NOR4_X2 U2144 (.ZN(haddr_o[0]), 
	.A4(n1612), 
	.A3(n1613), 
	.A2(n1670), 
	.A1(n1669));
   NAND4_X2 U2165 (.ZN(hprot_o[0]), 
	.A4(n2686), 
	.A3(n2685), 
	.A2(n2674), 
	.A1(n1876));
   INV_X4 U2174 (.ZN(hwdata_o[2]), 
	.A(n215));
   NAND2_X2 U2176 (.ZN(n215), 
	.A2(FE_OFN19_n1063), 
	.A1(n3177));
   INV_X4 U2177 (.ZN(hwdata_o[15]), 
	.A(n247));
   INV_X4 U2179 (.ZN(hwdata_o[14]), 
	.A(n245));
   OR4_X4 U2181 (.ZN(n969), 
	.A4(haddr_o[9]), 
	.A3(haddr_o[7]), 
	.A2(n963), 
	.A1(n948));
   INV_X4 U2203 (.ZN(haddr_o[7]), 
	.A(n1147));
   INV_X4 U2219 (.ZN(hwdata_o[11]), 
	.A(n238));
   AOI22_X2 U2240 (.ZN(n238), 
	.B2(n2246), 
	.B1(n4401), 
	.A2(n4239), 
	.A1(FE_OFN519_n2257));
   INV_X4 U2274 (.ZN(hwdata_o[9]), 
	.A(n234));
   AOI22_X2 U2309 (.ZN(n234), 
	.B2(n4239), 
	.B1(n2028), 
	.A2(n3287), 
	.A1(n4401));
   INV_X4 U2331 (.ZN(hwdata_o[22]), 
	.A(n19));
   OAI22_X2 U2332 (.ZN(n19), 
	.B2(n2251), 
	.B1(n4202), 
	.A2(n2250), 
	.A1(n4203));
   NOR3_X2 U2333 (.ZN(txev_o), 
	.A3(n1784), 
	.A2(n16824), 
	.A1(n1088));
   AOI211_X2 U2341 (.ZN(n2076), 
	.C2(n3213), 
	.C1(n2376), 
	.B(n3425), 
	.A(n3609));
   INV_X4 U2344 (.ZN(n3425), 
	.A(n3209));
   OAI21_X2 U2345 (.ZN(FE_OFN117_HADDR_31_), 
	.B2(n979), 
	.B1(n1618), 
	.A(n1871));
   OAI21_X2 U2346 (.ZN(haddr_o[8]), 
	.B2(n1622), 
	.B1(n1625), 
	.A(n1626));
   INV_X4 U2347 (.ZN(n16792), 
	.A(n16738));
   INV_X4 U2379 (.ZN(n17103), 
	.A(n17104));
   INV_X4 U2385 (.ZN(n17074), 
	.A(n17077));
   INV_X4 U2402 (.ZN(n17053), 
	.A(n17057));
   INV_X4 U2443 (.ZN(n17018), 
	.A(n17022));
   INV_X4 U2454 (.ZN(n17048), 
	.A(n17052));
   INV_X4 U2457 (.ZN(n17068), 
	.A(n17071));
   INV_X4 U2486 (.ZN(n17038), 
	.A(n17042));
   INV_X4 U2493 (.ZN(n17023), 
	.A(n17027));
   INV_X4 U2537 (.ZN(n17116), 
	.A(n16644));
   INV_X4 U2556 (.ZN(n17117), 
	.A(n36));
   INV_X4 U2569 (.ZN(n597), 
	.A(n532));
   INV_X4 U2571 (.ZN(n16956), 
	.A(n16957));
   INV_X4 U2593 (.ZN(n2337), 
	.A(n16788));
   INV_X4 U2605 (.ZN(n17088), 
	.A(n1632));
   INV_X4 U2607 (.ZN(n17090), 
	.A(n979));
   AND2_X2 U2641 (.ZN(n16738), 
	.A2(n527), 
	.A1(n17102));
   INV_X4 U2643 (.ZN(n17102), 
	.A(n866));
   INV_X4 U2644 (.ZN(n17104), 
	.A(n318));
   NAND2_X2 U2646 (.ZN(n699), 
	.A2(n17096), 
	.A1(n195));
   INV_X4 U2648 (.ZN(n17077), 
	.A(n16742));
   INV_X4 U2668 (.ZN(n17057), 
	.A(n16740));
   INV_X4 U2682 (.ZN(n17022), 
	.A(n16741));
   INV_X4 U2684 (.ZN(n17052), 
	.A(n16743));
   INV_X4 U2685 (.ZN(n17027), 
	.A(n16744));
   INV_X4 U2687 (.ZN(n17042), 
	.A(n16745));
   INV_X4 U2715 (.ZN(n17071), 
	.A(n16739));
   INV_X4 U2763 (.ZN(n17092), 
	.A(n200));
   INV_X4 U2798 (.ZN(n17043), 
	.A(n17046));
   INV_X4 U2821 (.ZN(n17028), 
	.A(n17031));
   INV_X4 U2833 (.ZN(n29), 
	.A(n54));
   INV_X4 U2867 (.ZN(n17058), 
	.A(n17062));
   INV_X4 U2870 (.ZN(n17078), 
	.A(n17082));
   INV_X4 U2880 (.ZN(n17063), 
	.A(n17067));
   INV_X4 U2910 (.ZN(n17013), 
	.A(n17017));
   INV_X4 U2936 (.ZN(n17033), 
	.A(n17037));
   NAND2_X2 U2971 (.ZN(n443), 
	.A2(n466), 
	.A1(n473));
   NAND2_X2 U2991 (.ZN(n532), 
	.A2(FE_OFN90_n16849), 
	.A1(n16870));
   NAND2_X2 U3000 (.ZN(n653), 
	.A2(n16860), 
	.A1(n16825));
   INV_X4 U3002 (.ZN(n991), 
	.A(FE_OFN106_n585));
   INV_X4 U3003 (.ZN(n16957), 
	.A(n2222));
   INV_X4 U3005 (.ZN(n16979), 
	.A(n2637));
   INV_X2 U3007 (.ZN(n16971), 
	.A(FE_PSN5237_n2184));
   INV_X4 U3034 (.ZN(n527), 
	.A(n640));
   INV_X4 U3037 (.ZN(n17096), 
	.A(n17097));
   INV_X4 U3071 (.ZN(n16988), 
	.A(n3180));
   INV_X2 U3078 (.ZN(n16970), 
	.A(FE_PSN5237_n2184));
   NAND2_X2 U3088 (.ZN(n696), 
	.A2(FE_OFN17_n16805), 
	.A1(n16825));
   NAND2_X2 U3094 (.ZN(n745), 
	.A2(n17096), 
	.A1(n16859));
   INV_X4 U3098 (.ZN(n526), 
	.A(FE_OFN104_n715));
   INV_X4 U3112 (.ZN(n1574), 
	.A(n1086));
   INV_X4 U3127 (.ZN(n827), 
	.A(n673));
   INV_X4 U3130 (.ZN(n529), 
	.A(n1519));
   INV_X4 U3141 (.ZN(n565), 
	.A(n918));
   INV_X4 U3148 (.ZN(n17083), 
	.A(n1514));
   INV_X2 U3159 (.ZN(n16972), 
	.A(FE_PSN5237_n2184));
   INV_X1 U3160 (.ZN(n16955), 
	.A(n16957));
   INV_X4 U3162 (.ZN(n16990), 
	.A(n16991));
   INV_X4 U3164 (.ZN(n16895), 
	.A(n16652));
   NOR2_X2 U3175 (.ZN(n2391), 
	.A2(n2233), 
	.A1(n1754));
   INV_X4 U3188 (.ZN(n16954), 
	.A(n16957));
   INV_X2 U3220 (.ZN(n16980), 
	.A(n2637));
   INV_X4 U3224 (.ZN(n16882), 
	.A(n16648));
   INV_X4 U3241 (.ZN(n16910), 
	.A(n16911));
   INV_X4 U3248 (.ZN(n16875), 
	.A(n16649));
   INV_X4 U3264 (.ZN(n16873), 
	.A(n16650));
   INV_X4 U3267 (.ZN(n17098), 
	.A(n17099));
   INV_X4 U3275 (.ZN(n592), 
	.A(n851));
   INV_X4 U3338 (.ZN(n16788), 
	.A(n16684));
   INV_X4 U3342 (.ZN(n16992), 
	.A(n2127));
   INV_X4 U3350 (.ZN(n16942), 
	.A(n3279));
   INV_X4 U3351 (.ZN(n16951), 
	.A(n3118));
   INV_X4 U3355 (.ZN(n16948), 
	.A(n3275));
   INV_X4 U3356 (.ZN(n16945), 
	.A(n3277));
   INV_X4 U3384 (.ZN(n1628), 
	.A(n1622));
   NAND2_X2 U3396 (.ZN(n650), 
	.A2(n16870), 
	.A1(n897));
   INV_X4 U3397 (.ZN(n195), 
	.A(n499));
   INV_X4 U3399 (.ZN(n17008), 
	.A(n2243));
   INV_X4 U3403 (.ZN(n16994), 
	.A(n2501));
   AND2_X2 U3406 (.ZN(n16739), 
	.A2(n3446), 
	.A1(n3438));
   AND2_X2 U3410 (.ZN(n16740), 
	.A2(n3435), 
	.A1(n3445));
   AND2_X2 U3412 (.ZN(n16741), 
	.A2(n3435), 
	.A1(n3442));
   AND2_X2 U3413 (.ZN(n16742), 
	.A2(n3446), 
	.A1(n3435));
   AND2_X2 U3415 (.ZN(n16743), 
	.A2(n3438), 
	.A1(n3445));
   AND2_X2 U3416 (.ZN(n16744), 
	.A2(n3438), 
	.A1(n3442));
   AND2_X2 U3418 (.ZN(n16745), 
	.A2(n3438), 
	.A1(n3437));
   INV_X4 U3419 (.ZN(n3215), 
	.A(n3213));
   INV_X4 U3423 (.ZN(n17017), 
	.A(n16750));
   INV_X4 U3424 (.ZN(n17037), 
	.A(n16748));
   INV_X4 U3427 (.ZN(n17062), 
	.A(n16749));
   INV_X4 U3428 (.ZN(n17082), 
	.A(n16751));
   INV_X4 U3447 (.ZN(n17046), 
	.A(n16746));
   INV_X4 U3448 (.ZN(n17031), 
	.A(n16747));
   INV_X4 U3450 (.ZN(n17001), 
	.A(n17005));
   INV_X4 U3454 (.ZN(n17067), 
	.A(n16752));
   NAND2_X2 U3494 (.ZN(n585), 
	.A2(n16864), 
	.A1(FE_OFN78_n16834));
   INV_X1 U3562 (.ZN(n16964), 
	.A(n2182));
   INV_X4 U3566 (.ZN(n16984), 
	.A(n16754));
   INV_X4 U3568 (.ZN(n16963), 
	.A(n2191));
   INV_X4 U3574 (.ZN(n16966), 
	.A(n2182));
   INV_X4 U3577 (.ZN(n16969), 
	.A(n16753));
   INV_X4 U3580 (.ZN(n16960), 
	.A(n2190));
   INV_X4 U3581 (.ZN(n16864), 
	.A(n16865));
   INV_X4 U3583 (.ZN(n16837), 
	.A(FE_OFN85_n16839));
   INV_X4 U3637 (.ZN(n16825), 
	.A(n16826));
   INV_X4 U3641 (.ZN(n16860), 
	.A(n16861));
   INV_X4 U3642 (.ZN(n16870), 
	.A(n16871));
   INV_X4 U3645 (.ZN(n16849), 
	.A(n16850));
   INV_X4 U3646 (.ZN(n17097), 
	.A(n797));
   NAND2_X2 U3649 (.ZN(n715), 
	.A2(FE_OFN82_n16856), 
	.A1(n16851));
   NAND2_X2 U3650 (.ZN(n1086), 
	.A2(FE_OFN85_n16839), 
	.A1(FE_OFN87_n16848));
   NAND2_X2 U3651 (.ZN(n640), 
	.A2(n17096), 
	.A1(FE_OFN79_n16834));
   NAND2_X2 U3652 (.ZN(n617), 
	.A2(n16860), 
	.A1(n16845));
   NAND2_X2 U3655 (.ZN(n1104), 
	.A2(n16842), 
	.A1(FE_OFN81_n16856));
   INV_X4 U3656 (.ZN(n16976), 
	.A(n16755));
   INV_X4 U3659 (.ZN(n16939), 
	.A(n16759));
   INV_X4 U3660 (.ZN(n16916), 
	.A(n16760));
   INV_X4 U3663 (.ZN(n16933), 
	.A(n16756));
   INV_X2 U3665 (.ZN(n16982), 
	.A(n16754));
   INV_X4 U3666 (.ZN(n16877), 
	.A(n16763));
   INV_X2 U3669 (.ZN(n16967), 
	.A(n16753));
   INV_X2 U3671 (.ZN(n16968), 
	.A(n16753));
   INV_X2 U3673 (.ZN(n16958), 
	.A(n2190));
   INV_X2 U3674 (.ZN(n16959), 
	.A(n2190));
   INV_X4 U3675 (.ZN(n16913), 
	.A(n16762));
   INV_X2 U3695 (.ZN(n16962), 
	.A(n2191));
   INV_X2 U3696 (.ZN(n16965), 
	.A(n2182));
   INV_X4 U3705 (.ZN(n16905), 
	.A(n16757));
   INV_X4 U3721 (.ZN(n16908), 
	.A(n16761));
   INV_X4 U3729 (.ZN(n16885), 
	.A(n16758));
   INV_X1 U3732 (.ZN(n16848), 
	.A(n16850));
   INV_X4 U3733 (.ZN(n16842), 
	.A(n16844));
   INV_X4 U3737 (.ZN(n16828), 
	.A(n16833));
   INV_X4 U3741 (.ZN(n16836), 
	.A(n16728));
   INV_X4 U3746 (.ZN(n16831), 
	.A(n16833));
   INV_X4 U3749 (.ZN(n16843), 
	.A(n16844));
   NAND2_X2 U3750 (.ZN(n1519), 
	.A2(n16855), 
	.A1(FE_OFN70_n16867));
   NAND2_X2 U3755 (.ZN(n673), 
	.A2(n16862), 
	.A1(n16838));
   NAND2_X2 U3758 (.ZN(n918), 
	.A2(FE_OFN85_n16839), 
	.A1(n16855));
   INV_X4 U3759 (.ZN(n2198), 
	.A(n2543));
   INV_X4 U3765 (.ZN(n16911), 
	.A(n4211));
   INV_X1 U3768 (.ZN(n16977), 
	.A(n16755));
   INV_X4 U3769 (.ZN(n16991), 
	.A(n2169));
   INV_X4 U3776 (.ZN(n16934), 
	.A(n16756));
   INV_X4 U3777 (.ZN(n16886), 
	.A(n16767));
   INV_X4 U3782 (.ZN(n16897), 
	.A(n16764));
   INV_X2 U3785 (.ZN(n16961), 
	.A(n2191));
   INV_X4 U3786 (.ZN(n16891), 
	.A(n16766));
   INV_X4 U3791 (.ZN(n16902), 
	.A(n16765));
   INV_X4 U3794 (.ZN(n16859), 
	.A(n16861));
   INV_X4 U3825 (.ZN(n16824), 
	.A(n16690));
   INV_X4 U3842 (.ZN(n16854), 
	.A(n16694));
   INV_X2 U3865 (.ZN(n16847), 
	.A(n16850));
   INV_X4 U3937 (.ZN(n16868), 
	.A(n16689));
   INV_X4 U3938 (.ZN(n16855), 
	.A(n16694));
   INV_X4 U3940 (.ZN(n16838), 
	.A(n16728));
   NOR2_X2 U3943 (.ZN(n1808), 
	.A2(n2078), 
	.A1(n2077));
   NAND2_X2 U3945 (.ZN(n499), 
	.A2(n16862), 
	.A1(n16851));
   INV_X2 U3948 (.ZN(n16983), 
	.A(n16754));
   INV_X4 U3976 (.ZN(n16893), 
	.A(n16651));
   INV_X4 U4010 (.ZN(n17099), 
	.A(n16686));
   AOI211_X2 U4027 (.ZN(n2519), 
	.C2(n17008), 
	.C1(n2250), 
	.B(n2521), 
	.A(n2520));
   NAND2_X2 U4041 (.ZN(n851), 
	.A2(n16820), 
	.A1(FE_OFN75_n16806));
   INV_X4 U4047 (.ZN(n16820), 
	.A(n16681));
   NAND2_X2 U4055 (.ZN(n379), 
	.A2(n1340), 
	.A1(n400));
   INV_X4 U4059 (.ZN(n16812), 
	.A(n16813));
   INV_X4 U4064 (.ZN(n2131), 
	.A(n2126));
   INV_X4 U4067 (.ZN(n2882), 
	.A(n2926));
   INV_X4 U4068 (.ZN(n2055), 
	.A(n2124));
   INV_X4 U4073 (.ZN(n2878), 
	.A(n2981));
   INV_X4 U4076 (.ZN(n4203), 
	.A(n4202));
   INV_X4 U4077 (.ZN(n2922), 
	.A(n2998));
   AND2_X2 U4087 (.ZN(n16746), 
	.A2(n3443), 
	.A1(n3445));
   AND2_X2 U4090 (.ZN(n16747), 
	.A2(n3443), 
	.A1(n3442));
   OAI21_X2 U4091 (.ZN(n3213), 
	.B2(n4070), 
	.B1(n17096), 
	.A(n3546));
   NOR2_X2 U4094 (.ZN(n37), 
	.A2(n1007), 
	.A1(FE_PHN675_n17126));
   NAND4_X2 U4114 (.ZN(n200), 
	.A4(FE_OFN81_n16856), 
	.A3(n16820), 
	.A2(n760), 
	.A1(n809));
   NAND2_X2 U4115 (.ZN(n819), 
	.A2(n16725), 
	.A1(n791));
   AND2_X2 U4118 (.ZN(n16748), 
	.A2(n3439), 
	.A1(n3437));
   AND2_X2 U4119 (.ZN(n16749), 
	.A2(n3439), 
	.A1(n3445));
   AND2_X2 U4123 (.ZN(n16750), 
	.A2(n3439), 
	.A1(n3442));
   AND2_X2 U4124 (.ZN(n16751), 
	.A2(n3439), 
	.A1(n3446));
   INV_X4 U4127 (.ZN(n17005), 
	.A(n16768));
   INV_X4 U4133 (.ZN(n16996), 
	.A(n17000));
   INV_X4 U4137 (.ZN(n16816), 
	.A(n16687));
   AND2_X2 U4143 (.ZN(n16752), 
	.A2(n3446), 
	.A1(n3443));
   NOR2_X2 U4144 (.ZN(n1317), 
	.A2(n1124), 
	.A1(n1125));
   INV_X4 U4147 (.ZN(n17109), 
	.A(n16769));
   INV_X4 U4154 (.ZN(n17124), 
	.A(FE_PHN674_n17127));
   INV_X4 U4155 (.ZN(n17094), 
	.A(n17095));
   INV_X4 U4159 (.ZN(n17122), 
	.A(FE_PHN675_n17126));
   INV_X4 U4164 (.ZN(n17106), 
	.A(n16647));
   NAND2_X2 U4174 (.ZN(n1131), 
	.A2(n1109), 
	.A1(n373));
   NAND3_X2 U4175 (.ZN(n16753), 
	.A3(n3593), 
	.A2(n3436), 
	.A1(n3592));
   NAND2_X2 U4178 (.ZN(n16754), 
	.A2(n3480), 
	.A1(n3593));
   INV_X4 U4179 (.ZN(n16985), 
	.A(n16770));
   INV_X4 U4194 (.ZN(n16839), 
	.A(n16840));
   INV_X4 U4197 (.ZN(n16826), 
	.A(n16827));
   OR2_X1 U4198 (.ZN(n16755), 
	.A2(n3601), 
	.A1(n16956));
   AND2_X2 U4204 (.ZN(n16756), 
	.A2(n3492), 
	.A1(n4162));
   AND2_X2 U4210 (.ZN(n16757), 
	.A2(n4658), 
	.A1(n4657));
   AND2_X2 U4224 (.ZN(n16758), 
	.A2(n4657), 
	.A1(n4662));
   NAND2_X2 U4226 (.ZN(n16759), 
	.A2(n3480), 
	.A1(n4163));
   NAND2_X2 U4230 (.ZN(n16760), 
	.A2(n4659), 
	.A1(n4663));
   AND2_X2 U4231 (.ZN(n16761), 
	.A2(n4658), 
	.A1(n4659));
   NAND2_X2 U4236 (.ZN(n16762), 
	.A2(n4659), 
	.A1(n4662));
   NAND2_X2 U4241 (.ZN(n16763), 
	.A2(n4657), 
	.A1(n4661));
   INV_X4 U4243 (.ZN(n16851), 
	.A(n16852));
   INV_X4 U4249 (.ZN(n16833), 
	.A(n16835));
   INV_X2 U4260 (.ZN(n16856), 
	.A(n16857));
   INV_X2 U4263 (.ZN(n16986), 
	.A(n16770));
   INV_X4 U4264 (.ZN(n16987), 
	.A(n16770));
   INV_X4 U4268 (.ZN(n16845), 
	.A(n16846));
   INV_X4 U4271 (.ZN(n16871), 
	.A(n16872));
   INV_X4 U4272 (.ZN(n16821), 
	.A(n16822));
   INV_X2 U4277 (.ZN(n16973), 
	.A(n16773));
   INV_X4 U4280 (.ZN(n16930), 
	.A(n16772));
   INV_X4 U4281 (.ZN(n16918), 
	.A(n16771));
   INV_X4 U4286 (.ZN(n16936), 
	.A(n16775));
   INV_X4 U4289 (.ZN(n16927), 
	.A(n16774));
   INV_X4 U4290 (.ZN(n16975), 
	.A(n16773));
   NAND2_X2 U4291 (.ZN(n16764), 
	.A2(n4658), 
	.A1(n4665));
   NAND3_X2 U4297 (.ZN(n16765), 
	.A3(n4660), 
	.A2(n3436), 
	.A1(n4662));
   NAND2_X2 U4300 (.ZN(n16766), 
	.A2(n4662), 
	.A1(n4665));
   NAND2_X2 U4301 (.ZN(n16767), 
	.A2(n4663), 
	.A1(n4660));
   INV_X4 U4302 (.ZN(n16862), 
	.A(n16863));
   INV_X4 U4307 (.ZN(n16924), 
	.A(n16777));
   INV_X2 U4310 (.ZN(n16925), 
	.A(n16777));
   INV_X4 U4311 (.ZN(n16921), 
	.A(n16776));
   INV_X2 U4312 (.ZN(n16922), 
	.A(n16776));
   INV_X4 U4315 (.ZN(n16931), 
	.A(n16772));
   INV_X4 U4320 (.ZN(n16919), 
	.A(n16771));
   INV_X2 U4325 (.ZN(n16974), 
	.A(n16773));
   NOR2_X2 U4343 (.ZN(n1750), 
	.A2(n2001), 
	.A1(n179));
   INV_X4 U4344 (.ZN(n16817), 
	.A(n16818));
   NOR2_X2 U4345 (.ZN(n475), 
	.A2(n16659), 
	.A1(FE_OFN21_n503));
   NAND2_X2 U4347 (.ZN(n616), 
	.A2(n16820), 
	.A1(n16680));
   INV_X4 U4348 (.ZN(n16804), 
	.A(n16802));
   INV_X4 U4350 (.ZN(n16813), 
	.A(n16814));
   NAND2_X2 U4351 (.ZN(n1900), 
	.A2(n2172), 
	.A1(n2231));
   NAND2_X2 U4355 (.ZN(n2948), 
	.A2(n2882), 
	.A1(n252));
   NAND2_X2 U4362 (.ZN(n3011), 
	.A2(n2882), 
	.A1(n3873));
   INV_X4 U4365 (.ZN(n2879), 
	.A(n2918));
   NAND2_X2 U4366 (.ZN(n334), 
	.A2(n1002), 
	.A1(n336));
   NAND2_X2 U4367 (.ZN(n2998), 
	.A2(n4077), 
	.A1(n1759));
   NAND2_X2 U4369 (.ZN(n4202), 
	.A2(n1612), 
	.A1(FE_OFN19_n1063));
   NAND2_X2 U4370 (.ZN(n226), 
	.A2(FE_OFN19_n1063), 
	.A1(n2250));
   NAND2_X2 U4374 (.ZN(n229), 
	.A2(FE_OFN19_n1063), 
	.A1(FE_OFN516_n2196));
   INV_X4 U4379 (.ZN(n17120), 
	.A(n16779));
   INV_X4 U4395 (.ZN(n1124), 
	.A(n1385));
   NAND2_X2 U4402 (.ZN(n478), 
	.A2(n16807), 
	.A1(n822));
   AND3_X2 U4404 (.ZN(n16768), 
	.A3(n3437), 
	.A2(n3436), 
	.A1(n3435));
   INV_X4 U4406 (.ZN(n17000), 
	.A(n16780));
   NAND2_X2 U4418 (.ZN(n1892), 
	.A2(n253), 
	.A1(n1893));
   NAND2_X2 U4419 (.ZN(n1895), 
	.A2(n253), 
	.A1(n1897));
   AND3_X2 U4424 (.ZN(n16769), 
	.A3(n314), 
	.A2(n315), 
	.A1(n17107));
   INV_X4 U4425 (.ZN(n17095), 
	.A(n16781));
   INV_X4 U4435 (.ZN(n17126), 
	.A(hready_i));
   INV_X4 U4436 (.ZN(n16799), 
	.A(n16798));
   NAND2_X2 U4440 (.ZN(n213), 
	.A2(n253), 
	.A1(n252));
   NAND2_X2 U4441 (.ZN(n1889), 
	.A2(n253), 
	.A1(n1890));
   NAND2_X2 U4444 (.ZN(n1886), 
	.A2(n253), 
	.A1(n1887));
   INV_X4 U4445 (.ZN(n17107), 
	.A(n17108));
   INV_X4 U4448 (.ZN(n17127), 
	.A(hready_i));
   OR4_X4 U4570 (.ZN(n16770), 
	.A4(n4959), 
	.A3(n4978), 
	.A2(n5036), 
	.A1(n2184));
   NAND3_X2 U4571 (.ZN(n16771), 
	.A3(n5252), 
	.A2(n3592), 
	.A1(n4959));
   AND2_X4 U4574 (.ZN(n16772), 
	.A2(n5252), 
	.A1(n4162));
   NAND3_X1 U4575 (.ZN(n16773), 
	.A3(n3593), 
	.A2(n4968), 
	.A1(n3592));
   NAND3_X2 U4578 (.ZN(n16774), 
	.A3(n4959), 
	.A2(n3492), 
	.A1(n3592));
   NAND2_X2 U4579 (.ZN(n16775), 
	.A2(n5036), 
	.A1(n4163));
   OR4_X4 U4582 (.ZN(n16776), 
	.A4(FE_OFN583_n5036), 
	.A3(n5252), 
	.A2(n3495), 
	.A1(n3488));
   INV_X4 U4583 (.ZN(n16989), 
	.A(FE_OFN559_n3180));
   OR4_X1 U4584 (.ZN(n16777), 
	.A4(n5252), 
	.A3(n3480), 
	.A2(n3495), 
	.A1(n3488));
   OAI21_X2 U4588 (.ZN(n422), 
	.B2(n1066), 
	.B1(n1341), 
	.A(n183));
   NAND2_X2 U4592 (.ZN(n1821), 
	.A2(n2172), 
	.A1(n5027));
   NAND2_X2 U4593 (.ZN(n3566), 
	.A2(n5120), 
	.A1(n5027));
   NAND2_X2 U4597 (.ZN(n1820), 
	.A2(n2231), 
	.A1(n5120));
   NAND3_X2 U4600 (.ZN(n2918), 
	.A3(n1111), 
	.A2(FE_PHN1894_n5149), 
	.A1(n2882));
   INV_X4 U4601 (.ZN(n16787), 
	.A(n16685));
   OR2_X1 U4607 (.ZN(n266), 
	.A2(n16647), 
	.A1(n16778));
   XOR2_X2 U4608 (.Z(n16778), 
	.B(sub_2068_carry_23_), 
	.A(sub_2068_A_23_));
   NAND2_X2 U4609 (.ZN(n16779), 
	.A2(n180), 
	.A1(n37));
   AND3_X2 U4610 (.ZN(n16780), 
	.A3(n3437), 
	.A2(n4968), 
	.A1(n3435));
   INV_X4 U4622 (.ZN(n17108), 
	.A(n265));
   OR3_X1 U4638 (.ZN(n16781), 
	.A3(n261), 
	.A2(n4905), 
	.A1(FE_PHN1037_n5007));
   XNOR2_X2 U4696 (.ZN(n16782), 
	.B(n16677), 
	.A(add_2073_A_7_));
   INV_X4 U4697 (.ZN(add_2073_SUM_7_), 
	.A(n16782));
   XNOR2_X1 U4698 (.ZN(n16783), 
	.B(n16654), 
	.A(add_2073_A_31_));
   INV_X4 U4701 (.ZN(add_2073_SUM_31_), 
	.A(n16783));
   NAND2_X1 U4702 (.ZN(n16784), 
	.A2(n16660), 
	.A1(add_2073_A_32_));
   XNOR2_X2 U4703 (.ZN(U4_DATA1_0), 
	.B(n16784), 
	.A(add_2082_carry[33]));
   XNOR2_X2 U4706 (.ZN(n16785), 
	.B(n16675), 
	.A(add_2073_B_1_));
   INV_X4 U4708 (.ZN(add_2073_SUM_1_), 
	.A(n16785));
   INV_X4 U4711 (.ZN(n731), 
	.A(n1963));
   INV_X4 U4713 (.ZN(n708), 
	.A(n1228));
   INV_X4 U4715 (.ZN(n483), 
	.A(n945));
   INV_X4 U4720 (.ZN(n897), 
	.A(n1882));
   INV_X4 U4721 (.ZN(n473), 
	.A(n1198));
   INV_X4 U4725 (.ZN(n466), 
	.A(n579));
   NAND3_X2 U4726 (.ZN(n610), 
	.A3(n4708), 
	.A2(n4707), 
	.A1(n4706));
   INV_X4 U4727 (.ZN(n2732), 
	.A(n2719));
   NAND2_X2 U4728 (.ZN(n4427), 
	.A2(n4657), 
	.A1(n4663));
   INV_X4 U4732 (.ZN(n4192), 
	.A(n4335));
   INV_X4 U4733 (.ZN(n563), 
	.A(n1234));
   INV_X4 U4736 (.ZN(n1314), 
	.A(n1125));
   INV_X4 U4774 (.ZN(n2074), 
	.A(n2723));
   NAND2_X2 U4778 (.ZN(n2126), 
	.A2(n3550), 
	.A1(n3549));
   NAND4_X2 U4779 (.ZN(n2501), 
	.A4(FE_OFN10_n1697), 
	.A3(n16826), 
	.A2(FE_OFN70_n16867), 
	.A1(n3532));
   INV_X4 U4780 (.ZN(n543), 
	.A(n713));
   AND2_X4 U4782 (.ZN(n3434), 
	.A2(n2103), 
	.A1(FE_PHN703_n44));
   AND3_X4 U4783 (.ZN(n3402), 
	.A3(n3404), 
	.A2(n3403), 
	.A1(n48));
   AND3_X4 U4796 (.ZN(n3351), 
	.A3(n3353), 
	.A2(n3352), 
	.A1(n144));
   INV_X4 U4797 (.ZN(n2912), 
	.A(n2875));
   AND2_X4 U4804 (.ZN(n3286), 
	.A2(n2113), 
	.A1(n127));
   AND2_X4 U4805 (.ZN(n3171), 
	.A2(n2115), 
	.A1(FE_PHN2916_n171));
   AND2_X4 U4813 (.ZN(n3144), 
	.A2(n2114), 
	.A1(FE_PHN770_n140));
   NOR4_X2 U4821 (.ZN(n3097), 
	.A4(n3098), 
	.A3(n2310), 
	.A2(n2055), 
	.A1(n2309));
   AND3_X4 U4822 (.ZN(n3030), 
	.A3(n3032), 
	.A2(n3031), 
	.A1(n136));
   AND4_X4 U4830 (.ZN(n2973), 
	.A4(n2975), 
	.A3(n2974), 
	.A2(n2306), 
	.A1(n2124));
   AND4_X4 U4831 (.ZN(n2866), 
	.A4(n2867), 
	.A3(n2285), 
	.A2(n2305), 
	.A1(n2124));
   AND4_X4 U4835 (.ZN(n2843), 
	.A4(n2846), 
	.A3(n2845), 
	.A2(n2844), 
	.A1(n2696));
   AND3_X4 U4836 (.ZN(n2820), 
	.A3(n2822), 
	.A2(n2696), 
	.A1(n2821));
   AND4_X4 U4839 (.ZN(n2797), 
	.A4(n2799), 
	.A3(FE_OFN382_n64), 
	.A2(n2798), 
	.A1(n2696));
   AND3_X4 U4840 (.ZN(n2775), 
	.A3(n2777), 
	.A2(n2696), 
	.A1(n2776));
   AND4_X4 U4843 (.ZN(n2750), 
	.A4(n2753), 
	.A3(n2752), 
	.A2(n2751), 
	.A1(n2696));
   AND3_X4 U4844 (.ZN(n2725), 
	.A3(n2726), 
	.A2(n2696), 
	.A1(n58));
   AND4_X4 U4847 (.ZN(n2694), 
	.A4(n2697), 
	.A3(n2696), 
	.A2(n2695), 
	.A1(n61));
   AND3_X4 U4848 (.ZN(n2597), 
	.A3(n2598), 
	.A2(n2111), 
	.A1(FE_PHN693_n166));
   AND4_X4 U4851 (.ZN(n2573), 
	.A4(n2283), 
	.A3(n2262), 
	.A2(n2112), 
	.A1(FE_PHN778_n160));
   AND4_X4 U4852 (.ZN(n2549), 
	.A4(n2281), 
	.A3(n2263), 
	.A2(n2107), 
	.A1(FE_PHN783_n152));
   AND2_X4 U4853 (.ZN(n2494), 
	.A2(n2109), 
	.A1(n109));
   AND4_X4 U4855 (.ZN(n2470), 
	.A4(n2471), 
	.A3(n2234), 
	.A2(n2291), 
	.A1(n2124));
   AND3_X4 U4856 (.ZN(n2442), 
	.A3(n2444), 
	.A2(n2443), 
	.A1(FE_PHN735_n100));
   NOR3_X2 U4858 (.ZN(n2416), 
	.A3(n99), 
	.A2(n2055), 
	.A1(n2110));
   NOR3_X2 U4859 (.ZN(n2079), 
	.A3(n2081), 
	.A2(n2080), 
	.A1(n117));
   AND4_X4 U4860 (.ZN(n1807), 
	.A4(n2065), 
	.A3(n2064), 
	.A2(n2063), 
	.A1(n76));
   NOR3_X2 U4865 (.ZN(n1809), 
	.A3(n2056), 
	.A2(n2055), 
	.A1(n2054));
   AND3_X4 U4866 (.ZN(n1810), 
	.A3(n2014), 
	.A2(n2013), 
	.A1(n192));
   INV_X4 U4869 (.ZN(n1109), 
	.A(FE_PHN776_n1108));
   INV_X4 U4870 (.ZN(n336), 
	.A(n376));
   INV_X4 U4871 (.ZN(n338), 
	.A(n378));
   AND4_X4 U4878 (.ZN(n341), 
	.A4(n375), 
	.A3(n374), 
	.A2(n336), 
	.A1(n373));
   OR2_X4 U4882 (.ZN(n211), 
	.A2(n251), 
	.A1(n213));
   NOR2_X2 U4883 (.ZN(n54), 
	.A2(n188), 
	.A1(n42));
   AOI211_X2 U198 (.ZN(n13870), 
	.C2(n1426), 
	.C1(n4964), 
	.B(n1428), 
	.A(n1427));
   AOI211_X2 U211 (.ZN(n13795), 
	.C2(n1442), 
	.C1(n5126), 
	.B(FE_PHN2970_n1444), 
	.A(n1443));
   AOI211_X2 U222 (.ZN(n13813), 
	.C2(n1438), 
	.C1(n5582), 
	.B(n1440), 
	.A(n1439));
   AOI211_X2 U225 (.ZN(n13989), 
	.C2(n1381), 
	.C1(n5118), 
	.B(n1383), 
	.A(n1382));
   AOI211_X2 U234 (.ZN(n13835), 
	.C2(n1433), 
	.C1(n5061), 
	.B(n1435), 
	.A(n1434));
   AOI211_X2 U237 (.ZN(n13919), 
	.C2(n1405), 
	.C1(n5531), 
	.B(n1407), 
	.A(n1406));
   AOI211_X2 U240 (.ZN(n13932), 
	.C2(n1399), 
	.C1(n5529), 
	.B(n1401), 
	.A(n1400));
   AOI211_X2 U572 (.ZN(n13894), 
	.C2(n1420), 
	.C1(n5524), 
	.B(n1422), 
	.A(n1421));
   AOI211_X2 U578 (.ZN(n13963), 
	.C2(n1387), 
	.C1(n5525), 
	.B(n1389), 
	.A(n1388));
   AOI211_X2 U814 (.ZN(n13951), 
	.C2(n1393), 
	.C1(n5527), 
	.B(n1395), 
	.A(n1394));
   OAI222_X2 U815 (.ZN(n4924), 
	.C2(n17102), 
	.C1(n4761), 
	.B2(n16792), 
	.B1(n4821), 
	.A2(n17103), 
	.A1(FE_OFN479_n1148));
   OAI222_X2 U817 (.ZN(n4926), 
	.C2(n17102), 
	.C1(n4763), 
	.B2(n16792), 
	.B1(n4819), 
	.A2(n17103), 
	.A1(n1150));
   OAI222_X2 U829 (.ZN(n4942), 
	.C2(n17102), 
	.C1(n4772), 
	.B2(n16792), 
	.B1(n4824), 
	.A2(n17103), 
	.A1(n973));
   OAI222_X2 U830 (.ZN(n4935), 
	.C2(n17102), 
	.C1(n4850), 
	.B2(n16792), 
	.B1(n4813), 
	.A2(n318), 
	.A1(n956));
   OAI222_X2 U832 (.ZN(n4936), 
	.C2(n17102), 
	.C1(n4832), 
	.B2(n16792), 
	.B1(n4816), 
	.A2(n318), 
	.A1(n957));
   OAI222_X2 U842 (.ZN(n4938), 
	.C2(n17102), 
	.C1(n4831), 
	.B2(n16792), 
	.B1(n4815), 
	.A2(n17103), 
	.A1(n963));
   OAI222_X2 U846 (.ZN(n4923), 
	.C2(n17102), 
	.C1(n4828), 
	.B2(n16792), 
	.B1(n4825), 
	.A2(n17103), 
	.A1(n1147));
   OAI221_X2 U987 (.ZN(n4943), 
	.C2(n17102), 
	.C1(FE_PHN3661_n4852), 
	.B2(n17103), 
	.B1(n968), 
	.A(n1164));
   OAI221_X2 U1058 (.ZN(n4944), 
	.C2(n17102), 
	.C1(FE_PHN3616_n4853), 
	.B2(n17103), 
	.B1(n967), 
	.A(n1165));
   OAI221_X2 U1062 (.ZN(n5784), 
	.C2(n17102), 
	.C1(n5501), 
	.B2(n17103), 
	.B1(n871), 
	.A(n872));
   OAI221_X2 U1066 (.ZN(n5786), 
	.C2(n17102), 
	.C1(FE_PHN3598_n5500), 
	.B2(n17103), 
	.B1(n876), 
	.A(n877));
   AOI211_X2 U1070 (.ZN(n14956), 
	.C2(n1311), 
	.C1(n1310), 
	.B(n1313), 
	.A(n1312));
   AOI211_X2 U1074 (.ZN(n13758), 
	.C2(n1448), 
	.C1(n1447), 
	.B(n1450), 
	.A(n1449));
   AOI211_X2 U1078 (.ZN(n13907), 
	.C2(n1412), 
	.C1(n1411), 
	.B(n1414), 
	.A(n1413));
   OAI221_X2 U1082 (.ZN(n5714), 
	.C2(n265), 
	.C1(n268), 
	.B2(n17109), 
	.B1(FE_PHN2140_n5515), 
	.A(n269));
   OAI221_X2 U1086 (.ZN(n5720), 
	.C2(n265), 
	.C1(n280), 
	.B2(n17109), 
	.B1(FE_PHN2254_n5074), 
	.A(n281));
   OAI221_X2 U1091 (.ZN(n5725), 
	.C2(n17107), 
	.C1(n290), 
	.B2(n17109), 
	.B1(FE_PHN2376_n5571), 
	.A(n291));
   OAI221_X2 U1095 (.ZN(n5726), 
	.C2(n17107), 
	.C1(n292), 
	.B2(n17109), 
	.B1(FE_PHN2223_n5508), 
	.A(n293));
   OAI221_X2 U1100 (.ZN(n5732), 
	.C2(n17107), 
	.C1(n304), 
	.B2(n17109), 
	.B1(FE_PHN2302_n5509), 
	.A(n305));
   OAI221_X2 U1103 (.ZN(n5731), 
	.C2(n17107), 
	.C1(n302), 
	.B2(n17109), 
	.B1(FE_PHN2240_n5514), 
	.A(n303));
   OAI221_X2 U4884 (.ZN(n5730), 
	.C2(n17107), 
	.C1(n300), 
	.B2(n17109), 
	.B1(FE_PHN2180_n5517), 
	.A(n301));
endmodule

module CORTEXM0DS (
	HCLK, 
	HRESETn, 
	HADDR, 
	HBURST, 
	HMASTLOCK, 
	HPROT, 
	HSIZE, 
	HTRANS, 
	HWDATA, 
	HWRITE, 
	HRDATA, 
	HREADY, 
	HRESP, 
	NMI, 
	IRQ, 
	TXEV, 
	RXEV, 
	LOCKUP, 
	SYSRESETREQ, 
	SLEEPING, 
	FE_OFN28_HRESETn, 
	FE_OFN29_HRESETn, 
	FE_OFN30_HRESETn, 
	FE_OFN34_HRESETn, 
	FE_OFN42_HRESETn, 
	FE_OFN43_HRESETn, 
	FE_OFN55_HRESETn, 
	SPCPT1_HADDR_29_, 
	HCLK__L5_N1, 
	HCLK__L5_N13, 
	HCLK__L5_N19, 
	HCLK__L5_N2, 
	HCLK__L5_N20, 
	HCLK__L5_N21, 
	HCLK__L5_N22, 
	HCLK__L5_N23, 
	HCLK__L5_N24, 
	HCLK__L5_N25, 
	HCLK__L5_N26, 
	HCLK__L5_N27, 
	HCLK__L5_N3, 
	HCLK__L5_N39, 
	HCLK__L5_N4, 
	HCLK__L5_N5, 
	HCLK__L5_N7, 
	HCLK__L5_N8, 
	HCLK__L5_N9);
   input HCLK;
   input HRESETn;
   output [31:0] HADDR;
   output [2:0] HBURST;
   output HMASTLOCK;
   output [3:0] HPROT;
   output [2:0] HSIZE;
   output [1:0] HTRANS;
   output [31:0] HWDATA;
   output HWRITE;
   input [31:0] HRDATA;
   input HREADY;
   input HRESP;
   input NMI;
   input [15:0] IRQ;
   output TXEV;
   input RXEV;
   output LOCKUP;
   output SYSRESETREQ;
   output SLEEPING;
   input FE_OFN28_HRESETn;
   input FE_OFN29_HRESETn;
   input FE_OFN30_HRESETn;
   input FE_OFN34_HRESETn;
   input FE_OFN42_HRESETn;
   input FE_OFN43_HRESETn;
   input FE_OFN55_HRESETn;
   input SPCPT1_HADDR_29_;
   input HCLK__L5_N1;
   input HCLK__L5_N13;
   input HCLK__L5_N19;
   input HCLK__L5_N2;
   input HCLK__L5_N20;
   input HCLK__L5_N21;
   input HCLK__L5_N22;
   input HCLK__L5_N23;
   input HCLK__L5_N24;
   input HCLK__L5_N25;
   input HCLK__L5_N26;
   input HCLK__L5_N27;
   input HCLK__L5_N3;
   input HCLK__L5_N39;
   input HCLK__L5_N4;
   input HCLK__L5_N5;
   input HCLK__L5_N7;
   input HCLK__L5_N8;
   input HCLK__L5_N9;

   // Internal wires
   wire FE_UNCONNECTED_11;
   wire FE_UNCONNECTED_10;
   wire FE_UNCONNECTED_9;
   wire FE_UNCONNECTED_8;
   wire FE_UNCONNECTED_7;
   wire FE_UNCONNECTED_6;
   wire SYNOPSYS_UNCONNECTED_7;
   wire SYNOPSYS_UNCONNECTED_8;
   wire SYNOPSYS_UNCONNECTED_9;
   wire SYNOPSYS_UNCONNECTED_10;
   wire SYNOPSYS_UNCONNECTED_11;
   wire SYNOPSYS_UNCONNECTED_12;
   wire SYNOPSYS_UNCONNECTED_13;
   wire SYNOPSYS_UNCONNECTED_14;
   wire SYNOPSYS_UNCONNECTED_15;
   wire SYNOPSYS_UNCONNECTED_16;
   wire SYNOPSYS_UNCONNECTED_17;
   wire SYNOPSYS_UNCONNECTED_18;
   wire SYNOPSYS_UNCONNECTED_19;
   wire SYNOPSYS_UNCONNECTED_20;
   wire SYNOPSYS_UNCONNECTED_21;
   wire SYNOPSYS_UNCONNECTED_22;
   wire SYNOPSYS_UNCONNECTED_23;
   wire SYNOPSYS_UNCONNECTED_24;
   wire SYNOPSYS_UNCONNECTED_25;
   wire SYNOPSYS_UNCONNECTED_26;
   wire SYNOPSYS_UNCONNECTED_27;
   wire SYNOPSYS_UNCONNECTED_28;
   wire SYNOPSYS_UNCONNECTED_29;
   wire SYNOPSYS_UNCONNECTED_30;
   wire SYNOPSYS_UNCONNECTED_31;
   wire SYNOPSYS_UNCONNECTED_32;
   wire SYNOPSYS_UNCONNECTED_33;
   wire SYNOPSYS_UNCONNECTED_34;
   wire SYNOPSYS_UNCONNECTED_35;
   wire SYNOPSYS_UNCONNECTED_36;
   wire SYNOPSYS_UNCONNECTED_37;
   wire SYNOPSYS_UNCONNECTED_38;
   wire SYNOPSYS_UNCONNECTED_39;
   wire SYNOPSYS_UNCONNECTED_40;
   wire SYNOPSYS_UNCONNECTED_41;
   wire SYNOPSYS_UNCONNECTED_42;
   wire SYNOPSYS_UNCONNECTED_43;
   wire SYNOPSYS_UNCONNECTED_44;
   wire SYNOPSYS_UNCONNECTED_45;
   wire SYNOPSYS_UNCONNECTED_46;
   wire SYNOPSYS_UNCONNECTED_47;
   wire SYNOPSYS_UNCONNECTED_48;
   wire SYNOPSYS_UNCONNECTED_49;
   wire SYNOPSYS_UNCONNECTED_50;
   wire SYNOPSYS_UNCONNECTED_51;
   wire SYNOPSYS_UNCONNECTED_52;
   wire SYNOPSYS_UNCONNECTED_53;
   wire SYNOPSYS_UNCONNECTED_54;
   wire SYNOPSYS_UNCONNECTED_55;
   wire SYNOPSYS_UNCONNECTED_56;
   wire SYNOPSYS_UNCONNECTED_57;
   wire SYNOPSYS_UNCONNECTED_58;
   wire SYNOPSYS_UNCONNECTED_59;
   wire SYNOPSYS_UNCONNECTED_60;
   wire SYNOPSYS_UNCONNECTED_61;
   wire SYNOPSYS_UNCONNECTED_62;
   wire SYNOPSYS_UNCONNECTED_63;
   wire SYNOPSYS_UNCONNECTED_64;
   wire SYNOPSYS_UNCONNECTED_65;
   wire SYNOPSYS_UNCONNECTED_66;
   wire SYNOPSYS_UNCONNECTED_67;
   wire SYNOPSYS_UNCONNECTED_68;
   wire SYNOPSYS_UNCONNECTED_69;
   wire SYNOPSYS_UNCONNECTED_70;
   wire SYNOPSYS_UNCONNECTED_71;
   wire SYNOPSYS_UNCONNECTED_72;
   wire SYNOPSYS_UNCONNECTED_73;
   wire SYNOPSYS_UNCONNECTED_74;
   wire SYNOPSYS_UNCONNECTED_75;
   wire SYNOPSYS_UNCONNECTED_76;
   wire SYNOPSYS_UNCONNECTED_77;
   wire SYNOPSYS_UNCONNECTED_78;
   wire SYNOPSYS_UNCONNECTED_79;
   wire SYNOPSYS_UNCONNECTED_80;
   wire SYNOPSYS_UNCONNECTED_81;
   wire SYNOPSYS_UNCONNECTED_82;
   wire SYNOPSYS_UNCONNECTED_83;
   wire SYNOPSYS_UNCONNECTED_84;
   wire SYNOPSYS_UNCONNECTED_85;
   wire SYNOPSYS_UNCONNECTED_86;
   wire SYNOPSYS_UNCONNECTED_87;
   wire SYNOPSYS_UNCONNECTED_88;
   wire SYNOPSYS_UNCONNECTED_89;
   wire SYNOPSYS_UNCONNECTED_90;
   wire SYNOPSYS_UNCONNECTED_91;
   wire SYNOPSYS_UNCONNECTED_92;
   wire SYNOPSYS_UNCONNECTED_93;
   wire SYNOPSYS_UNCONNECTED_94;
   wire SYNOPSYS_UNCONNECTED_95;
   wire SYNOPSYS_UNCONNECTED_96;
   wire SYNOPSYS_UNCONNECTED_97;
   wire SYNOPSYS_UNCONNECTED_98;
   wire SYNOPSYS_UNCONNECTED_99;
   wire SYNOPSYS_UNCONNECTED_100;
   wire SYNOPSYS_UNCONNECTED_101;
   wire SYNOPSYS_UNCONNECTED_102;
   wire SYNOPSYS_UNCONNECTED_103;
   wire SYNOPSYS_UNCONNECTED_104;
   wire SYNOPSYS_UNCONNECTED_105;
   wire SYNOPSYS_UNCONNECTED_106;
   wire SYNOPSYS_UNCONNECTED_107;
   wire SYNOPSYS_UNCONNECTED_108;
   wire SYNOPSYS_UNCONNECTED_109;
   wire SYNOPSYS_UNCONNECTED_110;
   wire SYNOPSYS_UNCONNECTED_111;
   wire SYNOPSYS_UNCONNECTED_112;
   wire SYNOPSYS_UNCONNECTED_113;
   wire SYNOPSYS_UNCONNECTED_114;
   wire SYNOPSYS_UNCONNECTED_115;
   wire SYNOPSYS_UNCONNECTED_116;
   wire SYNOPSYS_UNCONNECTED_117;
   wire SYNOPSYS_UNCONNECTED_118;
   wire SYNOPSYS_UNCONNECTED_119;
   wire SYNOPSYS_UNCONNECTED_120;
   wire SYNOPSYS_UNCONNECTED_121;
   wire SYNOPSYS_UNCONNECTED_122;
   wire SYNOPSYS_UNCONNECTED_123;
   wire SYNOPSYS_UNCONNECTED_124;
   wire SYNOPSYS_UNCONNECTED_125;
   wire SYNOPSYS_UNCONNECTED_126;
   wire SYNOPSYS_UNCONNECTED_127;
   wire SYNOPSYS_UNCONNECTED_128;
   wire SYNOPSYS_UNCONNECTED_129;
   wire SYNOPSYS_UNCONNECTED_130;
   wire SYNOPSYS_UNCONNECTED_131;
   wire SYNOPSYS_UNCONNECTED_132;
   wire SYNOPSYS_UNCONNECTED_133;
   wire SYNOPSYS_UNCONNECTED_134;
   wire SYNOPSYS_UNCONNECTED_135;
   wire SYNOPSYS_UNCONNECTED_136;
   wire SYNOPSYS_UNCONNECTED_137;
   wire SYNOPSYS_UNCONNECTED_138;
   wire SYNOPSYS_UNCONNECTED_139;
   wire SYNOPSYS_UNCONNECTED_140;
   wire SYNOPSYS_UNCONNECTED_141;
   wire SYNOPSYS_UNCONNECTED_142;
   wire SYNOPSYS_UNCONNECTED_143;
   wire SYNOPSYS_UNCONNECTED_144;
   wire SYNOPSYS_UNCONNECTED_145;
   wire SYNOPSYS_UNCONNECTED_146;
   wire SYNOPSYS_UNCONNECTED_147;
   wire SYNOPSYS_UNCONNECTED_148;
   wire SYNOPSYS_UNCONNECTED_149;
   wire SYNOPSYS_UNCONNECTED_150;
   wire SYNOPSYS_UNCONNECTED_151;
   wire SYNOPSYS_UNCONNECTED_152;
   wire SYNOPSYS_UNCONNECTED_153;
   wire SYNOPSYS_UNCONNECTED_154;
   wire SYNOPSYS_UNCONNECTED_155;
   wire SYNOPSYS_UNCONNECTED_156;
   wire SYNOPSYS_UNCONNECTED_157;
   wire SYNOPSYS_UNCONNECTED_158;
   wire SYNOPSYS_UNCONNECTED_159;
   wire SYNOPSYS_UNCONNECTED_160;
   wire SYNOPSYS_UNCONNECTED_161;
   wire SYNOPSYS_UNCONNECTED_162;
   wire SYNOPSYS_UNCONNECTED_163;
   wire SYNOPSYS_UNCONNECTED_164;
   wire SYNOPSYS_UNCONNECTED_165;
   wire SYNOPSYS_UNCONNECTED_166;
   wire SYNOPSYS_UNCONNECTED_167;
   wire SYNOPSYS_UNCONNECTED_168;
   wire SYNOPSYS_UNCONNECTED_169;
   wire SYNOPSYS_UNCONNECTED_170;
   wire SYNOPSYS_UNCONNECTED_171;
   wire SYNOPSYS_UNCONNECTED_172;
   wire SYNOPSYS_UNCONNECTED_173;
   wire SYNOPSYS_UNCONNECTED_174;
   wire SYNOPSYS_UNCONNECTED_175;
   wire SYNOPSYS_UNCONNECTED_176;
   wire SYNOPSYS_UNCONNECTED_177;
   wire SYNOPSYS_UNCONNECTED_178;
   wire SYNOPSYS_UNCONNECTED_179;
   wire SYNOPSYS_UNCONNECTED_180;
   wire SYNOPSYS_UNCONNECTED_181;
   wire SYNOPSYS_UNCONNECTED_182;
   wire SYNOPSYS_UNCONNECTED_183;
   wire SYNOPSYS_UNCONNECTED_184;
   wire SYNOPSYS_UNCONNECTED_185;
   wire SYNOPSYS_UNCONNECTED_186;
   wire SYNOPSYS_UNCONNECTED_187;
   wire SYNOPSYS_UNCONNECTED_188;
   wire SYNOPSYS_UNCONNECTED_189;
   wire SYNOPSYS_UNCONNECTED_190;
   wire SYNOPSYS_UNCONNECTED_191;
   wire SYNOPSYS_UNCONNECTED_192;
   wire SYNOPSYS_UNCONNECTED_193;
   wire SYNOPSYS_UNCONNECTED_194;
   wire SYNOPSYS_UNCONNECTED_195;
   wire SYNOPSYS_UNCONNECTED_196;
   wire SYNOPSYS_UNCONNECTED_197;
   wire SYNOPSYS_UNCONNECTED_198;
   wire SYNOPSYS_UNCONNECTED_199;
   wire SYNOPSYS_UNCONNECTED_200;
   wire SYNOPSYS_UNCONNECTED_201;
   wire SYNOPSYS_UNCONNECTED_202;
   wire SYNOPSYS_UNCONNECTED_203;
   wire SYNOPSYS_UNCONNECTED_204;
   wire SYNOPSYS_UNCONNECTED_205;
   wire SYNOPSYS_UNCONNECTED_206;
   wire SYNOPSYS_UNCONNECTED_207;
   wire SYNOPSYS_UNCONNECTED_208;
   wire SYNOPSYS_UNCONNECTED_209;
   wire SYNOPSYS_UNCONNECTED_210;
   wire SYNOPSYS_UNCONNECTED_211;
   wire SYNOPSYS_UNCONNECTED_212;
   wire SYNOPSYS_UNCONNECTED_213;
   wire SYNOPSYS_UNCONNECTED_214;
   wire SYNOPSYS_UNCONNECTED_215;
   wire SYNOPSYS_UNCONNECTED_216;
   wire SYNOPSYS_UNCONNECTED_217;
   wire SYNOPSYS_UNCONNECTED_218;
   wire SYNOPSYS_UNCONNECTED_219;
   wire SYNOPSYS_UNCONNECTED_220;
   wire SYNOPSYS_UNCONNECTED_221;
   wire SYNOPSYS_UNCONNECTED_222;
   wire SYNOPSYS_UNCONNECTED_223;
   wire SYNOPSYS_UNCONNECTED_224;
   wire SYNOPSYS_UNCONNECTED_225;
   wire SYNOPSYS_UNCONNECTED_226;
   wire SYNOPSYS_UNCONNECTED_227;
   wire SYNOPSYS_UNCONNECTED_228;
   wire SYNOPSYS_UNCONNECTED_229;
   wire SYNOPSYS_UNCONNECTED_230;
   wire SYNOPSYS_UNCONNECTED_231;
   wire SYNOPSYS_UNCONNECTED_232;
   wire SYNOPSYS_UNCONNECTED_233;
   wire SYNOPSYS_UNCONNECTED_234;
   wire SYNOPSYS_UNCONNECTED_235;
   wire SYNOPSYS_UNCONNECTED_236;
   wire SYNOPSYS_UNCONNECTED_237;
   wire SYNOPSYS_UNCONNECTED_238;
   wire SYNOPSYS_UNCONNECTED_239;
   wire SYNOPSYS_UNCONNECTED_240;
   wire SYNOPSYS_UNCONNECTED_241;
   wire SYNOPSYS_UNCONNECTED_242;
   wire SYNOPSYS_UNCONNECTED_243;
   wire SYNOPSYS_UNCONNECTED_244;
   wire SYNOPSYS_UNCONNECTED_245;
   wire SYNOPSYS_UNCONNECTED_246;
   wire SYNOPSYS_UNCONNECTED_247;
   wire SYNOPSYS_UNCONNECTED_248;
   wire SYNOPSYS_UNCONNECTED_249;
   wire SYNOPSYS_UNCONNECTED_250;
   wire SYNOPSYS_UNCONNECTED_251;
   wire SYNOPSYS_UNCONNECTED_252;
   wire SYNOPSYS_UNCONNECTED_253;
   wire SYNOPSYS_UNCONNECTED_254;
   wire SYNOPSYS_UNCONNECTED_255;
   wire SYNOPSYS_UNCONNECTED_256;
   wire SYNOPSYS_UNCONNECTED_257;
   wire SYNOPSYS_UNCONNECTED_258;
   wire SYNOPSYS_UNCONNECTED_259;
   wire SYNOPSYS_UNCONNECTED_260;
   wire SYNOPSYS_UNCONNECTED_261;
   wire SYNOPSYS_UNCONNECTED_262;
   wire SYNOPSYS_UNCONNECTED_263;
   wire SYNOPSYS_UNCONNECTED_264;
   wire SYNOPSYS_UNCONNECTED_265;
   wire SYNOPSYS_UNCONNECTED_266;
   wire SYNOPSYS_UNCONNECTED_267;
   wire SYNOPSYS_UNCONNECTED_268;
   wire SYNOPSYS_UNCONNECTED_269;
   wire SYNOPSYS_UNCONNECTED_270;
   wire SYNOPSYS_UNCONNECTED_271;
   wire SYNOPSYS_UNCONNECTED_272;
   wire SYNOPSYS_UNCONNECTED_273;
   wire SYNOPSYS_UNCONNECTED_274;
   wire SYNOPSYS_UNCONNECTED_275;
   wire SYNOPSYS_UNCONNECTED_276;
   wire SYNOPSYS_UNCONNECTED_277;
   wire SYNOPSYS_UNCONNECTED_278;
   wire SYNOPSYS_UNCONNECTED_279;
   wire SYNOPSYS_UNCONNECTED_280;
   wire SYNOPSYS_UNCONNECTED_281;
   wire SYNOPSYS_UNCONNECTED_282;
   wire SYNOPSYS_UNCONNECTED_283;
   wire SYNOPSYS_UNCONNECTED_284;
   wire SYNOPSYS_UNCONNECTED_285;
   wire SYNOPSYS_UNCONNECTED_286;
   wire SYNOPSYS_UNCONNECTED_287;
   wire SYNOPSYS_UNCONNECTED_288;
   wire SYNOPSYS_UNCONNECTED_289;
   wire SYNOPSYS_UNCONNECTED_290;
   wire SYNOPSYS_UNCONNECTED_291;
   wire SYNOPSYS_UNCONNECTED_292;
   wire SYNOPSYS_UNCONNECTED_293;
   wire SYNOPSYS_UNCONNECTED_294;
   wire SYNOPSYS_UNCONNECTED_295;
   wire SYNOPSYS_UNCONNECTED_296;
   wire SYNOPSYS_UNCONNECTED_297;
   wire SYNOPSYS_UNCONNECTED_298;
   wire SYNOPSYS_UNCONNECTED_299;
   wire SYNOPSYS_UNCONNECTED_300;
   wire SYNOPSYS_UNCONNECTED_301;
   wire SYNOPSYS_UNCONNECTED_302;
   wire SYNOPSYS_UNCONNECTED_303;
   wire SYNOPSYS_UNCONNECTED_304;
   wire SYNOPSYS_UNCONNECTED_305;
   wire SYNOPSYS_UNCONNECTED_306;
   wire SYNOPSYS_UNCONNECTED_307;
   wire SYNOPSYS_UNCONNECTED_308;
   wire SYNOPSYS_UNCONNECTED_309;
   wire SYNOPSYS_UNCONNECTED_310;
   wire SYNOPSYS_UNCONNECTED_311;
   wire SYNOPSYS_UNCONNECTED_312;
   wire SYNOPSYS_UNCONNECTED_313;
   wire SYNOPSYS_UNCONNECTED_314;
   wire SYNOPSYS_UNCONNECTED_315;
   wire SYNOPSYS_UNCONNECTED_316;
   wire SYNOPSYS_UNCONNECTED_317;
   wire SYNOPSYS_UNCONNECTED_318;
   wire SYNOPSYS_UNCONNECTED_319;
   wire SYNOPSYS_UNCONNECTED_320;
   wire SYNOPSYS_UNCONNECTED_321;
   wire SYNOPSYS_UNCONNECTED_322;
   wire SYNOPSYS_UNCONNECTED_323;
   wire SYNOPSYS_UNCONNECTED_324;
   wire SYNOPSYS_UNCONNECTED_325;
   wire SYNOPSYS_UNCONNECTED_326;
   wire SYNOPSYS_UNCONNECTED_327;
   wire SYNOPSYS_UNCONNECTED_328;
   wire SYNOPSYS_UNCONNECTED_329;
   wire SYNOPSYS_UNCONNECTED_330;
   wire SYNOPSYS_UNCONNECTED_331;
   wire SYNOPSYS_UNCONNECTED_332;
   wire SYNOPSYS_UNCONNECTED_333;
   wire SYNOPSYS_UNCONNECTED_334;
   wire SYNOPSYS_UNCONNECTED_335;
   wire SYNOPSYS_UNCONNECTED_336;
   wire SYNOPSYS_UNCONNECTED_337;
   wire SYNOPSYS_UNCONNECTED_338;
   wire SYNOPSYS_UNCONNECTED_339;
   wire SYNOPSYS_UNCONNECTED_340;
   wire SYNOPSYS_UNCONNECTED_341;
   wire SYNOPSYS_UNCONNECTED_342;
   wire SYNOPSYS_UNCONNECTED_343;
   wire SYNOPSYS_UNCONNECTED_344;
   wire SYNOPSYS_UNCONNECTED_345;
   wire SYNOPSYS_UNCONNECTED_346;
   wire SYNOPSYS_UNCONNECTED_347;
   wire SYNOPSYS_UNCONNECTED_348;
   wire SYNOPSYS_UNCONNECTED_349;
   wire SYNOPSYS_UNCONNECTED_350;
   wire SYNOPSYS_UNCONNECTED_351;
   wire SYNOPSYS_UNCONNECTED_352;
   wire SYNOPSYS_UNCONNECTED_353;
   wire SYNOPSYS_UNCONNECTED_354;
   wire SYNOPSYS_UNCONNECTED_355;
   wire SYNOPSYS_UNCONNECTED_356;
   wire SYNOPSYS_UNCONNECTED_357;
   wire SYNOPSYS_UNCONNECTED_358;
   wire SYNOPSYS_UNCONNECTED_359;
   wire SYNOPSYS_UNCONNECTED_360;
   wire SYNOPSYS_UNCONNECTED_361;
   wire SYNOPSYS_UNCONNECTED_362;
   wire SYNOPSYS_UNCONNECTED_363;
   wire SYNOPSYS_UNCONNECTED_364;
   wire SYNOPSYS_UNCONNECTED_365;
   wire SYNOPSYS_UNCONNECTED_366;
   wire SYNOPSYS_UNCONNECTED_367;
   wire SYNOPSYS_UNCONNECTED_368;
   wire SYNOPSYS_UNCONNECTED_369;
   wire SYNOPSYS_UNCONNECTED_370;
   wire SYNOPSYS_UNCONNECTED_371;
   wire SYNOPSYS_UNCONNECTED_372;
   wire SYNOPSYS_UNCONNECTED_373;
   wire SYNOPSYS_UNCONNECTED_374;
   wire SYNOPSYS_UNCONNECTED_375;
   wire SYNOPSYS_UNCONNECTED_376;
   wire SYNOPSYS_UNCONNECTED_377;
   wire SYNOPSYS_UNCONNECTED_378;
   wire SYNOPSYS_UNCONNECTED_379;
   wire SYNOPSYS_UNCONNECTED_380;
   wire SYNOPSYS_UNCONNECTED_381;
   wire SYNOPSYS_UNCONNECTED_382;
   wire SYNOPSYS_UNCONNECTED_383;
   wire SYNOPSYS_UNCONNECTED_384;
   wire SYNOPSYS_UNCONNECTED_385;
   wire SYNOPSYS_UNCONNECTED_386;
   wire SYNOPSYS_UNCONNECTED_387;
   wire SYNOPSYS_UNCONNECTED_388;
   wire SYNOPSYS_UNCONNECTED_389;
   wire SYNOPSYS_UNCONNECTED_390;
   wire SYNOPSYS_UNCONNECTED_391;
   wire SYNOPSYS_UNCONNECTED_392;
   wire SYNOPSYS_UNCONNECTED_393;
   wire SYNOPSYS_UNCONNECTED_394;
   wire SYNOPSYS_UNCONNECTED_395;
   wire SYNOPSYS_UNCONNECTED_396;
   wire SYNOPSYS_UNCONNECTED_397;
   wire SYNOPSYS_UNCONNECTED_398;
   wire SYNOPSYS_UNCONNECTED_399;
   wire SYNOPSYS_UNCONNECTED_400;
   wire SYNOPSYS_UNCONNECTED_401;
   wire SYNOPSYS_UNCONNECTED_402;
   wire SYNOPSYS_UNCONNECTED_403;
   wire SYNOPSYS_UNCONNECTED_404;
   wire SYNOPSYS_UNCONNECTED_405;
   wire SYNOPSYS_UNCONNECTED_406;
   wire SYNOPSYS_UNCONNECTED_407;
   wire SYNOPSYS_UNCONNECTED_408;
   wire SYNOPSYS_UNCONNECTED_409;
   wire SYNOPSYS_UNCONNECTED_410;
   wire SYNOPSYS_UNCONNECTED_411;
   wire SYNOPSYS_UNCONNECTED_412;
   wire SYNOPSYS_UNCONNECTED_413;
   wire SYNOPSYS_UNCONNECTED_414;
   wire SYNOPSYS_UNCONNECTED_415;
   wire SYNOPSYS_UNCONNECTED_416;
   wire SYNOPSYS_UNCONNECTED_417;
   wire SYNOPSYS_UNCONNECTED_418;
   wire SYNOPSYS_UNCONNECTED_419;
   wire SYNOPSYS_UNCONNECTED_420;
   wire SYNOPSYS_UNCONNECTED_421;
   wire SYNOPSYS_UNCONNECTED_422;
   wire SYNOPSYS_UNCONNECTED_423;
   wire SYNOPSYS_UNCONNECTED_424;
   wire SYNOPSYS_UNCONNECTED_425;
   wire SYNOPSYS_UNCONNECTED_426;
   wire SYNOPSYS_UNCONNECTED_427;
   wire SYNOPSYS_UNCONNECTED_428;
   wire SYNOPSYS_UNCONNECTED_429;
   wire SYNOPSYS_UNCONNECTED_430;
   wire SYNOPSYS_UNCONNECTED_431;
   wire SYNOPSYS_UNCONNECTED_432;
   wire SYNOPSYS_UNCONNECTED_433;
   wire SYNOPSYS_UNCONNECTED_434;
   wire SYNOPSYS_UNCONNECTED_435;
   wire SYNOPSYS_UNCONNECTED_436;
   wire SYNOPSYS_UNCONNECTED_437;
   wire SYNOPSYS_UNCONNECTED_438;
   wire SYNOPSYS_UNCONNECTED_439;
   wire SYNOPSYS_UNCONNECTED_440;
   wire SYNOPSYS_UNCONNECTED_441;
   wire SYNOPSYS_UNCONNECTED_442;
   wire SYNOPSYS_UNCONNECTED_443;
   wire SYNOPSYS_UNCONNECTED_444;
   wire SYNOPSYS_UNCONNECTED_445;
   wire SYNOPSYS_UNCONNECTED_446;
   wire SYNOPSYS_UNCONNECTED_447;
   wire SYNOPSYS_UNCONNECTED_448;
   wire SYNOPSYS_UNCONNECTED_449;
   wire SYNOPSYS_UNCONNECTED_450;
   wire SYNOPSYS_UNCONNECTED_451;
   wire SYNOPSYS_UNCONNECTED_452;
   wire SYNOPSYS_UNCONNECTED_453;
   wire SYNOPSYS_UNCONNECTED_454;
   wire SYNOPSYS_UNCONNECTED_455;
   wire SYNOPSYS_UNCONNECTED_456;
   wire SYNOPSYS_UNCONNECTED_457;
   wire SYNOPSYS_UNCONNECTED_458;
   wire SYNOPSYS_UNCONNECTED_459;
   wire SYNOPSYS_UNCONNECTED_460;
   wire SYNOPSYS_UNCONNECTED_461;
   wire SYNOPSYS_UNCONNECTED_462;
   wire SYNOPSYS_UNCONNECTED_463;
   wire SYNOPSYS_UNCONNECTED_464;
   wire SYNOPSYS_UNCONNECTED_465;
   wire SYNOPSYS_UNCONNECTED_466;
   wire SYNOPSYS_UNCONNECTED_467;
   wire SYNOPSYS_UNCONNECTED_468;
   wire SYNOPSYS_UNCONNECTED_469;
   wire SYNOPSYS_UNCONNECTED_470;
   wire SYNOPSYS_UNCONNECTED_471;
   wire SYNOPSYS_UNCONNECTED_472;
   wire SYNOPSYS_UNCONNECTED_473;
   wire SYNOPSYS_UNCONNECTED_474;
   wire SYNOPSYS_UNCONNECTED_475;
   wire SYNOPSYS_UNCONNECTED_476;
   wire SYNOPSYS_UNCONNECTED_477;
   wire SYNOPSYS_UNCONNECTED_478;
   wire SYNOPSYS_UNCONNECTED_479;
   wire SYNOPSYS_UNCONNECTED_480;
   wire SYNOPSYS_UNCONNECTED_481;
   wire SYNOPSYS_UNCONNECTED_482;
   wire SYNOPSYS_UNCONNECTED_483;
   wire SYNOPSYS_UNCONNECTED_484;
   wire SYNOPSYS_UNCONNECTED_485;
   wire SYNOPSYS_UNCONNECTED_486;
   wire SYNOPSYS_UNCONNECTED_487;
   wire SYNOPSYS_UNCONNECTED_488;
   wire SYNOPSYS_UNCONNECTED_489;
   wire SYNOPSYS_UNCONNECTED_490;
   wire SYNOPSYS_UNCONNECTED_491;
   wire SYNOPSYS_UNCONNECTED_492;
   wire SYNOPSYS_UNCONNECTED_493;
   wire SYNOPSYS_UNCONNECTED_494;
   wire SYNOPSYS_UNCONNECTED_495;
   wire SYNOPSYS_UNCONNECTED_496;
   wire SYNOPSYS_UNCONNECTED_497;
   wire SYNOPSYS_UNCONNECTED_498;
   wire SYNOPSYS_UNCONNECTED_499;
   wire SYNOPSYS_UNCONNECTED_500;
   wire SYNOPSYS_UNCONNECTED_501;
   wire SYNOPSYS_UNCONNECTED_502;
   wire SYNOPSYS_UNCONNECTED_503;
   wire SYNOPSYS_UNCONNECTED_504;
   wire SYNOPSYS_UNCONNECTED_505;
   wire SYNOPSYS_UNCONNECTED_506;
   wire SYNOPSYS_UNCONNECTED_507;
   wire SYNOPSYS_UNCONNECTED_508;
   wire SYNOPSYS_UNCONNECTED_509;
   wire SYNOPSYS_UNCONNECTED_510;
   wire SYNOPSYS_UNCONNECTED_511;
   wire SYNOPSYS_UNCONNECTED_512;
   wire SYNOPSYS_UNCONNECTED_513;
   wire SYNOPSYS_UNCONNECTED_514;
   wire SYNOPSYS_UNCONNECTED_515;
   wire SYNOPSYS_UNCONNECTED_516;
   wire SYNOPSYS_UNCONNECTED_517;
   wire SYNOPSYS_UNCONNECTED_518;
   wire SYNOPSYS_UNCONNECTED_519;
   wire SYNOPSYS_UNCONNECTED_520;
   wire SYNOPSYS_UNCONNECTED_521;
   wire SYNOPSYS_UNCONNECTED_522;
   wire SYNOPSYS_UNCONNECTED_523;
   wire SYNOPSYS_UNCONNECTED_524;
   wire SYNOPSYS_UNCONNECTED_525;
   wire SYNOPSYS_UNCONNECTED_526;
   wire SYNOPSYS_UNCONNECTED_527;
   wire SYNOPSYS_UNCONNECTED_528;
   wire SYNOPSYS_UNCONNECTED_529;
   wire SYNOPSYS_UNCONNECTED_530;
   wire SYNOPSYS_UNCONNECTED_531;
   wire SYNOPSYS_UNCONNECTED_532;
   wire SYNOPSYS_UNCONNECTED_533;
   wire SYNOPSYS_UNCONNECTED_534;
   wire SYNOPSYS_UNCONNECTED_535;
   wire SYNOPSYS_UNCONNECTED_536;
   wire SYNOPSYS_UNCONNECTED_537;
   wire SYNOPSYS_UNCONNECTED_538;
   wire SYNOPSYS_UNCONNECTED_539;
   wire SYNOPSYS_UNCONNECTED_540;
   wire SYNOPSYS_UNCONNECTED_541;
   wire SYNOPSYS_UNCONNECTED_542;
   wire SYNOPSYS_UNCONNECTED_543;
   wire SYNOPSYS_UNCONNECTED_544;
   wire SYNOPSYS_UNCONNECTED_545;
   wire SYNOPSYS_UNCONNECTED_546;
   wire SYNOPSYS_UNCONNECTED_547;
   wire SYNOPSYS_UNCONNECTED_548;
   wire SYNOPSYS_UNCONNECTED_549;
   wire SYNOPSYS_UNCONNECTED_550;
   wire SYNOPSYS_UNCONNECTED_551;
   wire SYNOPSYS_UNCONNECTED_552;
   wire SYNOPSYS_UNCONNECTED_553;
   wire SYNOPSYS_UNCONNECTED_554;
   wire SYNOPSYS_UNCONNECTED_555;

   assign HTRANS[0] = 1'b0 ;
   assign HSIZE[2] = 1'b0 ;
   assign HPROT[1] = 1'b1 ;
   assign HMASTLOCK = 1'b0 ;
   assign HBURST[0] = 1'b0 ;
   assign HBURST[1] = 1'b0 ;
   assign HBURST[2] = 1'b0 ;

   cortexm0ds_logic u_logic (.hclk(HCLK), 
	.hreset_n(HRESETn), 
	.haddr_o(HADDR), 
	.hburst_o({ FE_UNCONNECTED_6,
		FE_UNCONNECTED_7,
		FE_UNCONNECTED_8 }), 
	.hprot_o({ HPROT[3],
		HPROT[2],
		FE_UNCONNECTED_9,
		HPROT[0] }), 
	.hsize_o({ FE_UNCONNECTED_10,
		HSIZE[1],
		HSIZE[0] }), 
	.htrans_o({ HTRANS[1],
		FE_UNCONNECTED_11 }), 
	.hwdata_o(HWDATA), 
	.hwrite_o(HWRITE), 
	.hrdata_i(HRDATA), 
	.hready_i(HREADY), 
	.hresp_i(HRESP), 
	.nmi_i(NMI), 
	.irq_i(IRQ), 
	.txev_o(TXEV), 
	.rxev_i(RXEV), 
	.lockup_o(LOCKUP), 
	.sys_reset_req_o(SYSRESETREQ), 
	.sleeping_o(SLEEPING), 
	.vis_r0_o({ SYNOPSYS_UNCONNECTED_7,
		SYNOPSYS_UNCONNECTED_8,
		SYNOPSYS_UNCONNECTED_9,
		SYNOPSYS_UNCONNECTED_10,
		SYNOPSYS_UNCONNECTED_11,
		SYNOPSYS_UNCONNECTED_12,
		SYNOPSYS_UNCONNECTED_13,
		SYNOPSYS_UNCONNECTED_14,
		SYNOPSYS_UNCONNECTED_15,
		SYNOPSYS_UNCONNECTED_16,
		SYNOPSYS_UNCONNECTED_17,
		SYNOPSYS_UNCONNECTED_18,
		SYNOPSYS_UNCONNECTED_19,
		SYNOPSYS_UNCONNECTED_20,
		SYNOPSYS_UNCONNECTED_21,
		SYNOPSYS_UNCONNECTED_22,
		SYNOPSYS_UNCONNECTED_23,
		SYNOPSYS_UNCONNECTED_24,
		SYNOPSYS_UNCONNECTED_25,
		SYNOPSYS_UNCONNECTED_26,
		SYNOPSYS_UNCONNECTED_27,
		SYNOPSYS_UNCONNECTED_28,
		SYNOPSYS_UNCONNECTED_29,
		SYNOPSYS_UNCONNECTED_30,
		SYNOPSYS_UNCONNECTED_31,
		SYNOPSYS_UNCONNECTED_32,
		SYNOPSYS_UNCONNECTED_33,
		SYNOPSYS_UNCONNECTED_34,
		SYNOPSYS_UNCONNECTED_35,
		SYNOPSYS_UNCONNECTED_36,
		SYNOPSYS_UNCONNECTED_37,
		SYNOPSYS_UNCONNECTED_38 }), 
	.vis_r1_o({ SYNOPSYS_UNCONNECTED_39,
		SYNOPSYS_UNCONNECTED_40,
		SYNOPSYS_UNCONNECTED_41,
		SYNOPSYS_UNCONNECTED_42,
		SYNOPSYS_UNCONNECTED_43,
		SYNOPSYS_UNCONNECTED_44,
		SYNOPSYS_UNCONNECTED_45,
		SYNOPSYS_UNCONNECTED_46,
		SYNOPSYS_UNCONNECTED_47,
		SYNOPSYS_UNCONNECTED_48,
		SYNOPSYS_UNCONNECTED_49,
		SYNOPSYS_UNCONNECTED_50,
		SYNOPSYS_UNCONNECTED_51,
		SYNOPSYS_UNCONNECTED_52,
		SYNOPSYS_UNCONNECTED_53,
		SYNOPSYS_UNCONNECTED_54,
		SYNOPSYS_UNCONNECTED_55,
		SYNOPSYS_UNCONNECTED_56,
		SYNOPSYS_UNCONNECTED_57,
		SYNOPSYS_UNCONNECTED_58,
		SYNOPSYS_UNCONNECTED_59,
		SYNOPSYS_UNCONNECTED_60,
		SYNOPSYS_UNCONNECTED_61,
		SYNOPSYS_UNCONNECTED_62,
		SYNOPSYS_UNCONNECTED_63,
		SYNOPSYS_UNCONNECTED_64,
		SYNOPSYS_UNCONNECTED_65,
		SYNOPSYS_UNCONNECTED_66,
		SYNOPSYS_UNCONNECTED_67,
		SYNOPSYS_UNCONNECTED_68,
		SYNOPSYS_UNCONNECTED_69,
		SYNOPSYS_UNCONNECTED_70 }), 
	.vis_r2_o({ SYNOPSYS_UNCONNECTED_71,
		SYNOPSYS_UNCONNECTED_72,
		SYNOPSYS_UNCONNECTED_73,
		SYNOPSYS_UNCONNECTED_74,
		SYNOPSYS_UNCONNECTED_75,
		SYNOPSYS_UNCONNECTED_76,
		SYNOPSYS_UNCONNECTED_77,
		SYNOPSYS_UNCONNECTED_78,
		SYNOPSYS_UNCONNECTED_79,
		SYNOPSYS_UNCONNECTED_80,
		SYNOPSYS_UNCONNECTED_81,
		SYNOPSYS_UNCONNECTED_82,
		SYNOPSYS_UNCONNECTED_83,
		SYNOPSYS_UNCONNECTED_84,
		SYNOPSYS_UNCONNECTED_85,
		SYNOPSYS_UNCONNECTED_86,
		SYNOPSYS_UNCONNECTED_87,
		SYNOPSYS_UNCONNECTED_88,
		SYNOPSYS_UNCONNECTED_89,
		SYNOPSYS_UNCONNECTED_90,
		SYNOPSYS_UNCONNECTED_91,
		SYNOPSYS_UNCONNECTED_92,
		SYNOPSYS_UNCONNECTED_93,
		SYNOPSYS_UNCONNECTED_94,
		SYNOPSYS_UNCONNECTED_95,
		SYNOPSYS_UNCONNECTED_96,
		SYNOPSYS_UNCONNECTED_97,
		SYNOPSYS_UNCONNECTED_98,
		SYNOPSYS_UNCONNECTED_99,
		SYNOPSYS_UNCONNECTED_100,
		SYNOPSYS_UNCONNECTED_101,
		SYNOPSYS_UNCONNECTED_102 }), 
	.vis_r3_o({ SYNOPSYS_UNCONNECTED_103,
		SYNOPSYS_UNCONNECTED_104,
		SYNOPSYS_UNCONNECTED_105,
		SYNOPSYS_UNCONNECTED_106,
		SYNOPSYS_UNCONNECTED_107,
		SYNOPSYS_UNCONNECTED_108,
		SYNOPSYS_UNCONNECTED_109,
		SYNOPSYS_UNCONNECTED_110,
		SYNOPSYS_UNCONNECTED_111,
		SYNOPSYS_UNCONNECTED_112,
		SYNOPSYS_UNCONNECTED_113,
		SYNOPSYS_UNCONNECTED_114,
		SYNOPSYS_UNCONNECTED_115,
		SYNOPSYS_UNCONNECTED_116,
		SYNOPSYS_UNCONNECTED_117,
		SYNOPSYS_UNCONNECTED_118,
		SYNOPSYS_UNCONNECTED_119,
		SYNOPSYS_UNCONNECTED_120,
		SYNOPSYS_UNCONNECTED_121,
		SYNOPSYS_UNCONNECTED_122,
		SYNOPSYS_UNCONNECTED_123,
		SYNOPSYS_UNCONNECTED_124,
		SYNOPSYS_UNCONNECTED_125,
		SYNOPSYS_UNCONNECTED_126,
		SYNOPSYS_UNCONNECTED_127,
		SYNOPSYS_UNCONNECTED_128,
		SYNOPSYS_UNCONNECTED_129,
		SYNOPSYS_UNCONNECTED_130,
		SYNOPSYS_UNCONNECTED_131,
		SYNOPSYS_UNCONNECTED_132,
		SYNOPSYS_UNCONNECTED_133,
		SYNOPSYS_UNCONNECTED_134 }), 
	.vis_r4_o({ SYNOPSYS_UNCONNECTED_135,
		SYNOPSYS_UNCONNECTED_136,
		SYNOPSYS_UNCONNECTED_137,
		SYNOPSYS_UNCONNECTED_138,
		SYNOPSYS_UNCONNECTED_139,
		SYNOPSYS_UNCONNECTED_140,
		SYNOPSYS_UNCONNECTED_141,
		SYNOPSYS_UNCONNECTED_142,
		SYNOPSYS_UNCONNECTED_143,
		SYNOPSYS_UNCONNECTED_144,
		SYNOPSYS_UNCONNECTED_145,
		SYNOPSYS_UNCONNECTED_146,
		SYNOPSYS_UNCONNECTED_147,
		SYNOPSYS_UNCONNECTED_148,
		SYNOPSYS_UNCONNECTED_149,
		SYNOPSYS_UNCONNECTED_150,
		SYNOPSYS_UNCONNECTED_151,
		SYNOPSYS_UNCONNECTED_152,
		SYNOPSYS_UNCONNECTED_153,
		SYNOPSYS_UNCONNECTED_154,
		SYNOPSYS_UNCONNECTED_155,
		SYNOPSYS_UNCONNECTED_156,
		SYNOPSYS_UNCONNECTED_157,
		SYNOPSYS_UNCONNECTED_158,
		SYNOPSYS_UNCONNECTED_159,
		SYNOPSYS_UNCONNECTED_160,
		SYNOPSYS_UNCONNECTED_161,
		SYNOPSYS_UNCONNECTED_162,
		SYNOPSYS_UNCONNECTED_163,
		SYNOPSYS_UNCONNECTED_164,
		SYNOPSYS_UNCONNECTED_165,
		SYNOPSYS_UNCONNECTED_166 }), 
	.vis_r5_o({ SYNOPSYS_UNCONNECTED_167,
		SYNOPSYS_UNCONNECTED_168,
		SYNOPSYS_UNCONNECTED_169,
		SYNOPSYS_UNCONNECTED_170,
		SYNOPSYS_UNCONNECTED_171,
		SYNOPSYS_UNCONNECTED_172,
		SYNOPSYS_UNCONNECTED_173,
		SYNOPSYS_UNCONNECTED_174,
		SYNOPSYS_UNCONNECTED_175,
		SYNOPSYS_UNCONNECTED_176,
		SYNOPSYS_UNCONNECTED_177,
		SYNOPSYS_UNCONNECTED_178,
		SYNOPSYS_UNCONNECTED_179,
		SYNOPSYS_UNCONNECTED_180,
		SYNOPSYS_UNCONNECTED_181,
		SYNOPSYS_UNCONNECTED_182,
		SYNOPSYS_UNCONNECTED_183,
		SYNOPSYS_UNCONNECTED_184,
		SYNOPSYS_UNCONNECTED_185,
		SYNOPSYS_UNCONNECTED_186,
		SYNOPSYS_UNCONNECTED_187,
		SYNOPSYS_UNCONNECTED_188,
		SYNOPSYS_UNCONNECTED_189,
		SYNOPSYS_UNCONNECTED_190,
		SYNOPSYS_UNCONNECTED_191,
		SYNOPSYS_UNCONNECTED_192,
		SYNOPSYS_UNCONNECTED_193,
		SYNOPSYS_UNCONNECTED_194,
		SYNOPSYS_UNCONNECTED_195,
		SYNOPSYS_UNCONNECTED_196,
		SYNOPSYS_UNCONNECTED_197,
		SYNOPSYS_UNCONNECTED_198 }), 
	.vis_r6_o({ SYNOPSYS_UNCONNECTED_199,
		SYNOPSYS_UNCONNECTED_200,
		SYNOPSYS_UNCONNECTED_201,
		SYNOPSYS_UNCONNECTED_202,
		SYNOPSYS_UNCONNECTED_203,
		SYNOPSYS_UNCONNECTED_204,
		SYNOPSYS_UNCONNECTED_205,
		SYNOPSYS_UNCONNECTED_206,
		SYNOPSYS_UNCONNECTED_207,
		SYNOPSYS_UNCONNECTED_208,
		SYNOPSYS_UNCONNECTED_209,
		SYNOPSYS_UNCONNECTED_210,
		SYNOPSYS_UNCONNECTED_211,
		SYNOPSYS_UNCONNECTED_212,
		SYNOPSYS_UNCONNECTED_213,
		SYNOPSYS_UNCONNECTED_214,
		SYNOPSYS_UNCONNECTED_215,
		SYNOPSYS_UNCONNECTED_216,
		SYNOPSYS_UNCONNECTED_217,
		SYNOPSYS_UNCONNECTED_218,
		SYNOPSYS_UNCONNECTED_219,
		SYNOPSYS_UNCONNECTED_220,
		SYNOPSYS_UNCONNECTED_221,
		SYNOPSYS_UNCONNECTED_222,
		SYNOPSYS_UNCONNECTED_223,
		SYNOPSYS_UNCONNECTED_224,
		SYNOPSYS_UNCONNECTED_225,
		SYNOPSYS_UNCONNECTED_226,
		SYNOPSYS_UNCONNECTED_227,
		SYNOPSYS_UNCONNECTED_228,
		SYNOPSYS_UNCONNECTED_229,
		SYNOPSYS_UNCONNECTED_230 }), 
	.vis_r7_o({ SYNOPSYS_UNCONNECTED_231,
		SYNOPSYS_UNCONNECTED_232,
		SYNOPSYS_UNCONNECTED_233,
		SYNOPSYS_UNCONNECTED_234,
		SYNOPSYS_UNCONNECTED_235,
		SYNOPSYS_UNCONNECTED_236,
		SYNOPSYS_UNCONNECTED_237,
		SYNOPSYS_UNCONNECTED_238,
		SYNOPSYS_UNCONNECTED_239,
		SYNOPSYS_UNCONNECTED_240,
		SYNOPSYS_UNCONNECTED_241,
		SYNOPSYS_UNCONNECTED_242,
		SYNOPSYS_UNCONNECTED_243,
		SYNOPSYS_UNCONNECTED_244,
		SYNOPSYS_UNCONNECTED_245,
		SYNOPSYS_UNCONNECTED_246,
		SYNOPSYS_UNCONNECTED_247,
		SYNOPSYS_UNCONNECTED_248,
		SYNOPSYS_UNCONNECTED_249,
		SYNOPSYS_UNCONNECTED_250,
		SYNOPSYS_UNCONNECTED_251,
		SYNOPSYS_UNCONNECTED_252,
		SYNOPSYS_UNCONNECTED_253,
		SYNOPSYS_UNCONNECTED_254,
		SYNOPSYS_UNCONNECTED_255,
		SYNOPSYS_UNCONNECTED_256,
		SYNOPSYS_UNCONNECTED_257,
		SYNOPSYS_UNCONNECTED_258,
		SYNOPSYS_UNCONNECTED_259,
		SYNOPSYS_UNCONNECTED_260,
		SYNOPSYS_UNCONNECTED_261,
		SYNOPSYS_UNCONNECTED_262 }), 
	.vis_r8_o({ SYNOPSYS_UNCONNECTED_263,
		SYNOPSYS_UNCONNECTED_264,
		SYNOPSYS_UNCONNECTED_265,
		SYNOPSYS_UNCONNECTED_266,
		SYNOPSYS_UNCONNECTED_267,
		SYNOPSYS_UNCONNECTED_268,
		SYNOPSYS_UNCONNECTED_269,
		SYNOPSYS_UNCONNECTED_270,
		SYNOPSYS_UNCONNECTED_271,
		SYNOPSYS_UNCONNECTED_272,
		SYNOPSYS_UNCONNECTED_273,
		SYNOPSYS_UNCONNECTED_274,
		SYNOPSYS_UNCONNECTED_275,
		SYNOPSYS_UNCONNECTED_276,
		SYNOPSYS_UNCONNECTED_277,
		SYNOPSYS_UNCONNECTED_278,
		SYNOPSYS_UNCONNECTED_279,
		SYNOPSYS_UNCONNECTED_280,
		SYNOPSYS_UNCONNECTED_281,
		SYNOPSYS_UNCONNECTED_282,
		SYNOPSYS_UNCONNECTED_283,
		SYNOPSYS_UNCONNECTED_284,
		SYNOPSYS_UNCONNECTED_285,
		SYNOPSYS_UNCONNECTED_286,
		SYNOPSYS_UNCONNECTED_287,
		SYNOPSYS_UNCONNECTED_288,
		SYNOPSYS_UNCONNECTED_289,
		SYNOPSYS_UNCONNECTED_290,
		SYNOPSYS_UNCONNECTED_291,
		SYNOPSYS_UNCONNECTED_292,
		SYNOPSYS_UNCONNECTED_293,
		SYNOPSYS_UNCONNECTED_294 }), 
	.vis_r9_o({ SYNOPSYS_UNCONNECTED_295,
		SYNOPSYS_UNCONNECTED_296,
		SYNOPSYS_UNCONNECTED_297,
		SYNOPSYS_UNCONNECTED_298,
		SYNOPSYS_UNCONNECTED_299,
		SYNOPSYS_UNCONNECTED_300,
		SYNOPSYS_UNCONNECTED_301,
		SYNOPSYS_UNCONNECTED_302,
		SYNOPSYS_UNCONNECTED_303,
		SYNOPSYS_UNCONNECTED_304,
		SYNOPSYS_UNCONNECTED_305,
		SYNOPSYS_UNCONNECTED_306,
		SYNOPSYS_UNCONNECTED_307,
		SYNOPSYS_UNCONNECTED_308,
		SYNOPSYS_UNCONNECTED_309,
		SYNOPSYS_UNCONNECTED_310,
		SYNOPSYS_UNCONNECTED_311,
		SYNOPSYS_UNCONNECTED_312,
		SYNOPSYS_UNCONNECTED_313,
		SYNOPSYS_UNCONNECTED_314,
		SYNOPSYS_UNCONNECTED_315,
		SYNOPSYS_UNCONNECTED_316,
		SYNOPSYS_UNCONNECTED_317,
		SYNOPSYS_UNCONNECTED_318,
		SYNOPSYS_UNCONNECTED_319,
		SYNOPSYS_UNCONNECTED_320,
		SYNOPSYS_UNCONNECTED_321,
		SYNOPSYS_UNCONNECTED_322,
		SYNOPSYS_UNCONNECTED_323,
		SYNOPSYS_UNCONNECTED_324,
		SYNOPSYS_UNCONNECTED_325,
		SYNOPSYS_UNCONNECTED_326 }), 
	.vis_r10_o({ SYNOPSYS_UNCONNECTED_327,
		SYNOPSYS_UNCONNECTED_328,
		SYNOPSYS_UNCONNECTED_329,
		SYNOPSYS_UNCONNECTED_330,
		SYNOPSYS_UNCONNECTED_331,
		SYNOPSYS_UNCONNECTED_332,
		SYNOPSYS_UNCONNECTED_333,
		SYNOPSYS_UNCONNECTED_334,
		SYNOPSYS_UNCONNECTED_335,
		SYNOPSYS_UNCONNECTED_336,
		SYNOPSYS_UNCONNECTED_337,
		SYNOPSYS_UNCONNECTED_338,
		SYNOPSYS_UNCONNECTED_339,
		SYNOPSYS_UNCONNECTED_340,
		SYNOPSYS_UNCONNECTED_341,
		SYNOPSYS_UNCONNECTED_342,
		SYNOPSYS_UNCONNECTED_343,
		SYNOPSYS_UNCONNECTED_344,
		SYNOPSYS_UNCONNECTED_345,
		SYNOPSYS_UNCONNECTED_346,
		SYNOPSYS_UNCONNECTED_347,
		SYNOPSYS_UNCONNECTED_348,
		SYNOPSYS_UNCONNECTED_349,
		SYNOPSYS_UNCONNECTED_350,
		SYNOPSYS_UNCONNECTED_351,
		SYNOPSYS_UNCONNECTED_352,
		SYNOPSYS_UNCONNECTED_353,
		SYNOPSYS_UNCONNECTED_354,
		SYNOPSYS_UNCONNECTED_355,
		SYNOPSYS_UNCONNECTED_356,
		SYNOPSYS_UNCONNECTED_357,
		SYNOPSYS_UNCONNECTED_358 }), 
	.vis_r11_o({ SYNOPSYS_UNCONNECTED_359,
		SYNOPSYS_UNCONNECTED_360,
		SYNOPSYS_UNCONNECTED_361,
		SYNOPSYS_UNCONNECTED_362,
		SYNOPSYS_UNCONNECTED_363,
		SYNOPSYS_UNCONNECTED_364,
		SYNOPSYS_UNCONNECTED_365,
		SYNOPSYS_UNCONNECTED_366,
		SYNOPSYS_UNCONNECTED_367,
		SYNOPSYS_UNCONNECTED_368,
		SYNOPSYS_UNCONNECTED_369,
		SYNOPSYS_UNCONNECTED_370,
		SYNOPSYS_UNCONNECTED_371,
		SYNOPSYS_UNCONNECTED_372,
		SYNOPSYS_UNCONNECTED_373,
		SYNOPSYS_UNCONNECTED_374,
		SYNOPSYS_UNCONNECTED_375,
		SYNOPSYS_UNCONNECTED_376,
		SYNOPSYS_UNCONNECTED_377,
		SYNOPSYS_UNCONNECTED_378,
		SYNOPSYS_UNCONNECTED_379,
		SYNOPSYS_UNCONNECTED_380,
		SYNOPSYS_UNCONNECTED_381,
		SYNOPSYS_UNCONNECTED_382,
		SYNOPSYS_UNCONNECTED_383,
		SYNOPSYS_UNCONNECTED_384,
		SYNOPSYS_UNCONNECTED_385,
		SYNOPSYS_UNCONNECTED_386,
		SYNOPSYS_UNCONNECTED_387,
		SYNOPSYS_UNCONNECTED_388,
		SYNOPSYS_UNCONNECTED_389,
		SYNOPSYS_UNCONNECTED_390 }), 
	.vis_r12_o({ SYNOPSYS_UNCONNECTED_391,
		SYNOPSYS_UNCONNECTED_392,
		SYNOPSYS_UNCONNECTED_393,
		SYNOPSYS_UNCONNECTED_394,
		SYNOPSYS_UNCONNECTED_395,
		SYNOPSYS_UNCONNECTED_396,
		SYNOPSYS_UNCONNECTED_397,
		SYNOPSYS_UNCONNECTED_398,
		SYNOPSYS_UNCONNECTED_399,
		SYNOPSYS_UNCONNECTED_400,
		SYNOPSYS_UNCONNECTED_401,
		SYNOPSYS_UNCONNECTED_402,
		SYNOPSYS_UNCONNECTED_403,
		SYNOPSYS_UNCONNECTED_404,
		SYNOPSYS_UNCONNECTED_405,
		SYNOPSYS_UNCONNECTED_406,
		SYNOPSYS_UNCONNECTED_407,
		SYNOPSYS_UNCONNECTED_408,
		SYNOPSYS_UNCONNECTED_409,
		SYNOPSYS_UNCONNECTED_410,
		SYNOPSYS_UNCONNECTED_411,
		SYNOPSYS_UNCONNECTED_412,
		SYNOPSYS_UNCONNECTED_413,
		SYNOPSYS_UNCONNECTED_414,
		SYNOPSYS_UNCONNECTED_415,
		SYNOPSYS_UNCONNECTED_416,
		SYNOPSYS_UNCONNECTED_417,
		SYNOPSYS_UNCONNECTED_418,
		SYNOPSYS_UNCONNECTED_419,
		SYNOPSYS_UNCONNECTED_420,
		SYNOPSYS_UNCONNECTED_421,
		SYNOPSYS_UNCONNECTED_422 }), 
	.vis_r14_o({ SYNOPSYS_UNCONNECTED_423,
		SYNOPSYS_UNCONNECTED_424,
		SYNOPSYS_UNCONNECTED_425,
		SYNOPSYS_UNCONNECTED_426,
		SYNOPSYS_UNCONNECTED_427,
		SYNOPSYS_UNCONNECTED_428,
		SYNOPSYS_UNCONNECTED_429,
		SYNOPSYS_UNCONNECTED_430,
		SYNOPSYS_UNCONNECTED_431,
		SYNOPSYS_UNCONNECTED_432,
		SYNOPSYS_UNCONNECTED_433,
		SYNOPSYS_UNCONNECTED_434,
		SYNOPSYS_UNCONNECTED_435,
		SYNOPSYS_UNCONNECTED_436,
		SYNOPSYS_UNCONNECTED_437,
		SYNOPSYS_UNCONNECTED_438,
		SYNOPSYS_UNCONNECTED_439,
		SYNOPSYS_UNCONNECTED_440,
		SYNOPSYS_UNCONNECTED_441,
		SYNOPSYS_UNCONNECTED_442,
		SYNOPSYS_UNCONNECTED_443,
		SYNOPSYS_UNCONNECTED_444,
		SYNOPSYS_UNCONNECTED_445,
		SYNOPSYS_UNCONNECTED_446,
		SYNOPSYS_UNCONNECTED_447,
		SYNOPSYS_UNCONNECTED_448,
		SYNOPSYS_UNCONNECTED_449,
		SYNOPSYS_UNCONNECTED_450,
		SYNOPSYS_UNCONNECTED_451,
		SYNOPSYS_UNCONNECTED_452,
		SYNOPSYS_UNCONNECTED_453,
		SYNOPSYS_UNCONNECTED_454 }), 
	.vis_msp_o({ SYNOPSYS_UNCONNECTED_455,
		SYNOPSYS_UNCONNECTED_456,
		SYNOPSYS_UNCONNECTED_457,
		SYNOPSYS_UNCONNECTED_458,
		SYNOPSYS_UNCONNECTED_459,
		SYNOPSYS_UNCONNECTED_460,
		SYNOPSYS_UNCONNECTED_461,
		SYNOPSYS_UNCONNECTED_462,
		SYNOPSYS_UNCONNECTED_463,
		SYNOPSYS_UNCONNECTED_464,
		SYNOPSYS_UNCONNECTED_465,
		SYNOPSYS_UNCONNECTED_466,
		SYNOPSYS_UNCONNECTED_467,
		SYNOPSYS_UNCONNECTED_468,
		SYNOPSYS_UNCONNECTED_469,
		SYNOPSYS_UNCONNECTED_470,
		SYNOPSYS_UNCONNECTED_471,
		SYNOPSYS_UNCONNECTED_472,
		SYNOPSYS_UNCONNECTED_473,
		SYNOPSYS_UNCONNECTED_474,
		SYNOPSYS_UNCONNECTED_475,
		SYNOPSYS_UNCONNECTED_476,
		SYNOPSYS_UNCONNECTED_477,
		SYNOPSYS_UNCONNECTED_478,
		SYNOPSYS_UNCONNECTED_479,
		SYNOPSYS_UNCONNECTED_480,
		SYNOPSYS_UNCONNECTED_481,
		SYNOPSYS_UNCONNECTED_482,
		SYNOPSYS_UNCONNECTED_483,
		SYNOPSYS_UNCONNECTED_484 }), 
	.vis_psp_o({ SYNOPSYS_UNCONNECTED_485,
		SYNOPSYS_UNCONNECTED_486,
		SYNOPSYS_UNCONNECTED_487,
		SYNOPSYS_UNCONNECTED_488,
		SYNOPSYS_UNCONNECTED_489,
		SYNOPSYS_UNCONNECTED_490,
		SYNOPSYS_UNCONNECTED_491,
		SYNOPSYS_UNCONNECTED_492,
		SYNOPSYS_UNCONNECTED_493,
		SYNOPSYS_UNCONNECTED_494,
		SYNOPSYS_UNCONNECTED_495,
		SYNOPSYS_UNCONNECTED_496,
		SYNOPSYS_UNCONNECTED_497,
		SYNOPSYS_UNCONNECTED_498,
		SYNOPSYS_UNCONNECTED_499,
		SYNOPSYS_UNCONNECTED_500,
		SYNOPSYS_UNCONNECTED_501,
		SYNOPSYS_UNCONNECTED_502,
		SYNOPSYS_UNCONNECTED_503,
		SYNOPSYS_UNCONNECTED_504,
		SYNOPSYS_UNCONNECTED_505,
		SYNOPSYS_UNCONNECTED_506,
		SYNOPSYS_UNCONNECTED_507,
		SYNOPSYS_UNCONNECTED_508,
		SYNOPSYS_UNCONNECTED_509,
		SYNOPSYS_UNCONNECTED_510,
		SYNOPSYS_UNCONNECTED_511,
		SYNOPSYS_UNCONNECTED_512,
		SYNOPSYS_UNCONNECTED_513,
		SYNOPSYS_UNCONNECTED_514 }), 
	.vis_pc_o({ SYNOPSYS_UNCONNECTED_515,
		SYNOPSYS_UNCONNECTED_516,
		SYNOPSYS_UNCONNECTED_517,
		SYNOPSYS_UNCONNECTED_518,
		SYNOPSYS_UNCONNECTED_519,
		SYNOPSYS_UNCONNECTED_520,
		SYNOPSYS_UNCONNECTED_521,
		SYNOPSYS_UNCONNECTED_522,
		SYNOPSYS_UNCONNECTED_523,
		SYNOPSYS_UNCONNECTED_524,
		SYNOPSYS_UNCONNECTED_525,
		SYNOPSYS_UNCONNECTED_526,
		SYNOPSYS_UNCONNECTED_527,
		SYNOPSYS_UNCONNECTED_528,
		SYNOPSYS_UNCONNECTED_529,
		SYNOPSYS_UNCONNECTED_530,
		SYNOPSYS_UNCONNECTED_531,
		SYNOPSYS_UNCONNECTED_532,
		SYNOPSYS_UNCONNECTED_533,
		SYNOPSYS_UNCONNECTED_534,
		SYNOPSYS_UNCONNECTED_535,
		SYNOPSYS_UNCONNECTED_536,
		SYNOPSYS_UNCONNECTED_537,
		SYNOPSYS_UNCONNECTED_538,
		SYNOPSYS_UNCONNECTED_539,
		SYNOPSYS_UNCONNECTED_540,
		SYNOPSYS_UNCONNECTED_541,
		SYNOPSYS_UNCONNECTED_542,
		SYNOPSYS_UNCONNECTED_543,
		SYNOPSYS_UNCONNECTED_544,
		SYNOPSYS_UNCONNECTED_545 }), 
	.vis_apsr_o({ SYNOPSYS_UNCONNECTED_546,
		SYNOPSYS_UNCONNECTED_547,
		SYNOPSYS_UNCONNECTED_548,
		SYNOPSYS_UNCONNECTED_549 }), 
	.vis_ipsr_o({ SYNOPSYS_UNCONNECTED_550,
		SYNOPSYS_UNCONNECTED_551,
		SYNOPSYS_UNCONNECTED_552,
		SYNOPSYS_UNCONNECTED_553,
		SYNOPSYS_UNCONNECTED_554,
		SYNOPSYS_UNCONNECTED_555 }), 
	.FE_OFN28_HRESETn(FE_OFN28_HRESETn), 
	.FE_OFN29_HRESETn(FE_OFN29_HRESETn), 
	.FE_OFN30_HRESETn(FE_OFN30_HRESETn), 
	.FE_OFN34_HRESETn(FE_OFN34_HRESETn), 
	.FE_OFN42_HRESETn(FE_OFN42_HRESETn), 
	.FE_OFN43_HRESETn(FE_OFN43_HRESETn), 
	.FE_OFN55_HRESETn(FE_OFN55_HRESETn), 
	.SPCPT1_HADDR_29_(SPCPT1_HADDR_29_), 
	.HCLK__L5_N1(HCLK__L5_N1), 
	.HCLK__L5_N13(HCLK__L5_N13), 
	.HCLK__L5_N19(HCLK__L5_N19), 
	.HCLK__L5_N2(HCLK__L5_N2), 
	.HCLK__L5_N20(HCLK__L5_N20), 
	.HCLK__L5_N21(HCLK__L5_N21), 
	.HCLK__L5_N22(HCLK__L5_N22), 
	.HCLK__L5_N23(HCLK__L5_N23), 
	.HCLK__L5_N24(HCLK__L5_N24), 
	.HCLK__L5_N25(HCLK__L5_N25), 
	.HCLK__L5_N26(HCLK__L5_N26), 
	.HCLK__L5_N27(HCLK__L5_N27), 
	.HCLK__L5_N3(HCLK__L5_N3), 
	.HCLK__L5_N39(HCLK__L5_N39), 
	.HCLK__L5_N4(HCLK__L5_N4), 
	.HCLK__L5_N5(HCLK__L5_N5), 
	.HCLK__L5_N7(HCLK__L5_N7), 
	.HCLK__L5_N8(HCLK__L5_N8), 
	.HCLK__L5_N9(HCLK__L5_N9));
endmodule

module DW_ahb (
	hclk, 
	hresetn, 
	haddr_m1, 
	hburst_m1, 
	hlock_m1, 
	hprot_m1, 
	hsize_m1, 
	htrans_m1, 
	hwdata_m1, 
	hwrite_m1, 
	hsel_s1, 
	hready_resp_s1, 
	hresp_s1, 
	hrdata_s1, 
	hsel_s2, 
	hready_resp_s2, 
	hresp_s2, 
	hrdata_s2, 
	haddr, 
	hburst, 
	hprot, 
	hsize, 
	htrans, 
	hwdata, 
	hwrite, 
	hready, 
	hresp, 
	hrdata, 
	hmaster, 
	hmaster_data, 
	hmastlock);
   input hclk;
   input hresetn;
   input [31:0] haddr_m1;
   input [2:0] hburst_m1;
   input hlock_m1;
   input [3:0] hprot_m1;
   input [2:0] hsize_m1;
   input [1:0] htrans_m1;
   input [31:0] hwdata_m1;
   input hwrite_m1;
   output hsel_s1;
   input hready_resp_s1;
   input [1:0] hresp_s1;
   input [31:0] hrdata_s1;
   output hsel_s2;
   input hready_resp_s2;
   input [1:0] hresp_s2;
   input [31:0] hrdata_s2;
   output [31:0] haddr;
   output [2:0] hburst;
   output [3:0] hprot;
   output [2:0] hsize;
   output [1:0] htrans;
   output [31:0] hwdata;
   output hwrite;
   output hready;
   output [1:0] hresp;
   output [31:0] hrdata;
   output [3:0] hmaster;
   output [3:0] hmaster_data;
   output hmastlock;

   // Internal wires
   wire hsel_3_;
   wire hready_resp_none;
   wire hresp_none_0_;
   wire U_mux_n51;
   wire U_mux_n50;
   wire U_mux_n49;
   wire U_mux_n48;
   wire U_mux_n47;
   wire U_mux_n46;
   wire U_mux_n45;
   wire U_mux_n44;
   wire U_mux_n43;
   wire U_mux_n42;
   wire U_mux_n41;
   wire U_mux_n40;
   wire U_mux_n39;
   wire U_mux_n38;
   wire U_mux_n37;
   wire U_mux_n36;
   wire U_mux_n35;
   wire U_mux_n34;
   wire U_mux_n33;
   wire U_mux_n32;
   wire U_mux_n31;
   wire U_mux_n30;
   wire U_mux_n29;
   wire U_mux_n28;
   wire U_mux_n27;
   wire U_mux_n26;
   wire U_mux_n25;
   wire U_mux_n24;
   wire U_mux_n21;
   wire U_mux_n20;
   wire U_mux_n19;
   wire U_mux_n18;
   wire U_mux_n17;
   wire U_mux_n16;
   wire U_mux_n15;
   wire U_mux_n14;
   wire U_mux_n13;
   wire U_mux_n12;
   wire U_mux_n11;
   wire U_mux_n10;
   wire U_mux_n9;
   wire U_mux_n8;
   wire U_mux_n7;
   wire U_mux_n6;
   wire U_mux_n5;
   wire U_mux_n4;
   wire U_mux_n3;
   wire U_mux_n2;
   wire U_mux_n1;
   wire U_mux_n23;
   wire U_mux_n22;
   wire U_mux_hsel_prev_1_;
   wire U_dcdr_n1;
   wire U_arblite_n1;
   wire U_dfltslv_n3;
   wire U_dfltslv_n2;
   wire U_dfltslv_n1;
   wire U_dfltslv_N4;
   wire U_dfltslv_current_state;

   assign haddr[31] = haddr_m1[31] ;
   assign haddr[30] = haddr_m1[30] ;
   assign haddr[29] = haddr_m1[29] ;
   assign haddr[28] = haddr_m1[28] ;
   assign haddr[27] = haddr_m1[27] ;
   assign haddr[26] = haddr_m1[26] ;
   assign haddr[25] = haddr_m1[25] ;
   assign haddr[24] = haddr_m1[24] ;
   assign haddr[23] = haddr_m1[23] ;
   assign haddr[22] = haddr_m1[22] ;
   assign haddr[21] = haddr_m1[21] ;
   assign haddr[20] = haddr_m1[20] ;
   assign haddr[19] = haddr_m1[19] ;
   assign haddr[18] = haddr_m1[18] ;
   assign haddr[17] = haddr_m1[17] ;
   assign haddr[16] = haddr_m1[16] ;
   assign haddr[15] = haddr_m1[15] ;
   assign haddr[14] = haddr_m1[14] ;
   assign haddr[13] = haddr_m1[13] ;
   assign haddr[12] = haddr_m1[12] ;
   assign haddr[11] = haddr_m1[11] ;
   assign haddr[10] = haddr_m1[10] ;
   assign haddr[9] = haddr_m1[9] ;
   assign haddr[8] = haddr_m1[8] ;
   assign haddr[7] = haddr_m1[7] ;
   assign haddr[6] = haddr_m1[6] ;
   assign haddr[5] = haddr_m1[5] ;
   assign haddr[4] = haddr_m1[4] ;
   assign haddr[3] = haddr_m1[3] ;
   assign haddr[2] = haddr_m1[2] ;
   assign haddr[1] = haddr_m1[1] ;
   assign haddr[0] = haddr_m1[0] ;
   assign hburst[2] = hburst_m1[2] ;
   assign hburst[1] = hburst_m1[1] ;
   assign hburst[0] = hburst_m1[0] ;
   assign hprot[3] = hprot_m1[3] ;
   assign hprot[2] = hprot_m1[2] ;
   assign hprot[1] = hprot_m1[1] ;
   assign hprot[0] = hprot_m1[0] ;
   assign hsize[2] = hsize_m1[2] ;
   assign hsize[1] = hsize_m1[1] ;
   assign hsize[0] = hsize_m1[0] ;
   assign htrans[1] = htrans_m1[1] ;
   assign htrans[0] = htrans_m1[0] ;
   assign hwdata[31] = hwdata_m1[31] ;
   assign hwdata[30] = hwdata_m1[30] ;
   assign hwdata[29] = hwdata_m1[29] ;
   assign hwdata[28] = hwdata_m1[28] ;
   assign hwdata[27] = hwdata_m1[27] ;
   assign hwdata[26] = hwdata_m1[26] ;
   assign hwdata[25] = hwdata_m1[25] ;
   assign hwdata[24] = hwdata_m1[24] ;
   assign hwdata[23] = hwdata_m1[23] ;
   assign hwdata[22] = hwdata_m1[22] ;
   assign hwdata[21] = hwdata_m1[21] ;
   assign hwdata[20] = hwdata_m1[20] ;
   assign hwdata[19] = hwdata_m1[19] ;
   assign hwdata[18] = hwdata_m1[18] ;
   assign hwdata[17] = hwdata_m1[17] ;
   assign hwdata[16] = hwdata_m1[16] ;
   assign hwdata[15] = hwdata_m1[15] ;
   assign hwdata[14] = hwdata_m1[14] ;
   assign hwdata[13] = hwdata_m1[13] ;
   assign hwdata[12] = hwdata_m1[12] ;
   assign hwdata[11] = hwdata_m1[11] ;
   assign hwdata[10] = hwdata_m1[10] ;
   assign hwdata[9] = hwdata_m1[9] ;
   assign hwdata[8] = hwdata_m1[8] ;
   assign hwdata[7] = hwdata_m1[7] ;
   assign hwdata[6] = hwdata_m1[6] ;
   assign hwdata[5] = hwdata_m1[5] ;
   assign hwdata[4] = hwdata_m1[4] ;
   assign hwdata[3] = hwdata_m1[3] ;
   assign hwdata[2] = hwdata_m1[2] ;
   assign hwdata[1] = hwdata_m1[1] ;
   assign hwdata[0] = hwdata_m1[0] ;
   assign hwrite = hwrite_m1 ;
   assign hmaster_data[1] = 1'b0 ;
   assign hmaster_data[2] = 1'b0 ;
   assign hmaster_data[3] = 1'b0 ;
   assign hmaster[1] = 1'b0 ;
   assign hmaster[2] = 1'b0 ;
   assign hmaster[3] = 1'b0 ;
   assign hmaster_data[0] = 1'b1 ;
   assign hmaster[0] = 1'b1 ;

   AOI22_X1 U_mux_U88 (.ZN(U_mux_n51), 
	.B2(hready_resp_s1), 
	.B1(U_mux_n2), 
	.A2(U_mux_n49), 
	.A1(U_mux_n50));
   OAI21_X1 U_mux_U87 (.ZN(U_mux_n23), 
	.B2(U_mux_n47), 
	.B1(hready_resp_s1), 
	.A(U_mux_n46));
   OAI22_X1 U_mux_U86 (.ZN(U_mux_n46), 
	.B2(U_mux_hsel_prev_1_), 
	.B1(U_mux_n44), 
	.A2(hsel_s1), 
	.A1(U_mux_n45));
   NOR2_X1 U_mux_U85 (.ZN(U_mux_n44), 
	.A2(U_mux_n43), 
	.A1(U_mux_n45));
   NOR2_X1 U_mux_U84 (.ZN(U_mux_n43), 
	.A2(hready_resp_none), 
	.A1(U_mux_n3));
   NAND2_X1 U_mux_U83 (.ZN(U_mux_n22), 
	.A2(U_mux_n42), 
	.A1(U_mux_n50));
   OAI221_X1 U_mux_U82 (.ZN(U_mux_n42), 
	.C2(hready_resp_s1), 
	.C1(U_mux_n49), 
	.B2(U_mux_hsel_prev_1_), 
	.B1(U_mux_n49), 
	.A(hsel_s2));
   OAI21_X1 U_mux_U81 (.ZN(U_mux_n49), 
	.B2(U_mux_n41), 
	.B1(U_mux_hsel_prev_1_), 
	.A(U_mux_n1));
   INV_X1 U_mux_U79 (.ZN(U_mux_n50), 
	.A(U_mux_n45));
   NOR2_X1 U_mux_U78 (.ZN(U_mux_n45), 
	.A2(U_mux_n1), 
	.A1(hready_resp_s2));
   OAI21_X1 U_mux_U77 (.ZN(hresp[0]), 
	.B2(U_mux_n40), 
	.B1(U_mux_hsel_prev_1_), 
	.A(U_mux_n39));
   AOI22_X1 U_mux_U76 (.ZN(U_mux_n39), 
	.B2(hresp_s1[0]), 
	.B1(U_mux_n2), 
	.A2(hresp_s2[0]), 
	.A1(U_mux_n3));
   NAND2_X1 U_mux_U75 (.ZN(U_mux_n40), 
	.A2(hresp_none_0_), 
	.A1(U_mux_n1));
   INV_X1 U_mux_U72 (.ZN(hresp[1]), 
	.A(U_mux_n38));
   AOI22_X1 U_mux_U71 (.ZN(U_mux_n38), 
	.B2(hresp_s1[1]), 
	.B1(U_mux_n2), 
	.A2(hresp_s2[1]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U70 (.ZN(hrdata[31]), 
	.A(U_mux_n37));
   AOI22_X1 U_mux_U69 (.ZN(U_mux_n37), 
	.B2(hrdata_s1[31]), 
	.B1(U_mux_n2), 
	.A2(hrdata_s2[31]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U68 (.ZN(hrdata[30]), 
	.A(U_mux_n36));
   AOI22_X1 U_mux_U67 (.ZN(U_mux_n36), 
	.B2(hrdata_s1[30]), 
	.B1(U_mux_n2), 
	.A2(hrdata_s2[30]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U66 (.ZN(hrdata[29]), 
	.A(U_mux_n35));
   AOI22_X1 U_mux_U65 (.ZN(U_mux_n35), 
	.B2(hrdata_s1[29]), 
	.B1(U_mux_n2), 
	.A2(hrdata_s2[29]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U64 (.ZN(hrdata[28]), 
	.A(U_mux_n34));
   AOI22_X1 U_mux_U63 (.ZN(U_mux_n34), 
	.B2(hrdata_s1[28]), 
	.B1(U_mux_n2), 
	.A2(hrdata_s2[28]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U62 (.ZN(hrdata[27]), 
	.A(U_mux_n33));
   AOI22_X1 U_mux_U61 (.ZN(U_mux_n33), 
	.B2(hrdata_s1[27]), 
	.B1(U_mux_n2), 
	.A2(hrdata_s2[27]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U60 (.ZN(hrdata[26]), 
	.A(U_mux_n32));
   AOI22_X1 U_mux_U59 (.ZN(U_mux_n32), 
	.B2(hrdata_s1[26]), 
	.B1(U_mux_n2), 
	.A2(hrdata_s2[26]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U58 (.ZN(hrdata[25]), 
	.A(U_mux_n31));
   AOI22_X1 U_mux_U57 (.ZN(U_mux_n31), 
	.B2(hrdata_s1[25]), 
	.B1(U_mux_n2), 
	.A2(hrdata_s2[25]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U56 (.ZN(hrdata[24]), 
	.A(U_mux_n30));
   AOI22_X1 U_mux_U55 (.ZN(U_mux_n30), 
	.B2(hrdata_s1[24]), 
	.B1(U_mux_n2), 
	.A2(hrdata_s2[24]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U54 (.ZN(hrdata[23]), 
	.A(U_mux_n29));
   AOI22_X1 U_mux_U53 (.ZN(U_mux_n29), 
	.B2(hrdata_s1[23]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[23]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U52 (.ZN(hrdata[22]), 
	.A(U_mux_n28));
   AOI22_X1 U_mux_U51 (.ZN(U_mux_n28), 
	.B2(hrdata_s1[22]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[22]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U50 (.ZN(hrdata[21]), 
	.A(U_mux_n27));
   AOI22_X1 U_mux_U49 (.ZN(U_mux_n27), 
	.B2(hrdata_s1[21]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[21]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U48 (.ZN(hrdata[20]), 
	.A(U_mux_n26));
   AOI22_X1 U_mux_U47 (.ZN(U_mux_n26), 
	.B2(hrdata_s1[20]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[20]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U46 (.ZN(hrdata[19]), 
	.A(U_mux_n25));
   AOI22_X1 U_mux_U45 (.ZN(U_mux_n25), 
	.B2(hrdata_s1[19]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[19]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U44 (.ZN(hrdata[18]), 
	.A(U_mux_n24));
   AOI22_X1 U_mux_U43 (.ZN(U_mux_n24), 
	.B2(hrdata_s1[18]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[18]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U42 (.ZN(hrdata[17]), 
	.A(U_mux_n21));
   AOI22_X1 U_mux_U41 (.ZN(U_mux_n21), 
	.B2(hrdata_s1[17]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[17]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U40 (.ZN(hrdata[16]), 
	.A(U_mux_n20));
   AOI22_X1 U_mux_U39 (.ZN(U_mux_n20), 
	.B2(hrdata_s1[16]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[16]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U38 (.ZN(hrdata[15]), 
	.A(U_mux_n19));
   AOI22_X1 U_mux_U37 (.ZN(U_mux_n19), 
	.B2(hrdata_s1[15]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[15]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U36 (.ZN(hrdata[14]), 
	.A(U_mux_n18));
   AOI22_X1 U_mux_U35 (.ZN(U_mux_n18), 
	.B2(hrdata_s1[14]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[14]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U34 (.ZN(hrdata[13]), 
	.A(U_mux_n17));
   AOI22_X1 U_mux_U33 (.ZN(U_mux_n17), 
	.B2(hrdata_s1[13]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[13]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U32 (.ZN(hrdata[12]), 
	.A(U_mux_n16));
   AOI22_X1 U_mux_U31 (.ZN(U_mux_n16), 
	.B2(hrdata_s1[12]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[12]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U30 (.ZN(hrdata[11]), 
	.A(U_mux_n15));
   AOI22_X1 U_mux_U29 (.ZN(U_mux_n15), 
	.B2(hrdata_s1[11]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[11]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U28 (.ZN(hrdata[10]), 
	.A(U_mux_n14));
   AOI22_X1 U_mux_U27 (.ZN(U_mux_n14), 
	.B2(hrdata_s1[10]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[10]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U26 (.ZN(hrdata[9]), 
	.A(U_mux_n13));
   AOI22_X1 U_mux_U25 (.ZN(U_mux_n13), 
	.B2(hrdata_s1[9]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[9]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U24 (.ZN(hrdata[8]), 
	.A(U_mux_n12));
   AOI22_X1 U_mux_U23 (.ZN(U_mux_n12), 
	.B2(hrdata_s1[8]), 
	.B1(U_mux_n2), 
	.A2(hrdata_s2[8]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U22 (.ZN(hrdata[7]), 
	.A(U_mux_n11));
   AOI22_X1 U_mux_U21 (.ZN(U_mux_n11), 
	.B2(hrdata_s1[7]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[7]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U20 (.ZN(hrdata[6]), 
	.A(U_mux_n10));
   AOI22_X1 U_mux_U19 (.ZN(U_mux_n10), 
	.B2(hrdata_s1[6]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[6]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U18 (.ZN(hrdata[5]), 
	.A(U_mux_n9));
   AOI22_X1 U_mux_U17 (.ZN(U_mux_n9), 
	.B2(hrdata_s1[5]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[5]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U16 (.ZN(hrdata[4]), 
	.A(U_mux_n8));
   AOI22_X1 U_mux_U15 (.ZN(U_mux_n8), 
	.B2(hrdata_s1[4]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[4]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U14 (.ZN(hrdata[3]), 
	.A(U_mux_n7));
   AOI22_X1 U_mux_U13 (.ZN(U_mux_n7), 
	.B2(hrdata_s1[3]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[3]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U12 (.ZN(hrdata[2]), 
	.A(U_mux_n6));
   AOI22_X1 U_mux_U11 (.ZN(U_mux_n6), 
	.B2(hrdata_s1[2]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[2]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U10 (.ZN(hrdata[1]), 
	.A(U_mux_n5));
   AOI22_X1 U_mux_U9 (.ZN(U_mux_n5), 
	.B2(hrdata_s1[1]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[1]), 
	.A1(U_mux_n3));
   INV_X1 U_mux_U8 (.ZN(hrdata[0]), 
	.A(U_mux_n4));
   AOI22_X1 U_mux_U7 (.ZN(U_mux_n4), 
	.B2(hrdata_s1[0]), 
	.B1(U_mux_n48), 
	.A2(hrdata_s2[0]), 
	.A1(U_mux_n3));
   NAND2_X1 U_mux_U6 (.ZN(U_mux_n47), 
	.A2(U_mux_n1), 
	.A1(U_mux_hsel_prev_1_));
   BUF_X1 U_mux_U5 (.Z(U_mux_n2), 
	.A(U_mux_n48));
   INV_X1 U_mux_U4 (.ZN(hready), 
	.A(U_mux_n51));
   INV_X1 U_mux_U3 (.ZN(U_mux_n48), 
	.A(U_mux_n47));
   DFFR_X2 U_mux_hsel_prev_reg_2_ (.RN(hresetn), 
	.QN(U_mux_n1), 
	.Q(U_mux_n3), 
	.D(U_mux_n22), 
	.CK(hclk));
   DFFR_X1 U_mux_hsel_prev_reg_1_ (.RN(hresetn), 
	.Q(U_mux_hsel_prev_1_), 
	.D(U_mux_n23), 
	.CK(hclk));
   NOR2_X1 U_dcdr_U6 (.ZN(hsel_s1), 
	.A2(hsel_3_), 
	.A1(haddr[30]));
   NOR2_X1 U_dcdr_U5 (.ZN(hsel_s2), 
	.A2(U_dcdr_n1), 
	.A1(hsel_3_));
   INV_X1 U_dcdr_U4 (.ZN(U_dcdr_n1), 
	.A(haddr[30]));
   OR2_X1 U_dcdr_U3 (.ZN(hsel_3_), 
	.A2(haddr[29]), 
	.A1(haddr[31]));
   MUX2_X1 U_arblite_U3 (.Z(U_arblite_n1), 
	.S(hready), 
	.B(hlock_m1), 
	.A(hmastlock));
   DFFR_X1 U_arblite_hmastlock_reg (.RN(hresetn), 
	.Q(hmastlock), 
	.D(U_arblite_n1), 
	.CK(hclk));
   OR2_X1 U_dfltslv_U5 (.ZN(U_dfltslv_n1), 
	.A2(U_dfltslv_n3), 
	.A1(U_dfltslv_current_state));
   NAND2_X1 U_dfltslv_U4 (.ZN(U_dfltslv_N4), 
	.A2(U_dfltslv_n3), 
	.A1(U_dfltslv_n2));
   NAND3_X1 U_dfltslv_U3 (.ZN(U_dfltslv_n3), 
	.A3(hsel_3_), 
	.A2(hready), 
	.A1(htrans[1]));
   DFFR_X1 U_dfltslv_hresp_none_reg_0_ (.RN(hresetn), 
	.Q(hresp_none_0_), 
	.D(U_dfltslv_N4), 
	.CK(hclk));
   DFFS_X1 U_dfltslv_current_state_reg (.SN(hresetn), 
	.QN(U_dfltslv_current_state), 
	.Q(U_dfltslv_n2), 
	.D(U_dfltslv_n1), 
	.CK(hclk));
   DFFS_X1 U_dfltslv_hready_resp_none_reg (.SN(hresetn), 
	.QN(U_mux_n41), 
	.Q(hready_resp_none), 
	.D(U_dfltslv_n1), 
	.CK(hclk));
endmodule

module cortex_soc (
	HCLK, 
	HRESETn, 
	HADDR, 
	HBURST, 
	HMASTLOCK, 
	HPROT, 
	HSIZE, 
	HTRANS, 
	HWDATA, 
	HWRITE, 
	HRDATA, 
	HREADY, 
	HRESP, 
	NMI, 
	IRQ, 
	TXEV, 
	RXEV, 
	LOCKUP, 
	SYSRESETREQ, 
	SLEEPING, 
	htrans_s, 
	hwrite_s, 
	haddr_s, 
	hsize_s, 
	hwdata_s, 
	hsel_s2, 
	hresp_s2, 
	hready_resp_s2, 
	hready_resp_s1, 
	scan_mode, 
	remap, 
	power_down, 
	clear_sr_dp, 
	big_endian, 
	debug_ad_row_addr, 
	debug_ad_bank_addr, 
	debug_ad_col_addr, 
	hsel_s1, 
	hsel_reg, 
	s_rd_data, 
	s_rd_ready, 
	hclk_2x);
   input HCLK;
   input HRESETn;
   output [31:0] HADDR;
   output [2:0] HBURST;
   output HMASTLOCK;
   output [3:0] HPROT;
   output [2:0] HSIZE;
   output [1:0] HTRANS;
   output [31:0] HWDATA;
   output HWRITE;
   input [31:0] HRDATA;
   input HREADY;
   output HRESP;
   input NMI;
   input [15:0] IRQ;
   output TXEV;
   input RXEV;
   output LOCKUP;
   output SYSRESETREQ;
   output SLEEPING;
   output [1:0] htrans_s;
   output hwrite_s;
   output [31:0] haddr_s;
   output [2:0] hsize_s;
   output [31:0] hwdata_s;
   output hsel_s2;
   input [1:0] hresp_s2;
   input hready_resp_s2;
   output hready_resp_s1;
   input scan_mode;
   input remap;
   input power_down;
   input clear_sr_dp;
   input big_endian;
   output [15:0] debug_ad_row_addr;
   output [1:0] debug_ad_bank_addr;
   output [15:0] debug_ad_col_addr;
   output hsel_s1;
   input hsel_reg;
   input [31:0] s_rd_data;
   input s_rd_ready;
   input hclk_2x;

   // Internal wires
   wire FE_PHN5235_FE_OFN27_HRESETn;
   wire FE_PHN5172_FE_OFN27_HRESETn;
   wire FE_PHN4621_FE_OFN27_HRESETn;
   wire FE_PHN2906_FE_OFN27_HRESETn;
   wire FE_PHN670_FE_OFN27_HRESETn;
   wire HCLK__L5_N39;
   wire HCLK__L5_N38;
   wire HCLK__L5_N37;
   wire HCLK__L5_N36;
   wire HCLK__L5_N35;
   wire HCLK__L5_N34;
   wire HCLK__L5_N33;
   wire HCLK__L5_N32;
   wire HCLK__L5_N31;
   wire HCLK__L5_N30;
   wire HCLK__L5_N29;
   wire HCLK__L5_N28;
   wire HCLK__L5_N27;
   wire HCLK__L5_N26;
   wire HCLK__L5_N25;
   wire HCLK__L5_N24;
   wire HCLK__L5_N23;
   wire HCLK__L5_N22;
   wire HCLK__L5_N21;
   wire HCLK__L5_N20;
   wire HCLK__L5_N19;
   wire HCLK__L5_N18;
   wire HCLK__L5_N17;
   wire HCLK__L5_N16;
   wire HCLK__L5_N15;
   wire HCLK__L5_N14;
   wire HCLK__L5_N13;
   wire HCLK__L5_N12;
   wire HCLK__L5_N11;
   wire HCLK__L5_N10;
   wire HCLK__L5_N9;
   wire HCLK__L5_N8;
   wire HCLK__L5_N7;
   wire HCLK__L5_N6;
   wire HCLK__L5_N5;
   wire HCLK__L5_N4;
   wire HCLK__L5_N3;
   wire HCLK__L5_N2;
   wire HCLK__L5_N1;
   wire HCLK__L5_N0;
   wire HCLK__L4_N7;
   wire HCLK__L4_N6;
   wire HCLK__L4_N5;
   wire HCLK__L4_N4;
   wire HCLK__L4_N3;
   wire HCLK__L4_N2;
   wire HCLK__L4_N1;
   wire HCLK__L4_N0;
   wire HCLK__L3_N1;
   wire HCLK__L3_N0;
   wire HCLK__L2_N0;
   wire HCLK__L1_N0;
   wire FE_OFN119_HADDR_31_;
   wire FE_OFN114_HADDR_29_;
   wire FE_OFN55_HRESETn;
   wire FE_OFN43_HRESETn;
   wire FE_OFN42_HRESETn;
   wire FE_OFN34_HRESETn;
   wire FE_OFN30_HRESETn;
   wire FE_OFN29_HRESETn;
   wire FE_OFN28_HRESETn;
   wire FE_OFN27_HRESETn;
   wire FE_UNCONNECTED_20;
   wire FE_UNCONNECTED_19;
   wire FE_UNCONNECTED_18;
   wire FE_UNCONNECTED_17;
   wire FE_UNCONNECTED_16;
   wire FE_UNCONNECTED_15;
   wire FE_UNCONNECTED_14;
   wire FE_UNCONNECTED_13;
   wire FE_UNCONNECTED_12;
   wire FE_UNCONNECTED_11;
   wire [1:0] hresp_s1;
   wire [31:0] hrdata_s1;
   wire [31:0] hrdata_s2;
   wire [2:0] hburst_s;
   wire [3:0] hprot_s;
   wire hready;
   wire [1:0] hresp_ahb;
   wire [31:0] hrdata;
   wire [3:0] hmaster;
   wire [3:0] hmaster_data;
   wire [15:0] s_wr_data;
   wire [15:0] s_addr;
   wire [1:0] s_bank_addr;
   wire [1:0] s_dout_valid;
   wire [0:0] s_sel_n;
   wire [1:0] s_dqm;
   wire [1:0] s_dqs;
   wire [2:0] s_sa;
   wire s_scl;
   wire [2:0] s_cas_latency;
   wire [2:0] s_read_pipe;
   wire s_sda_oe_n;
   wire [7:0] gpo;
   wire [1:0] debug_ad_sf_bank_addr;
   wire [15:0] debug_ad_sf_row_addr;
   wire [15:0] debug_ad_sf_col_addr;
   wire [31:0] debug_hiu_addr;
   wire debug_sm_burst_done;
   wire debug_sm_pop_n;
   wire debug_sm_push_n;
   wire [3:0] debug_smc_cs;
   wire debug_ref_req;
   wire s_sda_in;
   wire [7:0] gpi;
   wire [31:0] hrdata_s1_2;
   wire hready_resp_s1_2;

   assign HRESP = 1'b0 ;

   BUF_X32 FE_PHC5235_FE_OFN27_HRESETn (.Z(FE_PHN5235_FE_OFN27_HRESETn), 
	.A(FE_PHN5172_FE_OFN27_HRESETn));
   BUF_X32 FE_PHC5172_FE_OFN27_HRESETn (.Z(FE_PHN5172_FE_OFN27_HRESETn), 
	.A(FE_PHN2906_FE_OFN27_HRESETn));
   BUF_X8 FE_PHC4621_FE_OFN27_HRESETn (.Z(FE_PHN4621_FE_OFN27_HRESETn), 
	.A(FE_PHN5235_FE_OFN27_HRESETn));
   BUF_X8 FE_PHC2906_FE_OFN27_HRESETn (.Z(FE_PHN2906_FE_OFN27_HRESETn), 
	.A(FE_PHN670_FE_OFN27_HRESETn));
   BUF_X8 FE_PHC670_FE_OFN27_HRESETn (.Z(FE_PHN670_FE_OFN27_HRESETn), 
	.A(FE_OFN27_HRESETn));
   INV_X16 HCLK__L5_I39 (.ZN(HCLK__L5_N39), 
	.A(HCLK__L4_N7));
   INV_X16 HCLK__L5_I38 (.ZN(HCLK__L5_N38), 
	.A(HCLK__L4_N7));
   INV_X16 HCLK__L5_I37 (.ZN(HCLK__L5_N37), 
	.A(HCLK__L4_N7));
   INV_X16 HCLK__L5_I36 (.ZN(HCLK__L5_N36), 
	.A(HCLK__L4_N7));
   INV_X16 HCLK__L5_I35 (.ZN(HCLK__L5_N35), 
	.A(HCLK__L4_N7));
   INV_X16 HCLK__L5_I34 (.ZN(HCLK__L5_N34), 
	.A(HCLK__L4_N7));
   INV_X16 HCLK__L5_I33 (.ZN(HCLK__L5_N33), 
	.A(HCLK__L4_N7));
   INV_X16 HCLK__L5_I32 (.ZN(HCLK__L5_N32), 
	.A(HCLK__L4_N7));
   INV_X16 HCLK__L5_I31 (.ZN(HCLK__L5_N31), 
	.A(HCLK__L4_N6));
   INV_X16 HCLK__L5_I30 (.ZN(HCLK__L5_N30), 
	.A(HCLK__L4_N6));
   INV_X16 HCLK__L5_I29 (.ZN(HCLK__L5_N29), 
	.A(HCLK__L4_N6));
   INV_X16 HCLK__L5_I28 (.ZN(HCLK__L5_N28), 
	.A(HCLK__L4_N6));
   INV_X16 HCLK__L5_I27 (.ZN(HCLK__L5_N27), 
	.A(HCLK__L4_N6));
   INV_X16 HCLK__L5_I26 (.ZN(HCLK__L5_N26), 
	.A(HCLK__L4_N5));
   INV_X16 HCLK__L5_I25 (.ZN(HCLK__L5_N25), 
	.A(HCLK__L4_N5));
   INV_X16 HCLK__L5_I24 (.ZN(HCLK__L5_N24), 
	.A(HCLK__L4_N5));
   INV_X16 HCLK__L5_I23 (.ZN(HCLK__L5_N23), 
	.A(HCLK__L4_N5));
   INV_X16 HCLK__L5_I22 (.ZN(HCLK__L5_N22), 
	.A(HCLK__L4_N5));
   INV_X16 HCLK__L5_I21 (.ZN(HCLK__L5_N21), 
	.A(HCLK__L4_N5));
   INV_X16 HCLK__L5_I20 (.ZN(HCLK__L5_N20), 
	.A(HCLK__L4_N5));
   INV_X16 HCLK__L5_I19 (.ZN(HCLK__L5_N19), 
	.A(HCLK__L4_N5));
   INV_X16 HCLK__L5_I18 (.ZN(HCLK__L5_N18), 
	.A(HCLK__L4_N4));
   INV_X16 HCLK__L5_I17 (.ZN(HCLK__L5_N17), 
	.A(HCLK__L4_N4));
   INV_X16 HCLK__L5_I16 (.ZN(HCLK__L5_N16), 
	.A(HCLK__L4_N4));
   INV_X16 HCLK__L5_I15 (.ZN(HCLK__L5_N15), 
	.A(HCLK__L4_N4));
   INV_X16 HCLK__L5_I14 (.ZN(HCLK__L5_N14), 
	.A(HCLK__L4_N4));
   INV_X16 HCLK__L5_I13 (.ZN(HCLK__L5_N13), 
	.A(HCLK__L4_N4));
   INV_X16 HCLK__L5_I12 (.ZN(HCLK__L5_N12), 
	.A(HCLK__L4_N3));
   INV_X16 HCLK__L5_I11 (.ZN(HCLK__L5_N11), 
	.A(HCLK__L4_N3));
   INV_X16 HCLK__L5_I10 (.ZN(HCLK__L5_N10), 
	.A(HCLK__L4_N3));
   INV_X16 HCLK__L5_I9 (.ZN(HCLK__L5_N9), 
	.A(HCLK__L4_N2));
   INV_X16 HCLK__L5_I8 (.ZN(HCLK__L5_N8), 
	.A(HCLK__L4_N2));
   INV_X16 HCLK__L5_I7 (.ZN(HCLK__L5_N7), 
	.A(HCLK__L4_N2));
   INV_X16 HCLK__L5_I6 (.ZN(HCLK__L5_N6), 
	.A(HCLK__L4_N1));
   INV_X16 HCLK__L5_I5 (.ZN(HCLK__L5_N5), 
	.A(HCLK__L4_N1));
   INV_X16 HCLK__L5_I4 (.ZN(HCLK__L5_N4), 
	.A(HCLK__L4_N1));
   INV_X16 HCLK__L5_I3 (.ZN(HCLK__L5_N3), 
	.A(HCLK__L4_N1));
   INV_X16 HCLK__L5_I2 (.ZN(HCLK__L5_N2), 
	.A(HCLK__L4_N0));
   INV_X16 HCLK__L5_I1 (.ZN(HCLK__L5_N1), 
	.A(HCLK__L4_N0));
   INV_X16 HCLK__L5_I0 (.ZN(HCLK__L5_N0), 
	.A(HCLK__L4_N0));
   INV_X32 HCLK__L4_I7 (.ZN(HCLK__L4_N7), 
	.A(HCLK__L3_N1));
   INV_X32 HCLK__L4_I6 (.ZN(HCLK__L4_N6), 
	.A(HCLK__L3_N1));
   INV_X32 HCLK__L4_I5 (.ZN(HCLK__L4_N5), 
	.A(HCLK__L3_N1));
   INV_X32 HCLK__L4_I4 (.ZN(HCLK__L4_N4), 
	.A(HCLK__L3_N0));
   INV_X32 HCLK__L4_I3 (.ZN(HCLK__L4_N3), 
	.A(HCLK__L3_N0));
   INV_X32 HCLK__L4_I2 (.ZN(HCLK__L4_N2), 
	.A(HCLK__L3_N0));
   INV_X32 HCLK__L4_I1 (.ZN(HCLK__L4_N1), 
	.A(HCLK__L3_N0));
   INV_X32 HCLK__L4_I0 (.ZN(HCLK__L4_N0), 
	.A(HCLK__L3_N0));
   INV_X32 HCLK__L3_I1 (.ZN(HCLK__L3_N1), 
	.A(HCLK__L2_N0));
   INV_X32 HCLK__L3_I0 (.ZN(HCLK__L3_N0), 
	.A(HCLK__L2_N0));
   BUF_X8 HCLK__L2_I0 (.Z(HCLK__L2_N0), 
	.A(HCLK__L1_N0));
   INV_X32 HCLK__L1_I0 (.ZN(HCLK__L1_N0), 
	.A(HCLK));
   INV_X1 FE_OFC120_HADDR_31_ (.ZN(HADDR[31]), 
	.A(FE_OFN119_HADDR_31_));
   INV_X4 FE_OFC115_HADDR_29_ (.ZN(HADDR[29]), 
	.A(FE_OFN114_HADDR_29_));
   BUF_X8 FE_OFC55_HRESETn (.Z(FE_OFN55_HRESETn), 
	.A(FE_OFN34_HRESETn));
   BUF_X8 FE_OFC43_HRESETn (.Z(FE_OFN43_HRESETn), 
	.A(FE_OFN28_HRESETn));
   BUF_X8 FE_OFC42_HRESETn (.Z(FE_OFN42_HRESETn), 
	.A(FE_OFN28_HRESETn));
   INV_X16 FE_OFC34_HRESETn (.ZN(FE_OFN34_HRESETn), 
	.A(FE_PHN4621_FE_OFN27_HRESETn));
   INV_X4 FE_OFC30_HRESETn (.ZN(FE_OFN30_HRESETn), 
	.A(FE_PHN4621_FE_OFN27_HRESETn));
   INV_X4 FE_OFC29_HRESETn (.ZN(FE_OFN29_HRESETn), 
	.A(FE_PHN4621_FE_OFN27_HRESETn));
   INV_X8 FE_OFC28_HRESETn (.ZN(FE_OFN28_HRESETn), 
	.A(FE_PHN4621_FE_OFN27_HRESETn));
   INV_X8 FE_OFC27_HRESETn (.ZN(FE_OFN27_HRESETn), 
	.A(HRESETn));
   AHB_Lite_2s ahb (.HCLK(HCLK), 
	.HRESETn(HRESETn), 
	.HADDR(HADDR), 
	.HBURST(HBURST), 
	.HMASTLOCK(HMASTLOCK), 
	.HPROT(HPROT), 
	.HSIZE(HSIZE), 
	.HTRANS(HTRANS), 
	.HWDATA(HWDATA), 
	.HWRITE(HWRITE), 
	.hsel_s1(hsel_s1), 
	.hready_resp_s1(hready_resp_s1), 
	.hresp_s1(hresp_s1), 
	.hrdata_s1(hrdata_s1), 
	.hsel_s2(hsel_s2), 
	.hready_resp_s2(hready_resp_s2), 
	.hresp_s2(hresp_s2), 
	.hrdata_s2(hrdata_s2), 
	.haddr_s(haddr_s), 
	.hburst_s(hburst_s), 
	.hprot_s(hprot_s), 
	.hsize_s(hsize_s), 
	.htrans_s(htrans_s), 
	.hwdata_s(hwdata_s), 
	.hwrite_s(hwrite_s), 
	.HREADY(HREADY), 
	.hresp_ahb(hresp_ahb), 
	.HRDATA(HRDATA), 
	.hmaster(hmaster), 
	.hmaster_data(hmaster_data), 
	.hmastlock_s(FE_UNCONNECTED_11), 
	.FE_OFN114_HADDR_29_(FE_OFN114_HADDR_29_), 
	.FE_OFN119_HADDR_31_(FE_OFN119_HADDR_31_));
   DW_memctl memctl_v4 (.hready_resp(hready_resp_s1), 
	.hresp(hresp_s1), 
	.hrdata(hrdata_s1), 
	.s_ras_n(FE_UNCONNECTED_12), 
	.s_cas_n(FE_UNCONNECTED_13), 
	.s_cke(FE_UNCONNECTED_14), 
	.s_wr_data(s_wr_data), 
	.s_addr(s_addr), 
	.s_bank_addr(s_bank_addr), 
	.s_dout_valid(s_dout_valid), 
	.s_sel_n(s_sel_n), 
	.s_dqm(s_dqm), 
	.s_we_n(FE_UNCONNECTED_15), 
	.s_dqs(s_dqs), 
	.s_sa(s_sa), 
	.s_scl(s_scl), 
	.s_rd_ready(s_rd_ready), 
	.s_rd_start(FE_UNCONNECTED_16), 
	.s_rd_pop(FE_UNCONNECTED_17), 
	.s_rd_end(FE_UNCONNECTED_18), 
	.s_rd_dqs_mask(FE_UNCONNECTED_19), 
	.s_cas_latency(s_cas_latency), 
	.s_read_pipe(s_read_pipe), 
	.s_sda_out(FE_UNCONNECTED_20), 
	.s_sda_oe_n(s_sda_oe_n), 
	.gpo(gpo), 
	.debug_ad_bank_addr(debug_ad_bank_addr), 
	.debug_ad_row_addr(debug_ad_row_addr), 
	.debug_ad_col_addr(debug_ad_col_addr), 
	.debug_ad_sf_bank_addr(debug_ad_sf_bank_addr), 
	.debug_ad_sf_row_addr(debug_ad_sf_row_addr), 
	.debug_ad_sf_col_addr(debug_ad_sf_col_addr), 
	.debug_hiu_addr(debug_hiu_addr), 
	.debug_sm_burst_done(debug_sm_burst_done), 
	.debug_sm_pop_n(debug_sm_pop_n), 
	.debug_sm_push_n(debug_sm_push_n), 
	.debug_smc_cs(debug_smc_cs), 
	.debug_ref_req(debug_ref_req), 
	.hclk(HCLK__L5_N10), 
	.hclk_2x(hclk_2x), 
	.hresetn(FE_PHN4621_FE_OFN27_HRESETn), 
	.scan_mode(scan_mode), 
	.haddr(haddr_s), 
	.hsel_mem(hsel_s1), 
	.hsel_reg(hsel_reg), 
	.hwrite(hwrite_s), 
	.htrans(htrans_s), 
	.hsize(hsize_s), 
	.hburst(hburst_s), 
	.hready(HREADY), 
	.hwdata(hwdata_s), 
	.s_rd_data(s_rd_data), 
	.s_sda_in(s_sda_in), 
	.gpi(gpi), 
	.remap(remap), 
	.power_down(power_down), 
	.clear_sr_dp(clear_sr_dp), 
	.big_endian(big_endian), 
	.FE_OFN28_HRESETn(FE_OFN28_HRESETn), 
	.FE_OFN29_HRESETn(FE_OFN29_HRESETn), 
	.FE_OFN30_HRESETn(FE_OFN30_HRESETn), 
	.FE_OFN34_HRESETn(FE_OFN34_HRESETn), 
	.FE_OFN42_HRESETn(FE_OFN42_HRESETn), 
	.FE_OFN43_HRESETn(FE_OFN43_HRESETn), 
	.FE_OFN55_HRESETn(FE_OFN55_HRESETn), 
	.HCLK__L5_N11(HCLK__L5_N11), 
	.HCLK__L5_N12(HCLK__L5_N12), 
	.HCLK__L5_N13(HCLK__L5_N13), 
	.HCLK__L5_N14(HCLK__L5_N14), 
	.HCLK__L5_N15(HCLK__L5_N15), 
	.HCLK__L5_N16(HCLK__L5_N16), 
	.HCLK__L5_N17(HCLK__L5_N17), 
	.HCLK__L5_N18(HCLK__L5_N18), 
	.HCLK__L5_N27(HCLK__L5_N27), 
	.HCLK__L5_N28(HCLK__L5_N28), 
	.HCLK__L5_N29(HCLK__L5_N29), 
	.HCLK__L5_N30(HCLK__L5_N30), 
	.HCLK__L5_N31(HCLK__L5_N31), 
	.HCLK__L5_N32(HCLK__L5_N32), 
	.HCLK__L5_N33(HCLK__L5_N33), 
	.HCLK__L5_N34(HCLK__L5_N34), 
	.HCLK__L5_N35(HCLK__L5_N35), 
	.HCLK__L5_N36(HCLK__L5_N36), 
	.HCLK__L5_N37(HCLK__L5_N37), 
	.HCLK__L5_N38(HCLK__L5_N38), 
	.HCLK__L5_N39(HCLK__L5_N39), 
	.HCLK__L5_N4(HCLK__L5_N4), 
	.HCLK__L5_N5(HCLK__L5_N5), 
	.HCLK__L5_N6(HCLK__L5_N6));
   CORTEXM0DS u_cortexm0ds (.HCLK(HCLK__L5_N0), 
	.HRESETn(FE_PHN4621_FE_OFN27_HRESETn), 
	.HADDR({ FE_OFN119_HADDR_31_,
		HADDR[30],
		FE_OFN114_HADDR_29_,
		HADDR[28],
		HADDR[27],
		HADDR[26],
		HADDR[25],
		HADDR[24],
		HADDR[23],
		HADDR[22],
		HADDR[21],
		HADDR[20],
		HADDR[19],
		HADDR[18],
		HADDR[17],
		HADDR[16],
		HADDR[15],
		HADDR[14],
		HADDR[13],
		HADDR[12],
		HADDR[11],
		HADDR[10],
		HADDR[9],
		HADDR[8],
		HADDR[7],
		HADDR[6],
		HADDR[5],
		HADDR[4],
		HADDR[3],
		HADDR[2],
		HADDR[1],
		HADDR[0] }), 
	.HBURST(HBURST), 
	.HMASTLOCK(HMASTLOCK), 
	.HPROT(HPROT), 
	.HSIZE(HSIZE), 
	.HTRANS(HTRANS), 
	.HWDATA(HWDATA), 
	.HWRITE(HWRITE), 
	.HRDATA(HRDATA), 
	.HREADY(HREADY), 
	.HRESP(HRESP), 
	.NMI(NMI), 
	.IRQ(IRQ), 
	.TXEV(TXEV), 
	.RXEV(RXEV), 
	.LOCKUP(LOCKUP), 
	.SYSRESETREQ(SYSRESETREQ), 
	.SLEEPING(SLEEPING), 
	.FE_OFN28_HRESETn(FE_OFN28_HRESETn), 
	.FE_OFN29_HRESETn(FE_OFN29_HRESETn), 
	.FE_OFN30_HRESETn(FE_OFN30_HRESETn), 
	.FE_OFN34_HRESETn(FE_OFN34_HRESETn), 
	.FE_OFN42_HRESETn(FE_OFN42_HRESETn), 
	.FE_OFN43_HRESETn(FE_OFN43_HRESETn), 
	.FE_OFN55_HRESETn(FE_OFN55_HRESETn), 
	.SPCPT1_HADDR_29_(HADDR[29]), 
	.HCLK__L5_N1(HCLK__L5_N1), 
	.HCLK__L5_N13(HCLK__L5_N13), 
	.HCLK__L5_N19(HCLK__L5_N19), 
	.HCLK__L5_N2(HCLK__L5_N2), 
	.HCLK__L5_N20(HCLK__L5_N20), 
	.HCLK__L5_N21(HCLK__L5_N21), 
	.HCLK__L5_N22(HCLK__L5_N22), 
	.HCLK__L5_N23(HCLK__L5_N23), 
	.HCLK__L5_N24(HCLK__L5_N24), 
	.HCLK__L5_N25(HCLK__L5_N25), 
	.HCLK__L5_N26(HCLK__L5_N26), 
	.HCLK__L5_N27(HCLK__L5_N27), 
	.HCLK__L5_N3(HCLK__L5_N3), 
	.HCLK__L5_N39(HCLK__L5_N39), 
	.HCLK__L5_N4(HCLK__L5_N4), 
	.HCLK__L5_N5(HCLK__L5_N5), 
	.HCLK__L5_N7(HCLK__L5_N7), 
	.HCLK__L5_N8(HCLK__L5_N8), 
	.HCLK__L5_N9(HCLK__L5_N9));
endmodule

