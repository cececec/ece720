
module DW_memctl_hiu ( hclk, hresetn, hsel_mem, hsel_reg, htrans, hwrite, 
        hsize, hburst, hready, hready_resp, hresp, haddr, hwdata, hrdata, 
        hiu_req, hiu_burst_size, hiu_wrap_burst, hiu_rw, hiu_terminate, 
        hiu_addr, hiu_data, hiu_haddr, hiu_hsize, miu_burst_done, miu_push_n, 
        miu_pop_n, miu_data, miu_data_width, miu_col_width, big_endian );
  input [1:0] htrans;
  input [2:0] hsize;
  input [2:0] hburst;
  output [1:0] hresp;
  input [31:0] haddr;
  input [31:0] hwdata;
  output [31:0] hrdata;
  output [1:0] hiu_req;
  output [5:0] hiu_burst_size;
  output [31:0] hiu_addr;
  output [31:0] hiu_data;
  output [3:0] hiu_haddr;
  output [2:0] hiu_hsize;
  input [31:0] miu_data;
  input [1:0] miu_data_width;
  input [3:0] miu_col_width;
  input hclk, hresetn, hsel_mem, hsel_reg, hwrite, hready, miu_burst_done,
         miu_push_n, miu_pop_n, big_endian;
  output hready_resp, hiu_wrap_burst, hiu_rw, hiu_terminate;
  wire   m_af_push1_n, m_af_data1_in_13_, m_af_data1_in_11_, m_af_data1_in_9_,
         m_af_data1_in_8_, m_af_data1_in_7_, m_af_data1_in_6_,
         m_af_data1_in_5_, m_af_data1_in_4_, m_af_data1_in_3_,
         m_af_data1_in_2_, m_af_data1_in_0_, m_af_ready, m_af_new_req,
         m_af_dummy_req, m_df_push_n, m_df_ready, m_df_wr_term, m_two_to_one,
         m_rb_start, m_rb_done, m_rb_busy, m_rb_pop_n, m_rb_sel_buf, m_double,
         m_rb_ready, m_rb_overflow, n7, n8, U_afifo_n259, U_afifo_n258,
         U_afifo_n257, U_afifo_n256, U_afifo_n255, U_afifo_n253, U_afifo_n252,
         U_afifo_n250, U_afifo_n248, U_afifo_n246, U_afifo_n245, U_afifo_n244,
         U_afifo_n243, U_afifo_n242, U_afifo_n241, U_afifo_n240, U_afifo_n239,
         U_afifo_n238, U_afifo_n237, U_afifo_n236, U_afifo_n235, U_afifo_n234,
         U_afifo_n233, U_afifo_n232, U_afifo_n231, U_afifo_n230, U_afifo_n229,
         U_afifo_n228, U_afifo_n227, U_afifo_n226, U_afifo_n225, U_afifo_n224,
         U_afifo_n223, U_afifo_n222, U_afifo_n221, U_afifo_n220, U_afifo_n219,
         U_afifo_n218, U_afifo_n217, U_afifo_n216, U_afifo_n215, U_afifo_n214,
         U_afifo_n213, U_afifo_n212, U_afifo_n211, U_afifo_n210, U_afifo_n209,
         U_afifo_n208, U_afifo_n207, U_afifo_n206, U_afifo_n205, U_afifo_n204,
         U_afifo_n203, U_afifo_n202, U_afifo_n201, U_afifo_n200, U_afifo_n198,
         U_afifo_n196, U_afifo_n195, U_afifo_n194, U_afifo_n192, U_afifo_n191,
         U_afifo_n190, U_afifo_n188, U_afifo_n187, U_afifo_n186, U_afifo_n185,
         U_afifo_n184, U_afifo_n183, U_afifo_n182, U_afifo_n181, U_afifo_n180,
         U_afifo_n179, U_afifo_n178, U_afifo_n176, U_afifo_n174, U_afifo_n173,
         U_afifo_n172, U_afifo_n171, U_afifo_n170, U_afifo_n169, U_afifo_n168,
         U_afifo_n167, U_afifo_n166, U_afifo_n165, U_afifo_n164, U_afifo_n163,
         U_afifo_n162, U_afifo_n161, U_afifo_n160, U_afifo_n159, U_afifo_n158,
         U_afifo_n157, U_afifo_n156, U_afifo_n155, U_afifo_n154, U_afifo_n153,
         U_afifo_n152, U_afifo_n151, U_afifo_n147, U_afifo_n140, U_afifo_n138,
         U_afifo_n137, U_afifo_n99, U_afifo_n98, U_afifo_n93, U_afifo_n85,
         U_afifo_n84, U_afifo_n76, U_afifo_n75, U_afifo_n54, U_afifo_n49,
         U_afifo_n15, U_afifo_n14, U_afifo_n13, U_afifo_n11, U_afifo_n10,
         U_afifo_n9, U_afifo_n7, U_afifo_n5, U_afifo_n1, U_afifo_n65,
         U_afifo_n55, U_afifo_n52, U_afifo_n51, U_afifo_n48, U_afifo_n47,
         U_afifo_n46, U_afifo_n45, U_afifo_n44, U_afifo_n43, U_afifo_n42,
         U_afifo_n41, U_afifo_n40, U_afifo_n39, U_afifo_n38, U_afifo_n37,
         U_afifo_n36, U_afifo_n35, U_afifo_n34, U_afifo_n33, U_afifo_n32,
         U_afifo_n31, U_afifo_n30, U_afifo_n29, U_afifo_n28, U_afifo_n27,
         U_afifo_n26, U_afifo_n25, U_afifo_n24, U_afifo_n23, U_afifo_n22,
         U_afifo_n21, U_afifo_n20, U_afifo_n19, U_afifo_n18, U_afifo_n17,
         U_afifo_n16, U_afifo_n12, U_afifo_n8, U_afifo_n6, U_afifo_n4,
         U_afifo_n3, U_afifo_n2, U_afifo_n_new_req, U_afifo_f_clr_pers,
         U_afifo_f_core_ready, U_afifo_f_data2_0_, U_afifo_f_data2_2_,
         U_afifo_f_data2_4_, U_afifo_f_data2_5_, U_afifo_f_data2_6_,
         U_afifo_f_data2_7_, U_afifo_f_data2_8_, U_afifo_f_data2_12_,
         U_afifo_f_data2_13_, U_afifo_f_data2_14_, U_afifo_f_data2_15_,
         U_afifo_f_data2_16_, U_afifo_f_data2_17_, U_afifo_f_data2_18_,
         U_afifo_f_data2_19_, U_afifo_f_data2_20_, U_afifo_f_data2_21_,
         U_afifo_f_data2_22_, U_afifo_f_data2_23_, U_afifo_f_data2_24_,
         U_afifo_f_data2_25_, U_afifo_f_data2_26_, U_afifo_f_data2_27_,
         U_afifo_f_data2_28_, U_afifo_f_data2_29_, U_afifo_f_data2_30_,
         U_afifo_f_data2_31_, U_afifo_f_data2_32_, U_afifo_f_data2_33_,
         U_afifo_f_data2_34_, U_afifo_f_data2_35_, U_afifo_f_data2_36_,
         U_afifo_f_data2_37_, U_afifo_f_data2_38_, U_afifo_f_data2_39_,
         U_afifo_f_data2_40_, U_afifo_f_data2_41_, U_afifo_f_data2_42_,
         U_afifo_f_data2_43_, U_afifo_f_data2_44_, U_afifo_f_data2_47_,
         U_afifo_f_data2_48_, U_afifo_f_push2_pending, U_afifo_m_data_out_0_,
         U_afifo_m_data_out_3, U_afifo_m_data_out_49, U_afifo_m_full,
         U_afifo_m_afull, U_afifo_m_aempty, U_afifo_m_empty, U_afifo_m_pop_n,
         U_dfifo_n4, U_dfifo_n2, U_dfifo_n5, U_dfifo_n3, U_dfifo_f_1st_half,
         U_dfifo_m_full, U_dfifo_m_afull, U_dfifo_m_aempty, U_dfifo_m_empty,
         U_dfifo_m_data_out_0_, U_dfifo_m_data_out_1_, U_rbuf_n198,
         U_rbuf_n197, U_rbuf_n196, U_rbuf_n195, U_rbuf_n194, U_rbuf_n193,
         U_rbuf_n192, U_rbuf_n191, U_rbuf_n190, U_rbuf_n189, U_rbuf_n188,
         U_rbuf_n187, U_rbuf_n186, U_rbuf_n185, U_rbuf_n184, U_rbuf_n183,
         U_rbuf_n182, U_rbuf_n181, U_rbuf_n180, U_rbuf_n179, U_rbuf_n178,
         U_rbuf_n177, U_rbuf_n176, U_rbuf_n175, U_rbuf_n174, U_rbuf_n173,
         U_rbuf_n172, U_rbuf_n171, U_rbuf_n170, U_rbuf_n169, U_rbuf_n168,
         U_rbuf_n167, U_rbuf_n166, U_rbuf_n165, U_rbuf_n164, U_rbuf_n163,
         U_rbuf_n162, U_rbuf_n161, U_rbuf_n160, U_rbuf_n159, U_rbuf_n158,
         U_rbuf_n157, U_rbuf_n156, U_rbuf_n155, U_rbuf_n154, U_rbuf_n152,
         U_rbuf_n151, U_rbuf_n150, U_rbuf_n149, U_rbuf_n148, U_rbuf_n146,
         U_rbuf_n145, U_rbuf_n143, U_rbuf_n142, U_rbuf_n141, U_rbuf_n140,
         U_rbuf_n139, U_rbuf_n138, U_rbuf_n137, U_rbuf_n136, U_rbuf_n135,
         U_rbuf_n134, U_rbuf_n133, U_rbuf_n132, U_rbuf_n131, U_rbuf_n130,
         U_rbuf_n129, U_rbuf_n128, U_rbuf_n127, U_rbuf_n126, U_rbuf_n125,
         U_rbuf_n124, U_rbuf_n123, U_rbuf_n120, U_rbuf_n119, U_rbuf_n118,
         U_rbuf_n117, U_rbuf_n116, U_rbuf_n115, U_rbuf_n114, U_rbuf_n113,
         U_rbuf_n112, U_rbuf_n111, U_rbuf_n110, U_rbuf_n109, U_rbuf_n108,
         U_rbuf_n107, U_rbuf_n106, U_rbuf_n105, U_rbuf_n104, U_rbuf_n103,
         U_rbuf_n102, U_rbuf_n101, U_rbuf_n100, U_rbuf_n99, U_rbuf_n98,
         U_rbuf_n97, U_rbuf_n96, U_rbuf_n95, U_rbuf_n94, U_rbuf_n93,
         U_rbuf_n92, U_rbuf_n91, U_rbuf_n90, U_rbuf_n54, U_rbuf_n53,
         U_rbuf_n52, U_rbuf_n51, U_rbuf_n50, U_rbuf_n49, U_rbuf_n48,
         U_rbuf_n47, U_rbuf_n46, U_rbuf_n45, U_rbuf_n44, U_rbuf_n43,
         U_rbuf_n42, U_rbuf_n41, U_rbuf_n40, U_rbuf_n39, U_rbuf_n38,
         U_rbuf_n35, U_rbuf_n34, U_rbuf_n33, U_rbuf_n32, U_rbuf_n31,
         U_rbuf_n30, U_rbuf_n29, U_rbuf_n28, U_rbuf_n27, U_rbuf_n26,
         U_rbuf_n25, U_rbuf_n24, U_rbuf_n23, U_rbuf_n22, U_rbuf_n21,
         U_rbuf_n20, U_rbuf_n19, U_rbuf_n18, U_rbuf_n17, U_rbuf_n16,
         U_rbuf_n15, U_rbuf_n9, U_rbuf_n8, U_rbuf_n7, U_rbuf_n6, U_rbuf_n4,
         U_rbuf_n3, U_rbuf_n89, U_rbuf_n88, U_rbuf_n87, U_rbuf_n86, U_rbuf_n85,
         U_rbuf_n84, U_rbuf_n83, U_rbuf_n82, U_rbuf_n81, U_rbuf_n80,
         U_rbuf_n79, U_rbuf_n78, U_rbuf_n77, U_rbuf_n76, U_rbuf_n75,
         U_rbuf_n74, U_rbuf_n73, U_rbuf_n72, U_rbuf_n71, U_rbuf_n70,
         U_rbuf_n69, U_rbuf_n68, U_rbuf_n67, U_rbuf_n66, U_rbuf_n65,
         U_rbuf_n64, U_rbuf_n63, U_rbuf_n62, U_rbuf_n61, U_rbuf_n60,
         U_rbuf_n59, U_rbuf_n58, U_rbuf_n57, U_rbuf_n56, U_rbuf_n55,
         U_rbuf_f_top_data_0_, U_rbuf_f_top_data_1_, U_rbuf_f_top_data_2_,
         U_rbuf_f_top_data_3_, U_rbuf_f_top_data_4_, U_rbuf_f_top_data_5_,
         U_rbuf_f_top_data_6_, U_rbuf_f_top_data_7_, U_rbuf_f_top_data_8_,
         U_rbuf_f_top_data_9_, U_rbuf_f_top_data_10_, U_rbuf_f_top_data_11_,
         U_rbuf_f_top_data_12_, U_rbuf_f_top_data_13_, U_rbuf_f_top_data_14_,
         U_rbuf_f_top_data_15_, U_rbuf_f_1st_half, U_rbuf_f_rbuf_state_0_,
         U_rbuf_f_rbuf_state_1_, U_ctl_n422, U_ctl_n421, U_ctl_n420,
         U_ctl_n419, U_ctl_n418, U_ctl_n417, U_ctl_n416, U_ctl_n415,
         U_ctl_n414, U_ctl_n413, U_ctl_n412, U_ctl_n411, U_ctl_n410,
         U_ctl_n409, U_ctl_n408, U_ctl_n407, U_ctl_n406, U_ctl_n405,
         U_ctl_n404, U_ctl_n403, U_ctl_n402, U_ctl_n401, U_ctl_n400,
         U_ctl_n399, U_ctl_n398, U_ctl_n397, U_ctl_n396, U_ctl_n395,
         U_ctl_n394, U_ctl_n393, U_ctl_n392, U_ctl_n391, U_ctl_n390,
         U_ctl_n389, U_ctl_n388, U_ctl_n387, U_ctl_n386, U_ctl_n385,
         U_ctl_n384, U_ctl_n383, U_ctl_n382, U_ctl_n381, U_ctl_n380,
         U_ctl_n379, U_ctl_n378, U_ctl_n376, U_ctl_n375, U_ctl_n374,
         U_ctl_n373, U_ctl_n372, U_ctl_n371, U_ctl_n370, U_ctl_n369,
         U_ctl_n368, U_ctl_n367, U_ctl_n366, U_ctl_n365, U_ctl_n364,
         U_ctl_n363, U_ctl_n362, U_ctl_n361, U_ctl_n360, U_ctl_n359,
         U_ctl_n358, U_ctl_n357, U_ctl_n356, U_ctl_n355, U_ctl_n354,
         U_ctl_n353, U_ctl_n352, U_ctl_n351, U_ctl_n350, U_ctl_n349,
         U_ctl_n348, U_ctl_n347, U_ctl_n346, U_ctl_n345, U_ctl_n344,
         U_ctl_n343, U_ctl_n342, U_ctl_n341, U_ctl_n340, U_ctl_n339,
         U_ctl_n338, U_ctl_n337, U_ctl_n336, U_ctl_n335, U_ctl_n332,
         U_ctl_n331, U_ctl_n330, U_ctl_n329, U_ctl_n328, U_ctl_n327,
         U_ctl_n326, U_ctl_n325, U_ctl_n324, U_ctl_n323, U_ctl_n320,
         U_ctl_n319, U_ctl_n318, U_ctl_n317, U_ctl_n316, U_ctl_n315,
         U_ctl_n314, U_ctl_n313, U_ctl_n312, U_ctl_n311, U_ctl_n310,
         U_ctl_n309, U_ctl_n308, U_ctl_n307, U_ctl_n306, U_ctl_n305,
         U_ctl_n304, U_ctl_n303, U_ctl_n302, U_ctl_n301, U_ctl_n300,
         U_ctl_n298, U_ctl_n297, U_ctl_n296, U_ctl_n295, U_ctl_n294,
         U_ctl_n293, U_ctl_n292, U_ctl_n291, U_ctl_n290, U_ctl_n289,
         U_ctl_n288, U_ctl_n287, U_ctl_n286, U_ctl_n285, U_ctl_n284,
         U_ctl_n283, U_ctl_n282, U_ctl_n281, U_ctl_n280, U_ctl_n279,
         U_ctl_n278, U_ctl_n277, U_ctl_n276, U_ctl_n275, U_ctl_n274,
         U_ctl_n273, U_ctl_n272, U_ctl_n271, U_ctl_n270, U_ctl_n269,
         U_ctl_n268, U_ctl_n267, U_ctl_n266, U_ctl_n265, U_ctl_n264,
         U_ctl_n263, U_ctl_n262, U_ctl_n261, U_ctl_n260, U_ctl_n259,
         U_ctl_n258, U_ctl_n257, U_ctl_n256, U_ctl_n255, U_ctl_n254,
         U_ctl_n253, U_ctl_n252, U_ctl_n251, U_ctl_n250, U_ctl_n249,
         U_ctl_n248, U_ctl_n247, U_ctl_n246, U_ctl_n245, U_ctl_n244,
         U_ctl_n243, U_ctl_n242, U_ctl_n241, U_ctl_n238, U_ctl_n237,
         U_ctl_n236, U_ctl_n235, U_ctl_n234, U_ctl_n233, U_ctl_n232,
         U_ctl_n231, U_ctl_n230, U_ctl_n229, U_ctl_n228, U_ctl_n227,
         U_ctl_n226, U_ctl_n225, U_ctl_n224, U_ctl_n223, U_ctl_n222,
         U_ctl_n221, U_ctl_n220, U_ctl_n219, U_ctl_n218, U_ctl_n217,
         U_ctl_n216, U_ctl_n215, U_ctl_n214, U_ctl_n213, U_ctl_n212,
         U_ctl_n211, U_ctl_n210, U_ctl_n209, U_ctl_n208, U_ctl_n207,
         U_ctl_n206, U_ctl_n205, U_ctl_n204, U_ctl_n203, U_ctl_n202,
         U_ctl_n201, U_ctl_n200, U_ctl_n199, U_ctl_n198, U_ctl_n197,
         U_ctl_n196, U_ctl_n195, U_ctl_n194, U_ctl_n193, U_ctl_n190,
         U_ctl_n189, U_ctl_n188, U_ctl_n187, U_ctl_n186, U_ctl_n185,
         U_ctl_n184, U_ctl_n183, U_ctl_n182, U_ctl_n181, U_ctl_n180,
         U_ctl_n179, U_ctl_n178, U_ctl_n177, U_ctl_n176, U_ctl_n175,
         U_ctl_n174, U_ctl_n173, U_ctl_n172, U_ctl_n171, U_ctl_n170,
         U_ctl_n169, U_ctl_n168, U_ctl_n167, U_ctl_n166, U_ctl_n165,
         U_ctl_n164, U_ctl_n163, U_ctl_n161, U_ctl_n160, U_ctl_n159,
         U_ctl_n158, U_ctl_n157, U_ctl_n156, U_ctl_n155, U_ctl_n154,
         U_ctl_n153, U_ctl_n151, U_ctl_n150, U_ctl_n148, U_ctl_n147,
         U_ctl_n146, U_ctl_n145, U_ctl_n144, U_ctl_n143, U_ctl_n142,
         U_ctl_n126, U_ctl_n99, U_ctl_n98, U_ctl_n97, U_ctl_n96, U_ctl_n95,
         U_ctl_n94, U_ctl_n92, U_ctl_n91, U_ctl_n90, U_ctl_n89, U_ctl_n88,
         U_ctl_n87, U_ctl_n86, U_ctl_n85, U_ctl_n84, U_ctl_n83, U_ctl_n82,
         U_ctl_n81, U_ctl_n80, U_ctl_n79, U_ctl_n78, U_ctl_n77, U_ctl_n76,
         U_ctl_n75, U_ctl_n74, U_ctl_n73, U_ctl_n70, U_ctl_n69, U_ctl_n68,
         U_ctl_n67, U_ctl_n66, U_ctl_n65, U_ctl_n64, U_ctl_n63, U_ctl_n62,
         U_ctl_n61, U_ctl_n60, U_ctl_n59, U_ctl_n58, U_ctl_n57, U_ctl_n56,
         U_ctl_n55, U_ctl_n54, U_ctl_n53, U_ctl_n50, U_ctl_n47, U_ctl_n45,
         U_ctl_n44, U_ctl_n43, U_ctl_n42, U_ctl_n41, U_ctl_n40, U_ctl_n39,
         U_ctl_n38, U_ctl_n37, U_ctl_n36, U_ctl_n35, U_ctl_n34, U_ctl_n33,
         U_ctl_n32, U_ctl_n30, U_ctl_n29, U_ctl_n28, U_ctl_n26, U_ctl_n25,
         U_ctl_n24, U_ctl_n23, U_ctl_n22, U_ctl_n21, U_ctl_n20, U_ctl_n19,
         U_ctl_n18, U_ctl_n16, U_ctl_n15, U_ctl_n14, U_ctl_n13, U_ctl_n11,
         U_ctl_n10, U_ctl_n9, U_ctl_n8, U_ctl_n7, U_ctl_n6, U_ctl_n5, U_ctl_n3,
         U_ctl_DP_OP_140_125_8947_n1, U_ctl_DP_OP_140_125_8947_n2,
         U_ctl_DP_OP_140_125_8947_n3, U_ctl_DP_OP_140_125_8947_n4,
         U_ctl_DP_OP_140_125_8947_n5, U_ctl_DP_OP_140_125_8947_n6,
         U_ctl_DP_OP_140_125_8947_n7, U_ctl_DP_OP_140_125_8947_n8,
         U_ctl_DP_OP_140_125_8947_n9, U_ctl_DP_OP_140_125_8947_n10,
         U_ctl_DP_OP_140_125_8947_n11, U_ctl_DP_OP_140_125_8947_n12,
         U_ctl_DP_OP_140_125_8947_n13, U_ctl_DP_OP_140_125_8947_n14,
         U_ctl_DP_OP_140_125_8947_n15, U_ctl_DP_OP_140_125_8947_n16,
         U_ctl_DP_OP_140_125_8947_n17, U_ctl_DP_OP_140_125_8947_n18,
         U_ctl_DP_OP_140_125_8947_n19, U_ctl_DP_OP_140_125_8947_n20,
         U_ctl_DP_OP_140_125_8947_n22, U_ctl_DP_OP_140_125_8947_n23,
         U_ctl_DP_OP_140_125_8947_n24, U_ctl_DP_OP_140_125_8947_n30,
         U_ctl_DP_OP_140_125_8947_n31, U_ctl_DP_OP_140_125_8947_n32,
         U_ctl_DP_OP_140_125_8947_n33, U_ctl_DP_OP_140_125_8947_n34,
         U_ctl_DP_OP_140_125_8947_n35, U_ctl_DP_OP_140_125_8947_I2, U_ctl_n299,
         U_ctl_n141, U_ctl_n140, U_ctl_n139, U_ctl_n138, U_ctl_n137,
         U_ctl_n136, U_ctl_n135, U_ctl_n134, U_ctl_n133, U_ctl_n132,
         U_ctl_n131, U_ctl_n130, U_ctl_n129, U_ctl_n128, U_ctl_n127,
         U_ctl_n125, U_ctl_n124, U_ctl_n123, U_ctl_n122, U_ctl_n121,
         U_ctl_n120, U_ctl_n119, U_ctl_n118, U_ctl_n117, U_ctl_n116,
         U_ctl_n115, U_ctl_n114, U_ctl_n113, U_ctl_n112, U_ctl_n111,
         U_ctl_n110, U_ctl_n109, U_ctl_n108, U_ctl_n107, U_ctl_n106,
         U_ctl_n105, U_ctl_n104, U_ctl_n103, U_ctl_n102, U_ctl_n101,
         U_ctl_n100, U_ctl_C64_DATA2_5, U_ctl_C64_DATA2_0, U_ctl_f_burst_done,
         U_ctl_f_burst_done2, U_ctl_n_sel_buf, U_ctl_N288, U_ctl_N287,
         U_ctl_N286, U_ctl_N285, U_ctl_N284, U_ctl_f_hiu_terminate,
         U_ctl_fr_wr_bcnt_0_, U_ctl_fr_wr_bcnt_1_, U_ctl_fr_wr_bcnt_2_,
         U_ctl_fr_wr_bcnt_3_, U_ctl_fr_wr_bcnt_4_, U_ctl_fr_wr_bcnt_5_,
         U_ctl_N237, U_ctl_fr_prv_1wrap_tm, U_ctl_fr_prv_1wrap, U_ctl_N236,
         U_ctl_f_bh_state_0_, U_ctl_f_bh_state_1_, U_ctl_f_bh_state_2_,
         U_ctl_fd_rd_ready, U_ctl_fd_amba_bcnt_0_, U_ctl_fd_amba_bcnt_1_,
         U_ctl_fd_amba_bcnt_2_, U_ctl_fd_amba_bcnt_3_, U_ctl_N89,
         U_ctl_fd_rd_bz, U_ctl_fd_haddr_1_, U_ctl_fd_narrow_trans,
         U_ctl_fd_non_single, U_ctl_fd_incr, U_ctl_f_offset_0_,
         U_ctl_f_offset_1_, U_ctl_f_offset_2_, U_ctl_f_offset_3_,
         U_ctl_fd_wr_bz, U_ctl_fd_hsel_mem, U_ctl_fd_miu_data_width_0_,
         U_ctl_fd_miu_data_width_1_, U_ctl_fd_miu_col_width_0_,
         U_ctl_fd_miu_col_width_1_, U_ctl_fd_miu_col_width_2_,
         U_ctl_fd_miu_col_width_3_, U_ctl_f_data_width_0_, U_ctl_fd_wr_width,
         U_afifo_U_acore_n211, U_afifo_U_acore_n210, U_afifo_U_acore_n209,
         U_afifo_U_acore_n208, U_afifo_U_acore_n207, U_afifo_U_acore_n206,
         U_afifo_U_acore_n205, U_afifo_U_acore_n204, U_afifo_U_acore_n203,
         U_afifo_U_acore_n202, U_afifo_U_acore_n201, U_afifo_U_acore_n200,
         U_afifo_U_acore_n199, U_afifo_U_acore_n198, U_afifo_U_acore_n197,
         U_afifo_U_acore_n196, U_afifo_U_acore_n195, U_afifo_U_acore_n194,
         U_afifo_U_acore_n193, U_afifo_U_acore_n192, U_afifo_U_acore_n191,
         U_afifo_U_acore_n190, U_afifo_U_acore_n189, U_afifo_U_acore_n188,
         U_afifo_U_acore_n187, U_afifo_U_acore_n186, U_afifo_U_acore_n185,
         U_afifo_U_acore_n184, U_afifo_U_acore_n183, U_afifo_U_acore_n182,
         U_afifo_U_acore_n181, U_afifo_U_acore_n180, U_afifo_U_acore_n179,
         U_afifo_U_acore_n178, U_afifo_U_acore_n177, U_afifo_U_acore_n176,
         U_afifo_U_acore_n175, U_afifo_U_acore_n174, U_afifo_U_acore_n173,
         U_afifo_U_acore_n172, U_afifo_U_acore_n171, U_afifo_U_acore_n170,
         U_afifo_U_acore_n169, U_afifo_U_acore_n168, U_afifo_U_acore_n167,
         U_afifo_U_acore_n164, U_afifo_U_acore_n163, U_afifo_U_acore_n162,
         U_afifo_U_acore_n161, U_afifo_U_acore_n160, U_afifo_U_acore_n159,
         U_afifo_U_acore_n158, U_afifo_U_acore_n157, U_afifo_U_acore_n156,
         U_afifo_U_acore_n155, U_afifo_U_acore_n153, U_afifo_U_acore_n143,
         U_afifo_U_acore_n104, U_afifo_U_acore_n103, U_afifo_U_acore_n102,
         U_afifo_U_acore_n101, U_afifo_U_acore_n100, U_afifo_U_acore_n99,
         U_afifo_U_acore_n98, U_afifo_U_acore_n97, U_afifo_U_acore_n96,
         U_afifo_U_acore_n95, U_afifo_U_acore_n94, U_afifo_U_acore_n93,
         U_afifo_U_acore_n92, U_afifo_U_acore_n91, U_afifo_U_acore_n90,
         U_afifo_U_acore_n89, U_afifo_U_acore_n88, U_afifo_U_acore_n87,
         U_afifo_U_acore_n86, U_afifo_U_acore_n85, U_afifo_U_acore_n84,
         U_afifo_U_acore_n83, U_afifo_U_acore_n82, U_afifo_U_acore_n81,
         U_afifo_U_acore_n80, U_afifo_U_acore_n79, U_afifo_U_acore_n78,
         U_afifo_U_acore_n77, U_afifo_U_acore_n76, U_afifo_U_acore_n75,
         U_afifo_U_acore_n74, U_afifo_U_acore_n73, U_afifo_U_acore_n72,
         U_afifo_U_acore_n71, U_afifo_U_acore_n70, U_afifo_U_acore_n69,
         U_afifo_U_acore_n68, U_afifo_U_acore_n67, U_afifo_U_acore_n66,
         U_afifo_U_acore_n65, U_afifo_U_acore_n64, U_afifo_U_acore_n63,
         U_afifo_U_acore_n62, U_afifo_U_acore_n61, U_afifo_U_acore_n60,
         U_afifo_U_acore_n59, U_afifo_U_acore_n58, U_afifo_U_acore_n57,
         U_afifo_U_acore_n56, U_afifo_U_acore_n55, U_afifo_U_acore_n54,
         U_afifo_U_acore_n53, U_afifo_U_acore_n51, U_afifo_U_acore_n49,
         U_afifo_U_acore_n48, U_afifo_U_acore_n47, U_afifo_U_acore_n46,
         U_afifo_U_acore_n45, U_afifo_U_acore_n44, U_afifo_U_acore_n43,
         U_afifo_U_acore_n42, U_afifo_U_acore_n41, U_afifo_U_acore_n40,
         U_afifo_U_acore_n39, U_afifo_U_acore_n38, U_afifo_U_acore_n37,
         U_afifo_U_acore_n36, U_afifo_U_acore_n35, U_afifo_U_acore_n34,
         U_afifo_U_acore_n33, U_afifo_U_acore_n32, U_afifo_U_acore_n31,
         U_afifo_U_acore_n30, U_afifo_U_acore_n29, U_afifo_U_acore_n28,
         U_afifo_U_acore_n27, U_afifo_U_acore_n26, U_afifo_U_acore_n25,
         U_afifo_U_acore_n24, U_afifo_U_acore_n23, U_afifo_U_acore_n22,
         U_afifo_U_acore_n21, U_afifo_U_acore_n20, U_afifo_U_acore_n19,
         U_afifo_U_acore_n18, U_afifo_U_acore_n17, U_afifo_U_acore_n16,
         U_afifo_U_acore_n15, U_afifo_U_acore_n14, U_afifo_U_acore_n13,
         U_afifo_U_acore_n12, U_afifo_U_acore_n11, U_afifo_U_acore_n10,
         U_afifo_U_acore_n9, U_afifo_U_acore_n8, U_afifo_U_acore_n7,
         U_afifo_U_acore_n6, U_afifo_U_acore_n5, U_afifo_U_acore_n4,
         U_afifo_U_acore_n3, U_afifo_U_acore_n2, U_afifo_U_acore_n1,
         U_afifo_U_acore_n166, U_afifo_U_acore_n165, U_afifo_U_acore_n154,
         U_afifo_U_acore_n152, U_afifo_U_acore_n151, U_afifo_U_acore_n150,
         U_afifo_U_acore_n149, U_afifo_U_acore_n148, U_afifo_U_acore_n147,
         U_afifo_U_acore_n146, U_afifo_U_acore_n145, U_afifo_U_acore_n144,
         U_afifo_U_acore_n142, U_afifo_U_acore_n141, U_afifo_U_acore_n140,
         U_afifo_U_acore_n139, U_afifo_U_acore_n138, U_afifo_U_acore_n137,
         U_afifo_U_acore_n136, U_afifo_U_acore_n135, U_afifo_U_acore_n134,
         U_afifo_U_acore_n133, U_afifo_U_acore_n132, U_afifo_U_acore_n131,
         U_afifo_U_acore_n130, U_afifo_U_acore_n129, U_afifo_U_acore_n128,
         U_afifo_U_acore_n127, U_afifo_U_acore_n126, U_afifo_U_acore_n125,
         U_afifo_U_acore_n124, U_afifo_U_acore_n123, U_afifo_U_acore_n122,
         U_afifo_U_acore_n121, U_afifo_U_acore_n120, U_afifo_U_acore_n119,
         U_afifo_U_acore_n118, U_afifo_U_acore_n117, U_afifo_U_acore_n116,
         U_afifo_U_acore_n115, U_afifo_U_acore_n114, U_afifo_U_acore_n113,
         U_afifo_U_acore_n112, U_afifo_U_acore_n111, U_afifo_U_acore_n110,
         U_afifo_U_acore_n109, U_afifo_U_acore_n108, U_afifo_U_acore_n107,
         U_afifo_U_acore_n106, U_afifo_U_acore_n105, U_afifo_U_acore_n_afull,
         U_afifo_U_acore_f_afull, U_afifo_U_acore_n_obuf_empty,
         U_afifo_U_acore_f_obuf_0_, U_afifo_U_acore_f_obuf_2_,
         U_afifo_U_acore_f_obuf_3_, U_afifo_U_acore_f_obuf_4_,
         U_afifo_U_acore_f_obuf_5_, U_afifo_U_acore_f_obuf_6_,
         U_afifo_U_acore_f_obuf_7_, U_afifo_U_acore_f_obuf_8_,
         U_afifo_U_acore_f_obuf_9_, U_afifo_U_acore_f_obuf_11_,
         U_afifo_U_acore_f_obuf_12_, U_afifo_U_acore_f_obuf_13_,
         U_afifo_U_acore_f_obuf_14_, U_afifo_U_acore_f_obuf_15_,
         U_afifo_U_acore_f_obuf_16_, U_afifo_U_acore_f_obuf_17_,
         U_afifo_U_acore_f_obuf_18_, U_afifo_U_acore_f_obuf_19_,
         U_afifo_U_acore_f_obuf_20_, U_afifo_U_acore_f_obuf_21_,
         U_afifo_U_acore_f_obuf_22_, U_afifo_U_acore_f_obuf_23_,
         U_afifo_U_acore_f_obuf_24_, U_afifo_U_acore_f_obuf_25_,
         U_afifo_U_acore_f_obuf_26_, U_afifo_U_acore_f_obuf_27_,
         U_afifo_U_acore_f_obuf_28_, U_afifo_U_acore_f_obuf_29_,
         U_afifo_U_acore_f_obuf_30_, U_afifo_U_acore_f_obuf_31_,
         U_afifo_U_acore_f_obuf_32_, U_afifo_U_acore_f_obuf_33_,
         U_afifo_U_acore_f_obuf_34_, U_afifo_U_acore_f_obuf_35_,
         U_afifo_U_acore_f_obuf_36_, U_afifo_U_acore_f_obuf_37_,
         U_afifo_U_acore_f_obuf_38_, U_afifo_U_acore_f_obuf_39_,
         U_afifo_U_acore_f_obuf_40_, U_afifo_U_acore_f_obuf_41_,
         U_afifo_U_acore_f_obuf_42_, U_afifo_U_acore_f_obuf_43_,
         U_afifo_U_acore_f_obuf_44_, U_afifo_U_acore_f_obuf_45_,
         U_afifo_U_acore_f_obuf_46_, U_afifo_U_acore_f_obuf_47_,
         U_afifo_U_acore_f_obuf_48_, U_afifo_U_acore_f_obuf_49_,
         U_afifo_U_acore_f_push_req_n, U_afifo_U_acore_m_sf_full,
         U_afifo_U_acore_f_ibuf_2_, U_afifo_U_acore_f_ibuf_18_,
         U_afifo_U_acore_f_ibuf_30_, U_afifo_U_acore_f_ibuf_31_,
         U_afifo_U_acore_f_ibuf_32_, U_afifo_U_acore_f_ibuf_33_,
         U_afifo_U_acore_f_ibuf_34_, U_afifo_U_acore_f_ibuf_35_,
         U_afifo_U_acore_f_ibuf_36_, U_afifo_U_acore_f_ibuf_37_,
         U_afifo_U_acore_f_ibuf_38_, U_afifo_U_acore_f_ibuf_39_,
         U_afifo_U_acore_f_ibuf_40_, U_afifo_U_acore_f_ibuf_41_,
         U_dfifo_U_dcore_n234, U_dfifo_U_dcore_n233, U_dfifo_U_dcore_n232,
         U_dfifo_U_dcore_n231, U_dfifo_U_dcore_n230, U_dfifo_U_dcore_n229,
         U_dfifo_U_dcore_n228, U_dfifo_U_dcore_n227, U_dfifo_U_dcore_n226,
         U_dfifo_U_dcore_n225, U_dfifo_U_dcore_n224, U_dfifo_U_dcore_n223,
         U_dfifo_U_dcore_n222, U_dfifo_U_dcore_n221, U_dfifo_U_dcore_n220,
         U_dfifo_U_dcore_n219, U_dfifo_U_dcore_n218, U_dfifo_U_dcore_n217,
         U_dfifo_U_dcore_n216, U_dfifo_U_dcore_n215, U_dfifo_U_dcore_n214,
         U_dfifo_U_dcore_n213, U_dfifo_U_dcore_n212, U_dfifo_U_dcore_n211,
         U_dfifo_U_dcore_n210, U_dfifo_U_dcore_n207, U_dfifo_U_dcore_n206,
         U_dfifo_U_dcore_n205, U_dfifo_U_dcore_n204, U_dfifo_U_dcore_n202,
         U_dfifo_U_dcore_n133, U_dfifo_U_dcore_n132, U_dfifo_U_dcore_n131,
         U_dfifo_U_dcore_n130, U_dfifo_U_dcore_n129, U_dfifo_U_dcore_n128,
         U_dfifo_U_dcore_n127, U_dfifo_U_dcore_n126, U_dfifo_U_dcore_n125,
         U_dfifo_U_dcore_n124, U_dfifo_U_dcore_n123, U_dfifo_U_dcore_n122,
         U_dfifo_U_dcore_n121, U_dfifo_U_dcore_n120, U_dfifo_U_dcore_n119,
         U_dfifo_U_dcore_n118, U_dfifo_U_dcore_n117, U_dfifo_U_dcore_n116,
         U_dfifo_U_dcore_n115, U_dfifo_U_dcore_n114, U_dfifo_U_dcore_n113,
         U_dfifo_U_dcore_n112, U_dfifo_U_dcore_n111, U_dfifo_U_dcore_n110,
         U_dfifo_U_dcore_n109, U_dfifo_U_dcore_n108, U_dfifo_U_dcore_n107,
         U_dfifo_U_dcore_n106, U_dfifo_U_dcore_n105, U_dfifo_U_dcore_n104,
         U_dfifo_U_dcore_n103, U_dfifo_U_dcore_n102, U_dfifo_U_dcore_n101,
         U_dfifo_U_dcore_n100, U_dfifo_U_dcore_n99, U_dfifo_U_dcore_n98,
         U_dfifo_U_dcore_n97, U_dfifo_U_dcore_n96, U_dfifo_U_dcore_n95,
         U_dfifo_U_dcore_n94, U_dfifo_U_dcore_n93, U_dfifo_U_dcore_n92,
         U_dfifo_U_dcore_n91, U_dfifo_U_dcore_n90, U_dfifo_U_dcore_n89,
         U_dfifo_U_dcore_n88, U_dfifo_U_dcore_n87, U_dfifo_U_dcore_n86,
         U_dfifo_U_dcore_n85, U_dfifo_U_dcore_n84, U_dfifo_U_dcore_n83,
         U_dfifo_U_dcore_n82, U_dfifo_U_dcore_n81, U_dfifo_U_dcore_n80,
         U_dfifo_U_dcore_n79, U_dfifo_U_dcore_n78, U_dfifo_U_dcore_n77,
         U_dfifo_U_dcore_n76, U_dfifo_U_dcore_n75, U_dfifo_U_dcore_n74,
         U_dfifo_U_dcore_n73, U_dfifo_U_dcore_n72, U_dfifo_U_dcore_n71,
         U_dfifo_U_dcore_n70, U_dfifo_U_dcore_n69, U_dfifo_U_dcore_n68,
         U_dfifo_U_dcore_n67, U_dfifo_U_dcore_n66, U_dfifo_U_dcore_n65,
         U_dfifo_U_dcore_n64, U_dfifo_U_dcore_n63, U_dfifo_U_dcore_n62,
         U_dfifo_U_dcore_n61, U_dfifo_U_dcore_n60, U_dfifo_U_dcore_n59,
         U_dfifo_U_dcore_n58, U_dfifo_U_dcore_n57, U_dfifo_U_dcore_n56,
         U_dfifo_U_dcore_n55, U_dfifo_U_dcore_n54, U_dfifo_U_dcore_n53,
         U_dfifo_U_dcore_n52, U_dfifo_U_dcore_n51, U_dfifo_U_dcore_n50,
         U_dfifo_U_dcore_n49, U_dfifo_U_dcore_n48, U_dfifo_U_dcore_n47,
         U_dfifo_U_dcore_n46, U_dfifo_U_dcore_n45, U_dfifo_U_dcore_n44,
         U_dfifo_U_dcore_n43, U_dfifo_U_dcore_n42, U_dfifo_U_dcore_n41,
         U_dfifo_U_dcore_n40, U_dfifo_U_dcore_n39, U_dfifo_U_dcore_n38,
         U_dfifo_U_dcore_n37, U_dfifo_U_dcore_n36, U_dfifo_U_dcore_n35,
         U_dfifo_U_dcore_n34, U_dfifo_U_dcore_n33, U_dfifo_U_dcore_n32,
         U_dfifo_U_dcore_n31, U_dfifo_U_dcore_n30, U_dfifo_U_dcore_n29,
         U_dfifo_U_dcore_n28, U_dfifo_U_dcore_n27, U_dfifo_U_dcore_n26,
         U_dfifo_U_dcore_n25, U_dfifo_U_dcore_n24, U_dfifo_U_dcore_n23,
         U_dfifo_U_dcore_n22, U_dfifo_U_dcore_n21, U_dfifo_U_dcore_n20,
         U_dfifo_U_dcore_n19, U_dfifo_U_dcore_n18, U_dfifo_U_dcore_n17,
         U_dfifo_U_dcore_n16, U_dfifo_U_dcore_n15, U_dfifo_U_dcore_n14,
         U_dfifo_U_dcore_n13, U_dfifo_U_dcore_n12, U_dfifo_U_dcore_n11,
         U_dfifo_U_dcore_n10, U_dfifo_U_dcore_n9, U_dfifo_U_dcore_n8,
         U_dfifo_U_dcore_n7, U_dfifo_U_dcore_n6, U_dfifo_U_dcore_n5,
         U_dfifo_U_dcore_n4, U_dfifo_U_dcore_n3, U_dfifo_U_dcore_n2,
         U_dfifo_U_dcore_n1, U_dfifo_U_dcore_n209, U_dfifo_U_dcore_n208,
         U_dfifo_U_dcore_n203, U_dfifo_U_dcore_n201, U_dfifo_U_dcore_n200,
         U_dfifo_U_dcore_n199, U_dfifo_U_dcore_n198, U_dfifo_U_dcore_n197,
         U_dfifo_U_dcore_n196, U_dfifo_U_dcore_n195, U_dfifo_U_dcore_n194,
         U_dfifo_U_dcore_n193, U_dfifo_U_dcore_n192, U_dfifo_U_dcore_n191,
         U_dfifo_U_dcore_n190, U_dfifo_U_dcore_n189, U_dfifo_U_dcore_n188,
         U_dfifo_U_dcore_n187, U_dfifo_U_dcore_n186, U_dfifo_U_dcore_n185,
         U_dfifo_U_dcore_n184, U_dfifo_U_dcore_n183, U_dfifo_U_dcore_n182,
         U_dfifo_U_dcore_n181, U_dfifo_U_dcore_n180, U_dfifo_U_dcore_n179,
         U_dfifo_U_dcore_n178, U_dfifo_U_dcore_n177, U_dfifo_U_dcore_n176,
         U_dfifo_U_dcore_n175, U_dfifo_U_dcore_n174, U_dfifo_U_dcore_n173,
         U_dfifo_U_dcore_n172, U_dfifo_U_dcore_n171, U_dfifo_U_dcore_n170,
         U_dfifo_U_dcore_n169, U_dfifo_U_dcore_n168, U_dfifo_U_dcore_n167,
         U_dfifo_U_dcore_n166, U_dfifo_U_dcore_n165, U_dfifo_U_dcore_n164,
         U_dfifo_U_dcore_n163, U_dfifo_U_dcore_n162, U_dfifo_U_dcore_n161,
         U_dfifo_U_dcore_n160, U_dfifo_U_dcore_n159, U_dfifo_U_dcore_n158,
         U_dfifo_U_dcore_n157, U_dfifo_U_dcore_n156, U_dfifo_U_dcore_n155,
         U_dfifo_U_dcore_n154, U_dfifo_U_dcore_n153, U_dfifo_U_dcore_n152,
         U_dfifo_U_dcore_n151, U_dfifo_U_dcore_n150, U_dfifo_U_dcore_n149,
         U_dfifo_U_dcore_n148, U_dfifo_U_dcore_n147, U_dfifo_U_dcore_n146,
         U_dfifo_U_dcore_n145, U_dfifo_U_dcore_n144, U_dfifo_U_dcore_n143,
         U_dfifo_U_dcore_n142, U_dfifo_U_dcore_n141, U_dfifo_U_dcore_n140,
         U_dfifo_U_dcore_n139, U_dfifo_U_dcore_n138, U_dfifo_U_dcore_n137,
         U_dfifo_U_dcore_n136, U_dfifo_U_dcore_n135, U_dfifo_U_dcore_n134,
         U_dfifo_U_dcore_n_empty, U_dfifo_U_dcore_f_buf_has_data,
         U_dfifo_U_dcore_m_sf_full, U_dfifo_U_dcore_m_sf_afull,
         U_dfifo_U_dcore_m_sf_empty, U_dfifo_U_dcore_f_buf_data_0_,
         U_dfifo_U_dcore_f_buf_data_1_, U_dfifo_U_dcore_f_buf_data_2_,
         U_dfifo_U_dcore_f_buf_data_3_, U_dfifo_U_dcore_f_buf_data_4_,
         U_dfifo_U_dcore_f_buf_data_5_, U_dfifo_U_dcore_f_buf_data_6_,
         U_dfifo_U_dcore_f_buf_data_7_, U_dfifo_U_dcore_f_buf_data_8_,
         U_dfifo_U_dcore_f_buf_data_9_, U_dfifo_U_dcore_f_buf_data_10_,
         U_dfifo_U_dcore_f_buf_data_11_, U_dfifo_U_dcore_f_buf_data_12_,
         U_dfifo_U_dcore_f_buf_data_13_, U_dfifo_U_dcore_f_buf_data_14_,
         U_dfifo_U_dcore_f_buf_data_15_, U_dfifo_U_dcore_f_buf_data_16_,
         U_dfifo_U_dcore_f_buf_data_17_, U_dfifo_U_dcore_f_buf_data_18_,
         U_dfifo_U_dcore_f_buf_data_19_, U_dfifo_U_dcore_f_buf_data_20_,
         U_dfifo_U_dcore_f_buf_data_21_, U_dfifo_U_dcore_f_buf_data_22_,
         U_dfifo_U_dcore_f_buf_data_23_, U_dfifo_U_dcore_f_buf_data_24_,
         U_dfifo_U_dcore_f_buf_data_25_, U_dfifo_U_dcore_f_buf_data_26_,
         U_dfifo_U_dcore_f_buf_data_27_, U_dfifo_U_dcore_f_buf_data_28_,
         U_dfifo_U_dcore_f_buf_data_29_, U_dfifo_U_dcore_f_buf_data_30_,
         U_dfifo_U_dcore_f_buf_data_31_, U_dfifo_U_dcore_f_buf_data_32_,
         U_dfifo_U_dcore_f_buf_data_33_, U_afifo_U_acore_U_sub_fifo_n373,
         U_afifo_U_acore_U_sub_fifo_n372, U_afifo_U_acore_U_sub_fifo_n371,
         U_afifo_U_acore_U_sub_fifo_n370, U_afifo_U_acore_U_sub_fifo_n369,
         U_afifo_U_acore_U_sub_fifo_n212, U_afifo_U_acore_U_sub_fifo_n169,
         U_afifo_U_acore_U_sub_fifo_n168, U_afifo_U_acore_U_sub_fifo_n167,
         U_afifo_U_acore_U_sub_fifo_n166, U_afifo_U_acore_U_sub_fifo_n165,
         U_afifo_U_acore_U_sub_fifo_n163, U_afifo_U_acore_U_sub_fifo_n162,
         U_afifo_U_acore_U_sub_fifo_n161, U_afifo_U_acore_U_sub_fifo_n160,
         U_afifo_U_acore_U_sub_fifo_n159, U_afifo_U_acore_U_sub_fifo_n158,
         U_afifo_U_acore_U_sub_fifo_n153, U_afifo_U_acore_U_sub_fifo_n152,
         U_afifo_U_acore_U_sub_fifo_n151, U_afifo_U_acore_U_sub_fifo_n150,
         U_afifo_U_acore_U_sub_fifo_n149, U_afifo_U_acore_U_sub_fifo_n148,
         U_afifo_U_acore_U_sub_fifo_n147, U_afifo_U_acore_U_sub_fifo_n146,
         U_afifo_U_acore_U_sub_fifo_n145, U_afifo_U_acore_U_sub_fifo_n144,
         U_afifo_U_acore_U_sub_fifo_n143, U_afifo_U_acore_U_sub_fifo_n142,
         U_afifo_U_acore_U_sub_fifo_n141, U_afifo_U_acore_U_sub_fifo_n140,
         U_afifo_U_acore_U_sub_fifo_n139, U_afifo_U_acore_U_sub_fifo_n138,
         U_afifo_U_acore_U_sub_fifo_n137, U_afifo_U_acore_U_sub_fifo_n136,
         U_afifo_U_acore_U_sub_fifo_n135, U_afifo_U_acore_U_sub_fifo_n134,
         U_afifo_U_acore_U_sub_fifo_n133, U_afifo_U_acore_U_sub_fifo_n132,
         U_afifo_U_acore_U_sub_fifo_n131, U_afifo_U_acore_U_sub_fifo_n130,
         U_afifo_U_acore_U_sub_fifo_n129, U_afifo_U_acore_U_sub_fifo_n128,
         U_afifo_U_acore_U_sub_fifo_n127, U_afifo_U_acore_U_sub_fifo_n126,
         U_afifo_U_acore_U_sub_fifo_n125, U_afifo_U_acore_U_sub_fifo_n124,
         U_afifo_U_acore_U_sub_fifo_n123, U_afifo_U_acore_U_sub_fifo_n122,
         U_afifo_U_acore_U_sub_fifo_n121, U_afifo_U_acore_U_sub_fifo_n120,
         U_afifo_U_acore_U_sub_fifo_n119, U_afifo_U_acore_U_sub_fifo_n118,
         U_afifo_U_acore_U_sub_fifo_n117, U_afifo_U_acore_U_sub_fifo_n116,
         U_afifo_U_acore_U_sub_fifo_n115, U_afifo_U_acore_U_sub_fifo_n114,
         U_afifo_U_acore_U_sub_fifo_n113, U_afifo_U_acore_U_sub_fifo_n112,
         U_afifo_U_acore_U_sub_fifo_n111, U_afifo_U_acore_U_sub_fifo_n110,
         U_afifo_U_acore_U_sub_fifo_n109, U_afifo_U_acore_U_sub_fifo_n108,
         U_afifo_U_acore_U_sub_fifo_n107, U_afifo_U_acore_U_sub_fifo_n106,
         U_afifo_U_acore_U_sub_fifo_n105, U_afifo_U_acore_U_sub_fifo_n104,
         U_afifo_U_acore_U_sub_fifo_n103, U_afifo_U_acore_U_sub_fifo_n102,
         U_afifo_U_acore_U_sub_fifo_n101, U_afifo_U_acore_U_sub_fifo_n100,
         U_afifo_U_acore_U_sub_fifo_n99, U_afifo_U_acore_U_sub_fifo_n98,
         U_afifo_U_acore_U_sub_fifo_n97, U_afifo_U_acore_U_sub_fifo_n96,
         U_afifo_U_acore_U_sub_fifo_n95, U_afifo_U_acore_U_sub_fifo_n94,
         U_afifo_U_acore_U_sub_fifo_n93, U_afifo_U_acore_U_sub_fifo_n92,
         U_afifo_U_acore_U_sub_fifo_n91, U_afifo_U_acore_U_sub_fifo_n90,
         U_afifo_U_acore_U_sub_fifo_n89, U_afifo_U_acore_U_sub_fifo_n88,
         U_afifo_U_acore_U_sub_fifo_n87, U_afifo_U_acore_U_sub_fifo_n86,
         U_afifo_U_acore_U_sub_fifo_n85, U_afifo_U_acore_U_sub_fifo_n84,
         U_afifo_U_acore_U_sub_fifo_n83, U_afifo_U_acore_U_sub_fifo_n82,
         U_afifo_U_acore_U_sub_fifo_n81, U_afifo_U_acore_U_sub_fifo_n80,
         U_afifo_U_acore_U_sub_fifo_n79, U_afifo_U_acore_U_sub_fifo_n78,
         U_afifo_U_acore_U_sub_fifo_n77, U_afifo_U_acore_U_sub_fifo_n76,
         U_afifo_U_acore_U_sub_fifo_n75, U_afifo_U_acore_U_sub_fifo_n74,
         U_afifo_U_acore_U_sub_fifo_n73, U_afifo_U_acore_U_sub_fifo_n72,
         U_afifo_U_acore_U_sub_fifo_n71, U_afifo_U_acore_U_sub_fifo_n70,
         U_afifo_U_acore_U_sub_fifo_n69, U_afifo_U_acore_U_sub_fifo_n68,
         U_afifo_U_acore_U_sub_fifo_n67, U_afifo_U_acore_U_sub_fifo_n66,
         U_afifo_U_acore_U_sub_fifo_n65, U_afifo_U_acore_U_sub_fifo_n64,
         U_afifo_U_acore_U_sub_fifo_n63, U_afifo_U_acore_U_sub_fifo_n62,
         U_afifo_U_acore_U_sub_fifo_n61, U_afifo_U_acore_U_sub_fifo_n60,
         U_afifo_U_acore_U_sub_fifo_n59, U_afifo_U_acore_U_sub_fifo_n58,
         U_afifo_U_acore_U_sub_fifo_n57, U_afifo_U_acore_U_sub_fifo_n56,
         U_afifo_U_acore_U_sub_fifo_n55, U_afifo_U_acore_U_sub_fifo_n54,
         U_afifo_U_acore_U_sub_fifo_n53, U_afifo_U_acore_U_sub_fifo_n52,
         U_afifo_U_acore_U_sub_fifo_n51, U_afifo_U_acore_U_sub_fifo_n50,
         U_afifo_U_acore_U_sub_fifo_n49, U_afifo_U_acore_U_sub_fifo_n48,
         U_afifo_U_acore_U_sub_fifo_n47, U_afifo_U_acore_U_sub_fifo_n46,
         U_afifo_U_acore_U_sub_fifo_n45, U_afifo_U_acore_U_sub_fifo_n44,
         U_afifo_U_acore_U_sub_fifo_n43, U_afifo_U_acore_U_sub_fifo_n42,
         U_afifo_U_acore_U_sub_fifo_n41, U_afifo_U_acore_U_sub_fifo_n40,
         U_afifo_U_acore_U_sub_fifo_n39, U_afifo_U_acore_U_sub_fifo_n38,
         U_afifo_U_acore_U_sub_fifo_n37, U_afifo_U_acore_U_sub_fifo_n36,
         U_afifo_U_acore_U_sub_fifo_n35, U_afifo_U_acore_U_sub_fifo_n34,
         U_afifo_U_acore_U_sub_fifo_n33, U_afifo_U_acore_U_sub_fifo_n32,
         U_afifo_U_acore_U_sub_fifo_n31, U_afifo_U_acore_U_sub_fifo_n30,
         U_afifo_U_acore_U_sub_fifo_n29, U_afifo_U_acore_U_sub_fifo_n28,
         U_afifo_U_acore_U_sub_fifo_n27, U_afifo_U_acore_U_sub_fifo_n26,
         U_afifo_U_acore_U_sub_fifo_n25, U_afifo_U_acore_U_sub_fifo_n24,
         U_afifo_U_acore_U_sub_fifo_n23, U_afifo_U_acore_U_sub_fifo_n22,
         U_afifo_U_acore_U_sub_fifo_n21, U_afifo_U_acore_U_sub_fifo_n20,
         U_afifo_U_acore_U_sub_fifo_n19, U_afifo_U_acore_U_sub_fifo_n18,
         U_afifo_U_acore_U_sub_fifo_n17, U_afifo_U_acore_U_sub_fifo_n16,
         U_afifo_U_acore_U_sub_fifo_n15, U_afifo_U_acore_U_sub_fifo_n14,
         U_afifo_U_acore_U_sub_fifo_n13, U_afifo_U_acore_U_sub_fifo_n12,
         U_afifo_U_acore_U_sub_fifo_n11, U_afifo_U_acore_U_sub_fifo_n10,
         U_afifo_U_acore_U_sub_fifo_n9, U_afifo_U_acore_U_sub_fifo_n8,
         U_afifo_U_acore_U_sub_fifo_n7, U_afifo_U_acore_U_sub_fifo_n6,
         U_afifo_U_acore_U_sub_fifo_n5, U_afifo_U_acore_U_sub_fifo_n4,
         U_afifo_U_acore_U_sub_fifo_n3, U_afifo_U_acore_U_sub_fifo_n2,
         U_afifo_U_acore_U_sub_fifo_n1, U_afifo_U_acore_U_sub_fifo_n325,
         U_afifo_U_acore_U_sub_fifo_n324, U_afifo_U_acore_U_sub_fifo_n323,
         U_afifo_U_acore_U_sub_fifo_n322, U_afifo_U_acore_U_sub_fifo_n320,
         U_afifo_U_acore_U_sub_fifo_n319, U_afifo_U_acore_U_sub_fifo_n318,
         U_afifo_U_acore_U_sub_fifo_n317, U_afifo_U_acore_U_sub_fifo_n316,
         U_afifo_U_acore_U_sub_fifo_n315, U_afifo_U_acore_U_sub_fifo_n314,
         U_afifo_U_acore_U_sub_fifo_n313, U_afifo_U_acore_U_sub_fifo_n311,
         U_afifo_U_acore_U_sub_fifo_n310, U_afifo_U_acore_U_sub_fifo_n309,
         U_afifo_U_acore_U_sub_fifo_n308, U_afifo_U_acore_U_sub_fifo_n307,
         U_afifo_U_acore_U_sub_fifo_n306, U_afifo_U_acore_U_sub_fifo_n305,
         U_afifo_U_acore_U_sub_fifo_n304, U_afifo_U_acore_U_sub_fifo_n303,
         U_afifo_U_acore_U_sub_fifo_n302, U_afifo_U_acore_U_sub_fifo_n301,
         U_afifo_U_acore_U_sub_fifo_n300, U_afifo_U_acore_U_sub_fifo_n299,
         U_afifo_U_acore_U_sub_fifo_n298, U_afifo_U_acore_U_sub_fifo_n297,
         U_afifo_U_acore_U_sub_fifo_n296, U_afifo_U_acore_U_sub_fifo_n295,
         U_afifo_U_acore_U_sub_fifo_n294, U_afifo_U_acore_U_sub_fifo_n293,
         U_afifo_U_acore_U_sub_fifo_n292, U_afifo_U_acore_U_sub_fifo_n291,
         U_afifo_U_acore_U_sub_fifo_n290, U_afifo_U_acore_U_sub_fifo_n289,
         U_afifo_U_acore_U_sub_fifo_n288, U_afifo_U_acore_U_sub_fifo_n287,
         U_afifo_U_acore_U_sub_fifo_n286, U_afifo_U_acore_U_sub_fifo_n285,
         U_afifo_U_acore_U_sub_fifo_n284, U_afifo_U_acore_U_sub_fifo_n283,
         U_afifo_U_acore_U_sub_fifo_n282, U_afifo_U_acore_U_sub_fifo_n281,
         U_afifo_U_acore_U_sub_fifo_n280, U_afifo_U_acore_U_sub_fifo_n279,
         U_afifo_U_acore_U_sub_fifo_n278, U_afifo_U_acore_U_sub_fifo_n277,
         U_afifo_U_acore_U_sub_fifo_n276, U_afifo_U_acore_U_sub_fifo_n275,
         U_afifo_U_acore_U_sub_fifo_n274, U_afifo_U_acore_U_sub_fifo_n273,
         U_afifo_U_acore_U_sub_fifo_n272, U_afifo_U_acore_U_sub_fifo_n270,
         U_afifo_U_acore_U_sub_fifo_n269, U_afifo_U_acore_U_sub_fifo_n268,
         U_afifo_U_acore_U_sub_fifo_n267, U_afifo_U_acore_U_sub_fifo_n266,
         U_afifo_U_acore_U_sub_fifo_n265, U_afifo_U_acore_U_sub_fifo_n264,
         U_afifo_U_acore_U_sub_fifo_n263, U_afifo_U_acore_U_sub_fifo_n261,
         U_afifo_U_acore_U_sub_fifo_n260, U_afifo_U_acore_U_sub_fifo_n259,
         U_afifo_U_acore_U_sub_fifo_n258, U_afifo_U_acore_U_sub_fifo_n257,
         U_afifo_U_acore_U_sub_fifo_n256, U_afifo_U_acore_U_sub_fifo_n255,
         U_afifo_U_acore_U_sub_fifo_n254, U_afifo_U_acore_U_sub_fifo_n253,
         U_afifo_U_acore_U_sub_fifo_n252, U_afifo_U_acore_U_sub_fifo_n251,
         U_afifo_U_acore_U_sub_fifo_n250, U_afifo_U_acore_U_sub_fifo_n249,
         U_afifo_U_acore_U_sub_fifo_n248, U_afifo_U_acore_U_sub_fifo_n247,
         U_afifo_U_acore_U_sub_fifo_n246, U_afifo_U_acore_U_sub_fifo_n245,
         U_afifo_U_acore_U_sub_fifo_n244, U_afifo_U_acore_U_sub_fifo_n243,
         U_afifo_U_acore_U_sub_fifo_n242, U_afifo_U_acore_U_sub_fifo_n241,
         U_afifo_U_acore_U_sub_fifo_n240, U_afifo_U_acore_U_sub_fifo_n239,
         U_afifo_U_acore_U_sub_fifo_n238, U_afifo_U_acore_U_sub_fifo_n237,
         U_afifo_U_acore_U_sub_fifo_n236, U_afifo_U_acore_U_sub_fifo_n235,
         U_afifo_U_acore_U_sub_fifo_n234, U_afifo_U_acore_U_sub_fifo_n233,
         U_afifo_U_acore_U_sub_fifo_n232, U_afifo_U_acore_U_sub_fifo_n231,
         U_afifo_U_acore_U_sub_fifo_n230, U_afifo_U_acore_U_sub_fifo_n229,
         U_afifo_U_acore_U_sub_fifo_n228, U_afifo_U_acore_U_sub_fifo_n227,
         U_afifo_U_acore_U_sub_fifo_n226, U_afifo_U_acore_U_sub_fifo_n225,
         U_afifo_U_acore_U_sub_fifo_n224, U_afifo_U_acore_U_sub_fifo_n223,
         U_afifo_U_acore_U_sub_fifo_n222, U_afifo_U_acore_U_sub_fifo_n220,
         U_afifo_U_acore_U_sub_fifo_n219, U_afifo_U_acore_U_sub_fifo_n218,
         U_afifo_U_acore_U_sub_fifo_n217, U_afifo_U_acore_U_sub_fifo_n216,
         U_afifo_U_acore_U_sub_fifo_n215, U_afifo_U_acore_U_sub_fifo_n214,
         U_afifo_U_acore_U_sub_fifo_n213, U_afifo_U_acore_U_sub_fifo_n211,
         U_afifo_U_acore_U_sub_fifo_n210, U_afifo_U_acore_U_sub_fifo_n209,
         U_afifo_U_acore_U_sub_fifo_n208, U_afifo_U_acore_U_sub_fifo_n207,
         U_afifo_U_acore_U_sub_fifo_n206, U_afifo_U_acore_U_sub_fifo_n205,
         U_afifo_U_acore_U_sub_fifo_n204, U_afifo_U_acore_U_sub_fifo_n203,
         U_afifo_U_acore_U_sub_fifo_n202, U_afifo_U_acore_U_sub_fifo_n201,
         U_afifo_U_acore_U_sub_fifo_n200, U_afifo_U_acore_U_sub_fifo_n199,
         U_afifo_U_acore_U_sub_fifo_n198, U_afifo_U_acore_U_sub_fifo_n197,
         U_afifo_U_acore_U_sub_fifo_n196, U_afifo_U_acore_U_sub_fifo_n195,
         U_afifo_U_acore_U_sub_fifo_n194, U_afifo_U_acore_U_sub_fifo_n193,
         U_afifo_U_acore_U_sub_fifo_n192, U_afifo_U_acore_U_sub_fifo_n191,
         U_afifo_U_acore_U_sub_fifo_n190, U_afifo_U_acore_U_sub_fifo_n189,
         U_afifo_U_acore_U_sub_fifo_n188, U_afifo_U_acore_U_sub_fifo_n187,
         U_afifo_U_acore_U_sub_fifo_n186, U_afifo_U_acore_U_sub_fifo_n185,
         U_afifo_U_acore_U_sub_fifo_n184, U_afifo_U_acore_U_sub_fifo_n183,
         U_afifo_U_acore_U_sub_fifo_n182, U_afifo_U_acore_U_sub_fifo_n181,
         U_afifo_U_acore_U_sub_fifo_n180, U_afifo_U_acore_U_sub_fifo_n179,
         U_afifo_U_acore_U_sub_fifo_n178, U_afifo_U_acore_U_sub_fifo_n177,
         U_afifo_U_acore_U_sub_fifo_n176, U_afifo_U_acore_U_sub_fifo_n175,
         U_afifo_U_acore_U_sub_fifo_n174, U_afifo_U_acore_U_sub_fifo_n173,
         U_afifo_U_acore_U_sub_fifo_n172, U_afifo_U_acore_U_sub_fifo_n171,
         U_afifo_U_acore_U_sub_fifo_n170, U_afifo_U_acore_U_sub_fifo_in_ptr_1_,
         U_afifo_U_acore_U_sub_fifo_count_0_,
         U_afifo_U_acore_U_sub_fifo_count_1_,
         U_afifo_U_acore_U_sub_fifo_out_ptr_0_,
         U_afifo_U_acore_U_sub_fifo_out_ptr_1_,
         U_dfifo_U_dcore_U_sub_fifo_n609, U_dfifo_U_dcore_U_sub_fifo_n608,
         U_dfifo_U_dcore_U_sub_fifo_n607, U_dfifo_U_dcore_U_sub_fifo_n606,
         U_dfifo_U_dcore_U_sub_fifo_n605, U_dfifo_U_dcore_U_sub_fifo_n604,
         U_dfifo_U_dcore_U_sub_fifo_n603, U_dfifo_U_dcore_U_sub_fifo_n602,
         U_dfifo_U_dcore_U_sub_fifo_n567, U_dfifo_U_dcore_U_sub_fifo_n566,
         U_dfifo_U_dcore_U_sub_fifo_n565, U_dfifo_U_dcore_U_sub_fifo_n564,
         U_dfifo_U_dcore_U_sub_fifo_n563, U_dfifo_U_dcore_U_sub_fifo_n562,
         U_dfifo_U_dcore_U_sub_fifo_n561, U_dfifo_U_dcore_U_sub_fifo_n560,
         U_dfifo_U_dcore_U_sub_fifo_n559, U_dfifo_U_dcore_U_sub_fifo_n558,
         U_dfifo_U_dcore_U_sub_fifo_n557, U_dfifo_U_dcore_U_sub_fifo_n556,
         U_dfifo_U_dcore_U_sub_fifo_n555, U_dfifo_U_dcore_U_sub_fifo_n554,
         U_dfifo_U_dcore_U_sub_fifo_n553, U_dfifo_U_dcore_U_sub_fifo_n552,
         U_dfifo_U_dcore_U_sub_fifo_n551, U_dfifo_U_dcore_U_sub_fifo_n550,
         U_dfifo_U_dcore_U_sub_fifo_n549, U_dfifo_U_dcore_U_sub_fifo_n548,
         U_dfifo_U_dcore_U_sub_fifo_n547, U_dfifo_U_dcore_U_sub_fifo_n546,
         U_dfifo_U_dcore_U_sub_fifo_n545, U_dfifo_U_dcore_U_sub_fifo_n544,
         U_dfifo_U_dcore_U_sub_fifo_n543, U_dfifo_U_dcore_U_sub_fifo_n542,
         U_dfifo_U_dcore_U_sub_fifo_n541, U_dfifo_U_dcore_U_sub_fifo_n540,
         U_dfifo_U_dcore_U_sub_fifo_n539, U_dfifo_U_dcore_U_sub_fifo_n538,
         U_dfifo_U_dcore_U_sub_fifo_n537, U_dfifo_U_dcore_U_sub_fifo_n536,
         U_dfifo_U_dcore_U_sub_fifo_n535, U_dfifo_U_dcore_U_sub_fifo_n534,
         U_dfifo_U_dcore_U_sub_fifo_n533, U_dfifo_U_dcore_U_sub_fifo_n532,
         U_dfifo_U_dcore_U_sub_fifo_n531, U_dfifo_U_dcore_U_sub_fifo_n530,
         U_dfifo_U_dcore_U_sub_fifo_n529, U_dfifo_U_dcore_U_sub_fifo_n528,
         U_dfifo_U_dcore_U_sub_fifo_n527, U_dfifo_U_dcore_U_sub_fifo_n526,
         U_dfifo_U_dcore_U_sub_fifo_n525, U_dfifo_U_dcore_U_sub_fifo_n524,
         U_dfifo_U_dcore_U_sub_fifo_n523, U_dfifo_U_dcore_U_sub_fifo_n522,
         U_dfifo_U_dcore_U_sub_fifo_n521, U_dfifo_U_dcore_U_sub_fifo_n520,
         U_dfifo_U_dcore_U_sub_fifo_n519, U_dfifo_U_dcore_U_sub_fifo_n518,
         U_dfifo_U_dcore_U_sub_fifo_n517, U_dfifo_U_dcore_U_sub_fifo_n516,
         U_dfifo_U_dcore_U_sub_fifo_n515, U_dfifo_U_dcore_U_sub_fifo_n514,
         U_dfifo_U_dcore_U_sub_fifo_n513, U_dfifo_U_dcore_U_sub_fifo_n512,
         U_dfifo_U_dcore_U_sub_fifo_n511, U_dfifo_U_dcore_U_sub_fifo_n510,
         U_dfifo_U_dcore_U_sub_fifo_n509, U_dfifo_U_dcore_U_sub_fifo_n508,
         U_dfifo_U_dcore_U_sub_fifo_n507, U_dfifo_U_dcore_U_sub_fifo_n506,
         U_dfifo_U_dcore_U_sub_fifo_n505, U_dfifo_U_dcore_U_sub_fifo_n504,
         U_dfifo_U_dcore_U_sub_fifo_n503, U_dfifo_U_dcore_U_sub_fifo_n502,
         U_dfifo_U_dcore_U_sub_fifo_n501, U_dfifo_U_dcore_U_sub_fifo_n500,
         U_dfifo_U_dcore_U_sub_fifo_n499, U_dfifo_U_dcore_U_sub_fifo_n498,
         U_dfifo_U_dcore_U_sub_fifo_n497, U_dfifo_U_dcore_U_sub_fifo_n496,
         U_dfifo_U_dcore_U_sub_fifo_n495, U_dfifo_U_dcore_U_sub_fifo_n494,
         U_dfifo_U_dcore_U_sub_fifo_n493, U_dfifo_U_dcore_U_sub_fifo_n492,
         U_dfifo_U_dcore_U_sub_fifo_n491, U_dfifo_U_dcore_U_sub_fifo_n490,
         U_dfifo_U_dcore_U_sub_fifo_n489, U_dfifo_U_dcore_U_sub_fifo_n488,
         U_dfifo_U_dcore_U_sub_fifo_n487, U_dfifo_U_dcore_U_sub_fifo_n486,
         U_dfifo_U_dcore_U_sub_fifo_n485, U_dfifo_U_dcore_U_sub_fifo_n484,
         U_dfifo_U_dcore_U_sub_fifo_n483, U_dfifo_U_dcore_U_sub_fifo_n482,
         U_dfifo_U_dcore_U_sub_fifo_n481, U_dfifo_U_dcore_U_sub_fifo_n480,
         U_dfifo_U_dcore_U_sub_fifo_n479, U_dfifo_U_dcore_U_sub_fifo_n478,
         U_dfifo_U_dcore_U_sub_fifo_n477, U_dfifo_U_dcore_U_sub_fifo_n476,
         U_dfifo_U_dcore_U_sub_fifo_n475, U_dfifo_U_dcore_U_sub_fifo_n474,
         U_dfifo_U_dcore_U_sub_fifo_n473, U_dfifo_U_dcore_U_sub_fifo_n472,
         U_dfifo_U_dcore_U_sub_fifo_n471, U_dfifo_U_dcore_U_sub_fifo_n470,
         U_dfifo_U_dcore_U_sub_fifo_n469, U_dfifo_U_dcore_U_sub_fifo_n468,
         U_dfifo_U_dcore_U_sub_fifo_n467, U_dfifo_U_dcore_U_sub_fifo_n466,
         U_dfifo_U_dcore_U_sub_fifo_n465, U_dfifo_U_dcore_U_sub_fifo_n464,
         U_dfifo_U_dcore_U_sub_fifo_n463, U_dfifo_U_dcore_U_sub_fifo_n462,
         U_dfifo_U_dcore_U_sub_fifo_n461, U_dfifo_U_dcore_U_sub_fifo_n460,
         U_dfifo_U_dcore_U_sub_fifo_n459, U_dfifo_U_dcore_U_sub_fifo_n458,
         U_dfifo_U_dcore_U_sub_fifo_n456, U_dfifo_U_dcore_U_sub_fifo_n455,
         U_dfifo_U_dcore_U_sub_fifo_n241, U_dfifo_U_dcore_U_sub_fifo_n235,
         U_dfifo_U_dcore_U_sub_fifo_n234, U_dfifo_U_dcore_U_sub_fifo_n233,
         U_dfifo_U_dcore_U_sub_fifo_n232, U_dfifo_U_dcore_U_sub_fifo_n231,
         U_dfifo_U_dcore_U_sub_fifo_n230, U_dfifo_U_dcore_U_sub_fifo_n229,
         U_dfifo_U_dcore_U_sub_fifo_n228, U_dfifo_U_dcore_U_sub_fifo_n227,
         U_dfifo_U_dcore_U_sub_fifo_n226, U_dfifo_U_dcore_U_sub_fifo_n225,
         U_dfifo_U_dcore_U_sub_fifo_n224, U_dfifo_U_dcore_U_sub_fifo_n223,
         U_dfifo_U_dcore_U_sub_fifo_n222, U_dfifo_U_dcore_U_sub_fifo_n221,
         U_dfifo_U_dcore_U_sub_fifo_n220, U_dfifo_U_dcore_U_sub_fifo_n219,
         U_dfifo_U_dcore_U_sub_fifo_n218, U_dfifo_U_dcore_U_sub_fifo_n217,
         U_dfifo_U_dcore_U_sub_fifo_n216, U_dfifo_U_dcore_U_sub_fifo_n215,
         U_dfifo_U_dcore_U_sub_fifo_n214, U_dfifo_U_dcore_U_sub_fifo_n213,
         U_dfifo_U_dcore_U_sub_fifo_n212, U_dfifo_U_dcore_U_sub_fifo_n211,
         U_dfifo_U_dcore_U_sub_fifo_n210, U_dfifo_U_dcore_U_sub_fifo_n209,
         U_dfifo_U_dcore_U_sub_fifo_n208, U_dfifo_U_dcore_U_sub_fifo_n207,
         U_dfifo_U_dcore_U_sub_fifo_n206, U_dfifo_U_dcore_U_sub_fifo_n205,
         U_dfifo_U_dcore_U_sub_fifo_n204, U_dfifo_U_dcore_U_sub_fifo_n203,
         U_dfifo_U_dcore_U_sub_fifo_n202, U_dfifo_U_dcore_U_sub_fifo_n201,
         U_dfifo_U_dcore_U_sub_fifo_n200, U_dfifo_U_dcore_U_sub_fifo_n199,
         U_dfifo_U_dcore_U_sub_fifo_n198, U_dfifo_U_dcore_U_sub_fifo_n197,
         U_dfifo_U_dcore_U_sub_fifo_n196, U_dfifo_U_dcore_U_sub_fifo_n195,
         U_dfifo_U_dcore_U_sub_fifo_n194, U_dfifo_U_dcore_U_sub_fifo_n193,
         U_dfifo_U_dcore_U_sub_fifo_n192, U_dfifo_U_dcore_U_sub_fifo_n191,
         U_dfifo_U_dcore_U_sub_fifo_n190, U_dfifo_U_dcore_U_sub_fifo_n189,
         U_dfifo_U_dcore_U_sub_fifo_n188, U_dfifo_U_dcore_U_sub_fifo_n187,
         U_dfifo_U_dcore_U_sub_fifo_n186, U_dfifo_U_dcore_U_sub_fifo_n185,
         U_dfifo_U_dcore_U_sub_fifo_n184, U_dfifo_U_dcore_U_sub_fifo_n183,
         U_dfifo_U_dcore_U_sub_fifo_n182, U_dfifo_U_dcore_U_sub_fifo_n181,
         U_dfifo_U_dcore_U_sub_fifo_n180, U_dfifo_U_dcore_U_sub_fifo_n179,
         U_dfifo_U_dcore_U_sub_fifo_n178, U_dfifo_U_dcore_U_sub_fifo_n177,
         U_dfifo_U_dcore_U_sub_fifo_n176, U_dfifo_U_dcore_U_sub_fifo_n175,
         U_dfifo_U_dcore_U_sub_fifo_n174, U_dfifo_U_dcore_U_sub_fifo_n173,
         U_dfifo_U_dcore_U_sub_fifo_n172, U_dfifo_U_dcore_U_sub_fifo_n171,
         U_dfifo_U_dcore_U_sub_fifo_n170, U_dfifo_U_dcore_U_sub_fifo_n169,
         U_dfifo_U_dcore_U_sub_fifo_n168, U_dfifo_U_dcore_U_sub_fifo_n167,
         U_dfifo_U_dcore_U_sub_fifo_n166, U_dfifo_U_dcore_U_sub_fifo_n165,
         U_dfifo_U_dcore_U_sub_fifo_n164, U_dfifo_U_dcore_U_sub_fifo_n163,
         U_dfifo_U_dcore_U_sub_fifo_n162, U_dfifo_U_dcore_U_sub_fifo_n161,
         U_dfifo_U_dcore_U_sub_fifo_n160, U_dfifo_U_dcore_U_sub_fifo_n159,
         U_dfifo_U_dcore_U_sub_fifo_n158, U_dfifo_U_dcore_U_sub_fifo_n157,
         U_dfifo_U_dcore_U_sub_fifo_n156, U_dfifo_U_dcore_U_sub_fifo_n155,
         U_dfifo_U_dcore_U_sub_fifo_n154, U_dfifo_U_dcore_U_sub_fifo_n153,
         U_dfifo_U_dcore_U_sub_fifo_n152, U_dfifo_U_dcore_U_sub_fifo_n151,
         U_dfifo_U_dcore_U_sub_fifo_n150, U_dfifo_U_dcore_U_sub_fifo_n149,
         U_dfifo_U_dcore_U_sub_fifo_n148, U_dfifo_U_dcore_U_sub_fifo_n147,
         U_dfifo_U_dcore_U_sub_fifo_n146, U_dfifo_U_dcore_U_sub_fifo_n145,
         U_dfifo_U_dcore_U_sub_fifo_n144, U_dfifo_U_dcore_U_sub_fifo_n143,
         U_dfifo_U_dcore_U_sub_fifo_n142, U_dfifo_U_dcore_U_sub_fifo_n141,
         U_dfifo_U_dcore_U_sub_fifo_n140, U_dfifo_U_dcore_U_sub_fifo_n139,
         U_dfifo_U_dcore_U_sub_fifo_n138, U_dfifo_U_dcore_U_sub_fifo_n137,
         U_dfifo_U_dcore_U_sub_fifo_n136, U_dfifo_U_dcore_U_sub_fifo_n135,
         U_dfifo_U_dcore_U_sub_fifo_n134, U_dfifo_U_dcore_U_sub_fifo_n133,
         U_dfifo_U_dcore_U_sub_fifo_n132, U_dfifo_U_dcore_U_sub_fifo_n131,
         U_dfifo_U_dcore_U_sub_fifo_n130, U_dfifo_U_dcore_U_sub_fifo_n129,
         U_dfifo_U_dcore_U_sub_fifo_n128, U_dfifo_U_dcore_U_sub_fifo_n127,
         U_dfifo_U_dcore_U_sub_fifo_n126, U_dfifo_U_dcore_U_sub_fifo_n125,
         U_dfifo_U_dcore_U_sub_fifo_n124, U_dfifo_U_dcore_U_sub_fifo_n123,
         U_dfifo_U_dcore_U_sub_fifo_n122, U_dfifo_U_dcore_U_sub_fifo_n121,
         U_dfifo_U_dcore_U_sub_fifo_n120, U_dfifo_U_dcore_U_sub_fifo_n119,
         U_dfifo_U_dcore_U_sub_fifo_n118, U_dfifo_U_dcore_U_sub_fifo_n117,
         U_dfifo_U_dcore_U_sub_fifo_n116, U_dfifo_U_dcore_U_sub_fifo_n115,
         U_dfifo_U_dcore_U_sub_fifo_n114, U_dfifo_U_dcore_U_sub_fifo_n113,
         U_dfifo_U_dcore_U_sub_fifo_n112, U_dfifo_U_dcore_U_sub_fifo_n111,
         U_dfifo_U_dcore_U_sub_fifo_n110, U_dfifo_U_dcore_U_sub_fifo_n109,
         U_dfifo_U_dcore_U_sub_fifo_n108, U_dfifo_U_dcore_U_sub_fifo_n107,
         U_dfifo_U_dcore_U_sub_fifo_n106, U_dfifo_U_dcore_U_sub_fifo_n105,
         U_dfifo_U_dcore_U_sub_fifo_n104, U_dfifo_U_dcore_U_sub_fifo_n103,
         U_dfifo_U_dcore_U_sub_fifo_n102, U_dfifo_U_dcore_U_sub_fifo_n101,
         U_dfifo_U_dcore_U_sub_fifo_n100, U_dfifo_U_dcore_U_sub_fifo_n99,
         U_dfifo_U_dcore_U_sub_fifo_n98, U_dfifo_U_dcore_U_sub_fifo_n97,
         U_dfifo_U_dcore_U_sub_fifo_n96, U_dfifo_U_dcore_U_sub_fifo_n95,
         U_dfifo_U_dcore_U_sub_fifo_n94, U_dfifo_U_dcore_U_sub_fifo_n93,
         U_dfifo_U_dcore_U_sub_fifo_n92, U_dfifo_U_dcore_U_sub_fifo_n91,
         U_dfifo_U_dcore_U_sub_fifo_n90, U_dfifo_U_dcore_U_sub_fifo_n89,
         U_dfifo_U_dcore_U_sub_fifo_n88, U_dfifo_U_dcore_U_sub_fifo_n87,
         U_dfifo_U_dcore_U_sub_fifo_n86, U_dfifo_U_dcore_U_sub_fifo_n85,
         U_dfifo_U_dcore_U_sub_fifo_n84, U_dfifo_U_dcore_U_sub_fifo_n83,
         U_dfifo_U_dcore_U_sub_fifo_n82, U_dfifo_U_dcore_U_sub_fifo_n81,
         U_dfifo_U_dcore_U_sub_fifo_n80, U_dfifo_U_dcore_U_sub_fifo_n79,
         U_dfifo_U_dcore_U_sub_fifo_n78, U_dfifo_U_dcore_U_sub_fifo_n77,
         U_dfifo_U_dcore_U_sub_fifo_n76, U_dfifo_U_dcore_U_sub_fifo_n75,
         U_dfifo_U_dcore_U_sub_fifo_n74, U_dfifo_U_dcore_U_sub_fifo_n73,
         U_dfifo_U_dcore_U_sub_fifo_n72, U_dfifo_U_dcore_U_sub_fifo_n71,
         U_dfifo_U_dcore_U_sub_fifo_n70, U_dfifo_U_dcore_U_sub_fifo_n69,
         U_dfifo_U_dcore_U_sub_fifo_n68, U_dfifo_U_dcore_U_sub_fifo_n67,
         U_dfifo_U_dcore_U_sub_fifo_n66, U_dfifo_U_dcore_U_sub_fifo_n65,
         U_dfifo_U_dcore_U_sub_fifo_n64, U_dfifo_U_dcore_U_sub_fifo_n63,
         U_dfifo_U_dcore_U_sub_fifo_n62, U_dfifo_U_dcore_U_sub_fifo_n61,
         U_dfifo_U_dcore_U_sub_fifo_n60, U_dfifo_U_dcore_U_sub_fifo_n59,
         U_dfifo_U_dcore_U_sub_fifo_n58, U_dfifo_U_dcore_U_sub_fifo_n57,
         U_dfifo_U_dcore_U_sub_fifo_n56, U_dfifo_U_dcore_U_sub_fifo_n55,
         U_dfifo_U_dcore_U_sub_fifo_n54, U_dfifo_U_dcore_U_sub_fifo_n53,
         U_dfifo_U_dcore_U_sub_fifo_n52, U_dfifo_U_dcore_U_sub_fifo_n51,
         U_dfifo_U_dcore_U_sub_fifo_n50, U_dfifo_U_dcore_U_sub_fifo_n49,
         U_dfifo_U_dcore_U_sub_fifo_n48, U_dfifo_U_dcore_U_sub_fifo_n47,
         U_dfifo_U_dcore_U_sub_fifo_n46, U_dfifo_U_dcore_U_sub_fifo_n45,
         U_dfifo_U_dcore_U_sub_fifo_n44, U_dfifo_U_dcore_U_sub_fifo_n43,
         U_dfifo_U_dcore_U_sub_fifo_n42, U_dfifo_U_dcore_U_sub_fifo_n41,
         U_dfifo_U_dcore_U_sub_fifo_n40, U_dfifo_U_dcore_U_sub_fifo_n39,
         U_dfifo_U_dcore_U_sub_fifo_n38, U_dfifo_U_dcore_U_sub_fifo_n37,
         U_dfifo_U_dcore_U_sub_fifo_n36, U_dfifo_U_dcore_U_sub_fifo_n35,
         U_dfifo_U_dcore_U_sub_fifo_n34, U_dfifo_U_dcore_U_sub_fifo_n33,
         U_dfifo_U_dcore_U_sub_fifo_n32, U_dfifo_U_dcore_U_sub_fifo_n31,
         U_dfifo_U_dcore_U_sub_fifo_n30, U_dfifo_U_dcore_U_sub_fifo_n29,
         U_dfifo_U_dcore_U_sub_fifo_n28, U_dfifo_U_dcore_U_sub_fifo_n27,
         U_dfifo_U_dcore_U_sub_fifo_n26, U_dfifo_U_dcore_U_sub_fifo_n25,
         U_dfifo_U_dcore_U_sub_fifo_n24, U_dfifo_U_dcore_U_sub_fifo_n23,
         U_dfifo_U_dcore_U_sub_fifo_n22, U_dfifo_U_dcore_U_sub_fifo_n21,
         U_dfifo_U_dcore_U_sub_fifo_n20, U_dfifo_U_dcore_U_sub_fifo_n19,
         U_dfifo_U_dcore_U_sub_fifo_n18, U_dfifo_U_dcore_U_sub_fifo_n17,
         U_dfifo_U_dcore_U_sub_fifo_n16, U_dfifo_U_dcore_U_sub_fifo_n15,
         U_dfifo_U_dcore_U_sub_fifo_n14, U_dfifo_U_dcore_U_sub_fifo_n13,
         U_dfifo_U_dcore_U_sub_fifo_n12, U_dfifo_U_dcore_U_sub_fifo_n11,
         U_dfifo_U_dcore_U_sub_fifo_n10, U_dfifo_U_dcore_U_sub_fifo_n9,
         U_dfifo_U_dcore_U_sub_fifo_n8, U_dfifo_U_dcore_U_sub_fifo_n7,
         U_dfifo_U_dcore_U_sub_fifo_n6, U_dfifo_U_dcore_U_sub_fifo_n5,
         U_dfifo_U_dcore_U_sub_fifo_n4, U_dfifo_U_dcore_U_sub_fifo_n3,
         U_dfifo_U_dcore_U_sub_fifo_n1, U_dfifo_U_dcore_U_sub_fifo_n454,
         U_dfifo_U_dcore_U_sub_fifo_n453, U_dfifo_U_dcore_U_sub_fifo_n452,
         U_dfifo_U_dcore_U_sub_fifo_n451, U_dfifo_U_dcore_U_sub_fifo_n450,
         U_dfifo_U_dcore_U_sub_fifo_n449, U_dfifo_U_dcore_U_sub_fifo_n448,
         U_dfifo_U_dcore_U_sub_fifo_n447, U_dfifo_U_dcore_U_sub_fifo_n446,
         U_dfifo_U_dcore_U_sub_fifo_n445, U_dfifo_U_dcore_U_sub_fifo_n444,
         U_dfifo_U_dcore_U_sub_fifo_n443, U_dfifo_U_dcore_U_sub_fifo_n442,
         U_dfifo_U_dcore_U_sub_fifo_n441, U_dfifo_U_dcore_U_sub_fifo_n440,
         U_dfifo_U_dcore_U_sub_fifo_n439, U_dfifo_U_dcore_U_sub_fifo_n438,
         U_dfifo_U_dcore_U_sub_fifo_n437, U_dfifo_U_dcore_U_sub_fifo_n436,
         U_dfifo_U_dcore_U_sub_fifo_n435, U_dfifo_U_dcore_U_sub_fifo_n434,
         U_dfifo_U_dcore_U_sub_fifo_n433, U_dfifo_U_dcore_U_sub_fifo_n432,
         U_dfifo_U_dcore_U_sub_fifo_n431, U_dfifo_U_dcore_U_sub_fifo_n430,
         U_dfifo_U_dcore_U_sub_fifo_n429, U_dfifo_U_dcore_U_sub_fifo_n428,
         U_dfifo_U_dcore_U_sub_fifo_n427, U_dfifo_U_dcore_U_sub_fifo_n426,
         U_dfifo_U_dcore_U_sub_fifo_n425, U_dfifo_U_dcore_U_sub_fifo_n424,
         U_dfifo_U_dcore_U_sub_fifo_n423, U_dfifo_U_dcore_U_sub_fifo_n422,
         U_dfifo_U_dcore_U_sub_fifo_n421, U_dfifo_U_dcore_U_sub_fifo_n420,
         U_dfifo_U_dcore_U_sub_fifo_n419, U_dfifo_U_dcore_U_sub_fifo_n418,
         U_dfifo_U_dcore_U_sub_fifo_n417, U_dfifo_U_dcore_U_sub_fifo_n416,
         U_dfifo_U_dcore_U_sub_fifo_n415, U_dfifo_U_dcore_U_sub_fifo_n414,
         U_dfifo_U_dcore_U_sub_fifo_n413, U_dfifo_U_dcore_U_sub_fifo_n412,
         U_dfifo_U_dcore_U_sub_fifo_n411, U_dfifo_U_dcore_U_sub_fifo_n410,
         U_dfifo_U_dcore_U_sub_fifo_n409, U_dfifo_U_dcore_U_sub_fifo_n408,
         U_dfifo_U_dcore_U_sub_fifo_n407, U_dfifo_U_dcore_U_sub_fifo_n406,
         U_dfifo_U_dcore_U_sub_fifo_n405, U_dfifo_U_dcore_U_sub_fifo_n404,
         U_dfifo_U_dcore_U_sub_fifo_n403, U_dfifo_U_dcore_U_sub_fifo_n402,
         U_dfifo_U_dcore_U_sub_fifo_n401, U_dfifo_U_dcore_U_sub_fifo_n400,
         U_dfifo_U_dcore_U_sub_fifo_n399, U_dfifo_U_dcore_U_sub_fifo_n398,
         U_dfifo_U_dcore_U_sub_fifo_n397, U_dfifo_U_dcore_U_sub_fifo_n396,
         U_dfifo_U_dcore_U_sub_fifo_n395, U_dfifo_U_dcore_U_sub_fifo_n394,
         U_dfifo_U_dcore_U_sub_fifo_n393, U_dfifo_U_dcore_U_sub_fifo_n392,
         U_dfifo_U_dcore_U_sub_fifo_n391, U_dfifo_U_dcore_U_sub_fifo_n390,
         U_dfifo_U_dcore_U_sub_fifo_n389, U_dfifo_U_dcore_U_sub_fifo_n388,
         U_dfifo_U_dcore_U_sub_fifo_n387, U_dfifo_U_dcore_U_sub_fifo_n386,
         U_dfifo_U_dcore_U_sub_fifo_n385, U_dfifo_U_dcore_U_sub_fifo_n384,
         U_dfifo_U_dcore_U_sub_fifo_n383, U_dfifo_U_dcore_U_sub_fifo_n382,
         U_dfifo_U_dcore_U_sub_fifo_n381, U_dfifo_U_dcore_U_sub_fifo_n380,
         U_dfifo_U_dcore_U_sub_fifo_n379, U_dfifo_U_dcore_U_sub_fifo_n378,
         U_dfifo_U_dcore_U_sub_fifo_n377, U_dfifo_U_dcore_U_sub_fifo_n376,
         U_dfifo_U_dcore_U_sub_fifo_n375, U_dfifo_U_dcore_U_sub_fifo_n374,
         U_dfifo_U_dcore_U_sub_fifo_n373, U_dfifo_U_dcore_U_sub_fifo_n372,
         U_dfifo_U_dcore_U_sub_fifo_n371, U_dfifo_U_dcore_U_sub_fifo_n370,
         U_dfifo_U_dcore_U_sub_fifo_n369, U_dfifo_U_dcore_U_sub_fifo_n368,
         U_dfifo_U_dcore_U_sub_fifo_n367, U_dfifo_U_dcore_U_sub_fifo_n366,
         U_dfifo_U_dcore_U_sub_fifo_n365, U_dfifo_U_dcore_U_sub_fifo_n364,
         U_dfifo_U_dcore_U_sub_fifo_n363, U_dfifo_U_dcore_U_sub_fifo_n362,
         U_dfifo_U_dcore_U_sub_fifo_n361, U_dfifo_U_dcore_U_sub_fifo_n360,
         U_dfifo_U_dcore_U_sub_fifo_n359, U_dfifo_U_dcore_U_sub_fifo_n358,
         U_dfifo_U_dcore_U_sub_fifo_n357, U_dfifo_U_dcore_U_sub_fifo_n356,
         U_dfifo_U_dcore_U_sub_fifo_n355, U_dfifo_U_dcore_U_sub_fifo_n354,
         U_dfifo_U_dcore_U_sub_fifo_n353, U_dfifo_U_dcore_U_sub_fifo_n352,
         U_dfifo_U_dcore_U_sub_fifo_n351, U_dfifo_U_dcore_U_sub_fifo_n350,
         U_dfifo_U_dcore_U_sub_fifo_n349, U_dfifo_U_dcore_U_sub_fifo_n348,
         U_dfifo_U_dcore_U_sub_fifo_n347, U_dfifo_U_dcore_U_sub_fifo_n346,
         U_dfifo_U_dcore_U_sub_fifo_n345, U_dfifo_U_dcore_U_sub_fifo_n344,
         U_dfifo_U_dcore_U_sub_fifo_n343, U_dfifo_U_dcore_U_sub_fifo_n342,
         U_dfifo_U_dcore_U_sub_fifo_n341, U_dfifo_U_dcore_U_sub_fifo_n340,
         U_dfifo_U_dcore_U_sub_fifo_n339, U_dfifo_U_dcore_U_sub_fifo_n338,
         U_dfifo_U_dcore_U_sub_fifo_n337, U_dfifo_U_dcore_U_sub_fifo_n336,
         U_dfifo_U_dcore_U_sub_fifo_n335, U_dfifo_U_dcore_U_sub_fifo_n334,
         U_dfifo_U_dcore_U_sub_fifo_n333, U_dfifo_U_dcore_U_sub_fifo_n332,
         U_dfifo_U_dcore_U_sub_fifo_n331, U_dfifo_U_dcore_U_sub_fifo_n330,
         U_dfifo_U_dcore_U_sub_fifo_n329, U_dfifo_U_dcore_U_sub_fifo_n328,
         U_dfifo_U_dcore_U_sub_fifo_n327, U_dfifo_U_dcore_U_sub_fifo_n326,
         U_dfifo_U_dcore_U_sub_fifo_n325, U_dfifo_U_dcore_U_sub_fifo_n324,
         U_dfifo_U_dcore_U_sub_fifo_n323, U_dfifo_U_dcore_U_sub_fifo_n322,
         U_dfifo_U_dcore_U_sub_fifo_n321, U_dfifo_U_dcore_U_sub_fifo_n320,
         U_dfifo_U_dcore_U_sub_fifo_n319, U_dfifo_U_dcore_U_sub_fifo_n318,
         U_dfifo_U_dcore_U_sub_fifo_n317, U_dfifo_U_dcore_U_sub_fifo_n316,
         U_dfifo_U_dcore_U_sub_fifo_n315, U_dfifo_U_dcore_U_sub_fifo_n314,
         U_dfifo_U_dcore_U_sub_fifo_n313, U_dfifo_U_dcore_U_sub_fifo_n312,
         U_dfifo_U_dcore_U_sub_fifo_n311, U_dfifo_U_dcore_U_sub_fifo_n310,
         U_dfifo_U_dcore_U_sub_fifo_n309, U_dfifo_U_dcore_U_sub_fifo_n308,
         U_dfifo_U_dcore_U_sub_fifo_n307, U_dfifo_U_dcore_U_sub_fifo_n306,
         U_dfifo_U_dcore_U_sub_fifo_n305, U_dfifo_U_dcore_U_sub_fifo_n304,
         U_dfifo_U_dcore_U_sub_fifo_n303, U_dfifo_U_dcore_U_sub_fifo_n302,
         U_dfifo_U_dcore_U_sub_fifo_n301, U_dfifo_U_dcore_U_sub_fifo_n300,
         U_dfifo_U_dcore_U_sub_fifo_n299, U_dfifo_U_dcore_U_sub_fifo_n298,
         U_dfifo_U_dcore_U_sub_fifo_n297, U_dfifo_U_dcore_U_sub_fifo_n296,
         U_dfifo_U_dcore_U_sub_fifo_n295, U_dfifo_U_dcore_U_sub_fifo_n294,
         U_dfifo_U_dcore_U_sub_fifo_n293, U_dfifo_U_dcore_U_sub_fifo_n292,
         U_dfifo_U_dcore_U_sub_fifo_n291, U_dfifo_U_dcore_U_sub_fifo_n290,
         U_dfifo_U_dcore_U_sub_fifo_n289, U_dfifo_U_dcore_U_sub_fifo_n288,
         U_dfifo_U_dcore_U_sub_fifo_n287, U_dfifo_U_dcore_U_sub_fifo_n286,
         U_dfifo_U_dcore_U_sub_fifo_n285, U_dfifo_U_dcore_U_sub_fifo_n284,
         U_dfifo_U_dcore_U_sub_fifo_n283, U_dfifo_U_dcore_U_sub_fifo_n282,
         U_dfifo_U_dcore_U_sub_fifo_n281, U_dfifo_U_dcore_U_sub_fifo_n280,
         U_dfifo_U_dcore_U_sub_fifo_n279, U_dfifo_U_dcore_U_sub_fifo_n278,
         U_dfifo_U_dcore_U_sub_fifo_n277, U_dfifo_U_dcore_U_sub_fifo_n276,
         U_dfifo_U_dcore_U_sub_fifo_n275, U_dfifo_U_dcore_U_sub_fifo_n274,
         U_dfifo_U_dcore_U_sub_fifo_n273, U_dfifo_U_dcore_U_sub_fifo_n272,
         U_dfifo_U_dcore_U_sub_fifo_n271, U_dfifo_U_dcore_U_sub_fifo_n270,
         U_dfifo_U_dcore_U_sub_fifo_n269, U_dfifo_U_dcore_U_sub_fifo_n268,
         U_dfifo_U_dcore_U_sub_fifo_n267, U_dfifo_U_dcore_U_sub_fifo_n266,
         U_dfifo_U_dcore_U_sub_fifo_n265, U_dfifo_U_dcore_U_sub_fifo_n264,
         U_dfifo_U_dcore_U_sub_fifo_n263, U_dfifo_U_dcore_U_sub_fifo_n262,
         U_dfifo_U_dcore_U_sub_fifo_n261, U_dfifo_U_dcore_U_sub_fifo_n260,
         U_dfifo_U_dcore_U_sub_fifo_n259, U_dfifo_U_dcore_U_sub_fifo_n258,
         U_dfifo_U_dcore_U_sub_fifo_n257, U_dfifo_U_dcore_U_sub_fifo_n256,
         U_dfifo_U_dcore_U_sub_fifo_n255, U_dfifo_U_dcore_U_sub_fifo_n254,
         U_dfifo_U_dcore_U_sub_fifo_n253, U_dfifo_U_dcore_U_sub_fifo_n252,
         U_dfifo_U_dcore_U_sub_fifo_n251, U_dfifo_U_dcore_U_sub_fifo_n250,
         U_dfifo_U_dcore_U_sub_fifo_n249, U_dfifo_U_dcore_U_sub_fifo_n248,
         U_dfifo_U_dcore_U_sub_fifo_n247, U_dfifo_U_dcore_U_sub_fifo_n246,
         U_dfifo_U_dcore_U_sub_fifo_n245, U_dfifo_U_dcore_U_sub_fifo_n244,
         U_dfifo_U_dcore_U_sub_fifo_n243, U_dfifo_U_dcore_U_sub_fifo_n242,
         U_dfifo_U_dcore_U_sub_fifo_in_ptr_0_,
         U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_,
         U_dfifo_U_dcore_U_sub_fifo_in_ptr_2_,
         U_dfifo_U_dcore_U_sub_fifo_count_0_,
         U_dfifo_U_dcore_U_sub_fifo_count_1_,
         U_dfifo_U_dcore_U_sub_fifo_count_2_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__0_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__1_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__2_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__3_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__4_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__5_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__6_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__7_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__8_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__9_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__10_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__11_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__12_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__13_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__14_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__15_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__16_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__17_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__18_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__19_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__20_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__21_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__22_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__23_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__24_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__25_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__26_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__27_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__28_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__29_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__30_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__31_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__32_,
         U_dfifo_U_dcore_U_sub_fifo_mem_0__33_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__0_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__1_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__2_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__3_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__4_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__5_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__6_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__7_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__8_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__9_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__10_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__11_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__12_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__13_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__14_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__15_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__16_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__17_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__18_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__19_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__20_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__21_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__22_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__23_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__24_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__25_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__26_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__27_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__28_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__29_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__30_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__31_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__32_,
         U_dfifo_U_dcore_U_sub_fifo_mem_2__33_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__0_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__1_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__2_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__3_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__4_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__5_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__6_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__7_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__8_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__9_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__10_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__11_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__12_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__13_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__14_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__15_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__16_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__17_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__18_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__19_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__20_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__21_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__22_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__23_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__24_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__25_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__26_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__27_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__28_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__29_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__30_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__31_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__32_,
         U_dfifo_U_dcore_U_sub_fifo_mem_3__33_,
         U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_,
         U_dfifo_U_dcore_U_sub_fifo_out_ptr_1_,
         U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;
  wire   [16:4] m_af_data2_in;
  wire   [33:0] m_df_data_in;
  wire   [49:0] U_afifo_m_data_in;
  wire   [15:0] U_dfifo_m_btm_data;
  wire   [2:0] U_ctl_n_bh_state;
  wire   [3:0] U_ctl_f_amba_bsz2;
  wire   [3:0] U_ctl_f_col_width;
  wire   [49:0] U_afifo_U_acore_m_sf_data_out;
  wire   [33:0] U_dfifo_U_dcore_m_sf_data_out;

  INV_X4 U1 ( .A(n7), .ZN(n8) );
  INV_X4 U2 ( .A(hsel_mem), .ZN(n7) );
  NAND2_X2 U_afifo_U299 ( .A1(U_afifo_m_data_out_49), .A2(U_afifo_n153), .ZN(
        U_afifo_n259) );
  AND2_X4 U_afifo_U298 ( .A1(U_afifo_m_pop_n), .A2(U_afifo_m_full), .ZN(
        U_afifo_n156) );
  NAND2_X1 U_afifo_U297 ( .A1(U_afifo_m_pop_n), .A2(U_afifo_m_afull), .ZN(
        U_afifo_n168) );
  AOI22_X2 U_afifo_U293 ( .A1(m_af_data1_in_7_), .A2(U_afifo_n98), .B1(
        U_afifo_f_data2_7_), .B2(U_afifo_n54), .ZN(U_afifo_n181) );
  INV_X4 U_afifo_U292 ( .A(U_afifo_n181), .ZN(U_afifo_m_data_in[7]) );
  AOI21_X2 U_afifo_U291 ( .B1(m_af_data1_in_8_), .B2(U_afifo_n99), .A(
        U_afifo_n152), .ZN(U_afifo_n182) );
  INV_X4 U_afifo_U290 ( .A(U_afifo_n182), .ZN(U_afifo_m_data_in[8]) );
  NAND2_X2 U_afifo_U289 ( .A1(n47), .A2(m_af_data2_in[12]), .ZN(U_afifo_n252)
         );
  OAI21_X2 U_afifo_U288 ( .B1(n47), .B2(U_afifo_n165), .A(U_afifo_n252), .ZN(
        U_afifo_n51) );
  OAI21_X2 U_afifo_U287 ( .B1(n47), .B2(U_afifo_n159), .A(U_afifo_n252), .ZN(
        U_afifo_n16) );
  NAND2_X2 U_afifo_U286 ( .A1(n47), .A2(m_af_data2_in[13]), .ZN(U_afifo_n253)
         );
  OAI21_X2 U_afifo_U285 ( .B1(n47), .B2(U_afifo_n166), .A(U_afifo_n253), .ZN(
        U_afifo_n52) );
  OAI21_X2 U_afifo_U284 ( .B1(n47), .B2(U_afifo_n160), .A(U_afifo_n253), .ZN(
        U_afifo_n17) );
  NAND2_X2 U_afifo_U283 ( .A1(m_af_data2_in[5]), .A2(n47), .ZN(U_afifo_n172)
         );
  NAND2_X2 U_afifo_U282 ( .A1(U_afifo_f_data2_5_), .A2(U_afifo_n176), .ZN(
        U_afifo_n173) );
  NAND2_X2 U_afifo_U281 ( .A1(U_afifo_n172), .A2(U_afifo_n173), .ZN(
        U_afifo_n154) );
  OAI21_X2 U_afifo_U280 ( .B1(U_afifo_f_core_ready), .B2(U_afifo_n157), .A(
        U_afifo_n176), .ZN(U_afifo_n3) );
  NAND2_X2 U_afifo_U279 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_0_), .ZN(
        U_afifo_n186) );
  OAI21_X2 U_afifo_U278 ( .B1(U_afifo_n174), .B2(U_afifo_n187), .A(
        U_afifo_n186), .ZN(U_afifo_n4) );
  NAND2_X2 U_afifo_U277 ( .A1(m_af_data2_in[4]), .A2(n47), .ZN(U_afifo_n190)
         );
  OAI21_X2 U_afifo_U276 ( .B1(n47), .B2(U_afifo_n191), .A(U_afifo_n190), .ZN(
        U_afifo_n8) );
  NAND2_X2 U_afifo_U275 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_31_), .ZN(
        U_afifo_n224) );
  OAI21_X2 U_afifo_U274 ( .B1(U_afifo_n174), .B2(U_afifo_n225), .A(
        U_afifo_n224), .ZN(U_afifo_n35) );
  NAND2_X2 U_afifo_U273 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_44_), .ZN(
        U_afifo_n250) );
  OAI21_X2 U_afifo_U272 ( .B1(U_afifo_n174), .B2(U_ctl_n381), .A(U_afifo_n250), 
        .ZN(U_afifo_n48) );
  NAND2_X2 U_afifo_U271 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_20_), .ZN(
        U_afifo_n202) );
  OAI21_X2 U_afifo_U270 ( .B1(U_afifo_n174), .B2(U_afifo_n203), .A(
        U_afifo_n202), .ZN(U_afifo_n24) );
  NAND2_X2 U_afifo_U269 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_27_), .ZN(
        U_afifo_n216) );
  OAI21_X2 U_afifo_U268 ( .B1(U_afifo_n174), .B2(U_afifo_n217), .A(
        U_afifo_n216), .ZN(U_afifo_n31) );
  NAND2_X2 U_afifo_U267 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_18_), .ZN(
        U_afifo_n198) );
  OAI21_X2 U_afifo_U266 ( .B1(U_afifo_n174), .B2(U_ctl_n16), .A(U_afifo_n198), 
        .ZN(U_afifo_n22) );
  NAND2_X2 U_afifo_U265 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_26_), .ZN(
        U_afifo_n214) );
  OAI21_X2 U_afifo_U264 ( .B1(U_afifo_n174), .B2(U_afifo_n215), .A(
        U_afifo_n214), .ZN(U_afifo_n30) );
  NAND2_X2 U_afifo_U263 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_33_), .ZN(
        U_afifo_n228) );
  OAI21_X2 U_afifo_U262 ( .B1(U_afifo_n174), .B2(U_afifo_n229), .A(
        U_afifo_n228), .ZN(U_afifo_n37) );
  NAND2_X2 U_afifo_U261 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_19_), .ZN(
        U_afifo_n200) );
  OAI21_X2 U_afifo_U260 ( .B1(U_afifo_n174), .B2(U_afifo_n201), .A(
        U_afifo_n200), .ZN(U_afifo_n23) );
  NAND2_X2 U_afifo_U259 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_32_), .ZN(
        U_afifo_n226) );
  OAI21_X2 U_afifo_U258 ( .B1(U_afifo_n174), .B2(U_afifo_n227), .A(
        U_afifo_n226), .ZN(U_afifo_n36) );
  NAND2_X2 U_afifo_U257 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_22_), .ZN(
        U_afifo_n206) );
  OAI21_X2 U_afifo_U256 ( .B1(U_afifo_n174), .B2(U_afifo_n207), .A(
        U_afifo_n206), .ZN(U_afifo_n26) );
  NAND2_X2 U_afifo_U255 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_30_), .ZN(
        U_afifo_n222) );
  OAI21_X2 U_afifo_U254 ( .B1(U_afifo_n174), .B2(U_afifo_n223), .A(
        U_afifo_n222), .ZN(U_afifo_n34) );
  NAND2_X2 U_afifo_U253 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_2_), .ZN(
        U_afifo_n188) );
  OAI21_X2 U_afifo_U252 ( .B1(U_afifo_n174), .B2(hwrite), .A(U_afifo_n188), 
        .ZN(U_afifo_n6) );
  NAND2_X2 U_afifo_U251 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_29_), .ZN(
        U_afifo_n220) );
  OAI21_X2 U_afifo_U250 ( .B1(U_afifo_n174), .B2(U_afifo_n221), .A(
        U_afifo_n220), .ZN(U_afifo_n33) );
  NAND2_X2 U_afifo_U249 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_28_), .ZN(
        U_afifo_n218) );
  OAI21_X2 U_afifo_U248 ( .B1(U_afifo_n174), .B2(U_afifo_n219), .A(
        U_afifo_n218), .ZN(U_afifo_n32) );
  NAND2_X2 U_afifo_U247 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_23_), .ZN(
        U_afifo_n208) );
  OAI21_X2 U_afifo_U246 ( .B1(U_afifo_n174), .B2(U_afifo_n209), .A(
        U_afifo_n208), .ZN(U_afifo_n27) );
  NAND2_X2 U_afifo_U245 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_21_), .ZN(
        U_afifo_n204) );
  OAI21_X2 U_afifo_U244 ( .B1(U_afifo_n174), .B2(U_afifo_n205), .A(
        U_afifo_n204), .ZN(U_afifo_n25) );
  NAND2_X2 U_afifo_U243 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_25_), .ZN(
        U_afifo_n212) );
  OAI21_X2 U_afifo_U242 ( .B1(U_afifo_n174), .B2(U_afifo_n213), .A(
        U_afifo_n212), .ZN(U_afifo_n29) );
  NAND2_X2 U_afifo_U241 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_24_), .ZN(
        U_afifo_n210) );
  OAI21_X2 U_afifo_U240 ( .B1(U_afifo_n174), .B2(U_afifo_n211), .A(
        U_afifo_n210), .ZN(U_afifo_n28) );
  NAND2_X2 U_afifo_U239 ( .A1(n47), .A2(m_af_data2_in[15]), .ZN(U_afifo_n195)
         );
  OAI21_X2 U_afifo_U238 ( .B1(n47), .B2(U_afifo_n162), .A(U_afifo_n195), .ZN(
        U_afifo_n19) );
  NAND2_X2 U_afifo_U237 ( .A1(n47), .A2(m_af_data2_in[14]), .ZN(U_afifo_n194)
         );
  OAI21_X2 U_afifo_U236 ( .B1(n47), .B2(U_afifo_n161), .A(U_afifo_n194), .ZN(
        U_afifo_n18) );
  NAND2_X2 U_afifo_U235 ( .A1(n47), .A2(m_af_data2_in[16]), .ZN(U_afifo_n196)
         );
  OAI21_X2 U_afifo_U234 ( .B1(n47), .B2(U_afifo_n163), .A(U_afifo_n196), .ZN(
        U_afifo_n20) );
  NAND2_X2 U_afifo_U231 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_36_), .ZN(
        U_afifo_n234) );
  OAI21_X2 U_afifo_U230 ( .B1(U_afifo_n176), .B2(U_afifo_n235), .A(
        U_afifo_n234), .ZN(U_afifo_n40) );
  NAND2_X2 U_afifo_U229 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_38_), .ZN(
        U_afifo_n238) );
  OAI21_X2 U_afifo_U228 ( .B1(U_afifo_n176), .B2(U_afifo_n239), .A(
        U_afifo_n238), .ZN(U_afifo_n42) );
  NAND2_X2 U_afifo_U227 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_42_), .ZN(
        U_afifo_n246) );
  OAI21_X2 U_afifo_U226 ( .B1(U_afifo_n176), .B2(U_ctl_n227), .A(U_afifo_n246), 
        .ZN(U_afifo_n46) );
  NAND2_X2 U_afifo_U225 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_43_), .ZN(
        U_afifo_n248) );
  OAI21_X2 U_afifo_U224 ( .B1(U_afifo_n176), .B2(U_ctl_n230), .A(U_afifo_n248), 
        .ZN(U_afifo_n47) );
  NAND2_X2 U_afifo_U223 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_34_), .ZN(
        U_afifo_n230) );
  OAI21_X2 U_afifo_U222 ( .B1(U_afifo_n176), .B2(U_afifo_n231), .A(
        U_afifo_n230), .ZN(U_afifo_n38) );
  NAND2_X2 U_afifo_U221 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_39_), .ZN(
        U_afifo_n240) );
  OAI21_X2 U_afifo_U220 ( .B1(U_afifo_n176), .B2(U_afifo_n241), .A(
        U_afifo_n240), .ZN(U_afifo_n43) );
  NAND2_X2 U_afifo_U219 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_41_), .ZN(
        U_afifo_n244) );
  OAI21_X2 U_afifo_U218 ( .B1(U_afifo_n176), .B2(U_afifo_n245), .A(
        U_afifo_n244), .ZN(U_afifo_n45) );
  NAND2_X2 U_afifo_U217 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_35_), .ZN(
        U_afifo_n232) );
  OAI21_X2 U_afifo_U216 ( .B1(U_afifo_n176), .B2(U_afifo_n233), .A(
        U_afifo_n232), .ZN(U_afifo_n39) );
  NAND2_X2 U_afifo_U215 ( .A1(U_afifo_n174), .A2(U_afifo_f_data2_40_), .ZN(
        U_afifo_n242) );
  OAI21_X2 U_afifo_U214 ( .B1(U_afifo_n176), .B2(U_afifo_n243), .A(
        U_afifo_n242), .ZN(U_afifo_n44) );
  NAND2_X2 U_afifo_U213 ( .A1(U_afifo_n176), .A2(U_afifo_f_data2_37_), .ZN(
        U_afifo_n236) );
  OAI21_X2 U_afifo_U212 ( .B1(U_afifo_n176), .B2(U_afifo_n237), .A(
        U_afifo_n236), .ZN(U_afifo_n41) );
  NAND2_X2 U_afifo_U211 ( .A1(m_af_data2_in[6]), .A2(n47), .ZN(U_afifo_n170)
         );
  NAND2_X2 U_afifo_U210 ( .A1(U_afifo_f_data2_6_), .A2(U_afifo_n176), .ZN(
        U_afifo_n171) );
  NAND2_X2 U_afifo_U209 ( .A1(U_afifo_n170), .A2(U_afifo_n171), .ZN(
        U_afifo_n155) );
  INV_X4 U_afifo_U208 ( .A(U_afifo_m_data_out_0_), .ZN(U_afifo_n256) );
  NOR3_X2 U_afifo_U207 ( .A1(m_af_dummy_req), .A2(U_afifo_m_empty), .A3(
        U_afifo_n256), .ZN(hiu_req[1]) );
  AOI21_X2 U_afifo_U206 ( .B1(U_afifo_m_afull), .B2(U_afifo_f_push2_pending), 
        .A(U_afifo_n151), .ZN(m_af_ready) );
  AOI22_X2 U_afifo_U205 ( .A1(m_af_data1_in_5_), .A2(U_afifo_n140), .B1(
        U_afifo_f_data2_5_), .B2(U_afifo_n54), .ZN(U_afifo_n179) );
  INV_X4 U_afifo_U204 ( .A(U_afifo_n179), .ZN(U_afifo_m_data_in[5]) );
  AOI22_X2 U_afifo_U203 ( .A1(m_af_data1_in_6_), .A2(U_afifo_n93), .B1(
        U_afifo_f_data2_6_), .B2(U_afifo_n54), .ZN(U_afifo_n180) );
  INV_X4 U_afifo_U202 ( .A(U_afifo_n180), .ZN(U_afifo_m_data_in[6]) );
  OAI21_X2 U_afifo_U201 ( .B1(U_afifo_m_aempty), .B2(U_afifo_n255), .A(
        U_afifo_n184), .ZN(U_afifo_n_new_req) );
  NAND2_X2 U_afifo_U200 ( .A1(U_afifo_n168), .A2(U_afifo_n167), .ZN(
        U_afifo_n169) );
  OAI21_X2 U_afifo_U199 ( .B1(U_afifo_n185), .B2(U_afifo_n156), .A(
        U_afifo_n169), .ZN(U_afifo_n65) );
  NOR3_X2 U_afifo_U198 ( .A1(m_af_dummy_req), .A2(U_afifo_m_empty), .A3(
        U_afifo_m_data_out_0_), .ZN(hiu_req[0]) );
  INV_X1 U_afifo_U197 ( .A(m_af_data1_in_0_), .ZN(U_afifo_n187) );
  INV_X1 U_afifo_U196 ( .A(miu_burst_done), .ZN(U_afifo_n255) );
  OAI21_X1 U_afifo_U195 ( .B1(miu_burst_done), .B2(U_afifo_m_empty), .A(
        U_afifo_n185), .ZN(U_afifo_n184) );
  INV_X4 U_afifo_U194 ( .A(U_afifo_n259), .ZN(m_af_dummy_req) );
  INV_X1 U_afifo_U189 ( .A(U_afifo_n54), .ZN(U_afifo_n147) );
  INV_X1 U_afifo_U184 ( .A(U_afifo_n54), .ZN(U_afifo_n140) );
  NAND2_X2 U_afifo_U182 ( .A1(U_afifo_n54), .A2(U_afifo_f_data2_42_), .ZN(
        U_afifo_n137) );
  INV_X1 U_afifo_U156 ( .A(U_afifo_n54), .ZN(U_afifo_n99) );
  INV_X1 U_afifo_U155 ( .A(U_afifo_n54), .ZN(U_afifo_n98) );
  INV_X1 U_afifo_U151 ( .A(U_afifo_n54), .ZN(U_afifo_n93) );
  NAND2_X2 U_afifo_U145 ( .A1(U_afifo_n54), .A2(U_afifo_f_data2_38_), .ZN(
        U_afifo_n84) );
  NAND2_X2 U_afifo_U139 ( .A1(U_afifo_n54), .A2(U_afifo_f_data2_32_), .ZN(
        U_afifo_n75) );
  NAND2_X1 U_afifo_U125 ( .A1(U_afifo_f_core_ready), .A2(
        U_afifo_f_push2_pending), .ZN(U_afifo_n183) );
  INV_X2 U_afifo_U123 ( .A(U_afifo_m_full), .ZN(U_afifo_n167) );
  INV_X1 U_afifo_U122 ( .A(U_afifo_m_data_out_49), .ZN(U_afifo_n257) );
  NAND2_X2 U_afifo_U121 ( .A1(miu_burst_done), .A2(U_afifo_n259), .ZN(
        U_afifo_m_pop_n) );
  OAI21_X1 U_afifo_U120 ( .B1(U_afifo_n255), .B2(U_afifo_n259), .A(
        U_afifo_n258), .ZN(U_afifo_n2) );
  INV_X1 U_afifo_U116 ( .A(U_afifo_n185), .ZN(U_afifo_n55) );
  AND2_X2 U_afifo_U112 ( .A1(U_afifo_n99), .A2(m_af_data1_in_3_), .ZN(
        U_afifo_m_data_in[3]) );
  NAND2_X2 U_afifo_U107 ( .A1(U_afifo_n147), .A2(haddr[28]), .ZN(U_afifo_n85)
         );
  AND2_X2 U_afifo_U103 ( .A1(U_afifo_n147), .A2(haddr[0]), .ZN(
        U_afifo_m_data_in[45]) );
  NAND2_X2 U_afifo_U96 ( .A1(U_afifo_n147), .A2(haddr[22]), .ZN(U_afifo_n76)
         );
  AND2_X2 U_afifo_U92 ( .A1(U_afifo_n140), .A2(haddr[1]), .ZN(
        U_afifo_m_data_in[46]) );
  AND2_X2 U_afifo_U91 ( .A1(m_af_data1_in_11_), .A2(U_afifo_n99), .ZN(
        U_afifo_m_data_in[11]) );
  AND2_X2 U_afifo_U89 ( .A1(m_af_data1_in_9_), .A2(U_afifo_n147), .ZN(
        U_afifo_m_data_in[9]) );
  NAND2_X2 U_afifo_U81 ( .A1(U_afifo_n85), .A2(U_afifo_n84), .ZN(
        U_afifo_m_data_in[38]) );
  NAND2_X2 U_afifo_U64 ( .A1(U_afifo_n76), .A2(U_afifo_n75), .ZN(
        U_afifo_m_data_in[32]) );
  NAND2_X2 U_afifo_U62 ( .A1(U_afifo_n138), .A2(U_afifo_n137), .ZN(
        U_afifo_m_data_in[42]) );
  AOI22_X2 U_afifo_U59 ( .A1(m_af_data2_in[7]), .A2(n47), .B1(
        U_afifo_f_data2_7_), .B2(U_afifo_n176), .ZN(U_afifo_n192) );
  INV_X2 U_afifo_U58 ( .A(haddr[17]), .ZN(U_afifo_n217) );
  INV_X2 U_afifo_U57 ( .A(haddr[11]), .ZN(U_afifo_n205) );
  INV_X2 U_afifo_U56 ( .A(haddr[18]), .ZN(U_afifo_n219) );
  INV_X2 U_afifo_U55 ( .A(haddr[12]), .ZN(U_afifo_n207) );
  INV_X2 U_afifo_U54 ( .A(haddr[13]), .ZN(U_afifo_n209) );
  INV_X2 U_afifo_U53 ( .A(haddr[9]), .ZN(U_afifo_n201) );
  INV_X2 U_afifo_U52 ( .A(haddr[15]), .ZN(U_afifo_n213) );
  INV_X2 U_afifo_U51 ( .A(haddr[16]), .ZN(U_afifo_n215) );
  INV_X2 U_afifo_U50 ( .A(haddr[14]), .ZN(U_afifo_n211) );
  INV_X2 U_afifo_U49 ( .A(haddr[10]), .ZN(U_afifo_n203) );
  INV_X2 U_afifo_U48 ( .A(haddr[30]), .ZN(U_afifo_n243) );
  INV_X2 U_afifo_U47 ( .A(haddr[31]), .ZN(U_afifo_n245) );
  INV_X2 U_afifo_U46 ( .A(haddr[26]), .ZN(U_afifo_n235) );
  INV_X2 U_afifo_U45 ( .A(haddr[27]), .ZN(U_afifo_n237) );
  INV_X2 U_afifo_U44 ( .A(haddr[28]), .ZN(U_afifo_n239) );
  INV_X2 U_afifo_U43 ( .A(haddr[29]), .ZN(U_afifo_n241) );
  INV_X2 U_afifo_U42 ( .A(haddr[23]), .ZN(U_afifo_n229) );
  INV_X2 U_afifo_U41 ( .A(haddr[21]), .ZN(U_afifo_n225) );
  INV_X2 U_afifo_U40 ( .A(haddr[24]), .ZN(U_afifo_n231) );
  INV_X2 U_afifo_U39 ( .A(haddr[20]), .ZN(U_afifo_n223) );
  INV_X2 U_afifo_U38 ( .A(haddr[22]), .ZN(U_afifo_n227) );
  INV_X2 U_afifo_U37 ( .A(haddr[25]), .ZN(U_afifo_n233) );
  INV_X2 U_afifo_U36 ( .A(haddr[19]), .ZN(U_afifo_n221) );
  OAI21_X1 U_afifo_U35 ( .B1(U_afifo_n255), .B2(U_afifo_n257), .A(
        U_afifo_f_clr_pers), .ZN(U_afifo_n258) );
  NAND2_X2 U_afifo_U33 ( .A1(U_afifo_n54), .A2(U_afifo_n183), .ZN(U_afifo_n185) );
  AND2_X2 U_afifo_U32 ( .A1(U_afifo_n54), .A2(U_afifo_f_data2_8_), .ZN(
        U_afifo_n152) );
  NAND2_X2 U_afifo_U29 ( .A1(U_afifo_n98), .A2(hsize[0]), .ZN(U_afifo_n138) );
  NOR2_X2 U_afifo_U28 ( .A1(U_afifo_n54), .A2(U_afifo_n157), .ZN(
        U_afifo_m_data_in[49]) );
  INV_X16 U_afifo_U26 ( .A(U_afifo_n178), .ZN(U_afifo_n54) );
  INV_X1 U_afifo_U25 ( .A(U_afifo_n49), .ZN(U_afifo_m_data_in[13]) );
  AOI22_X1 U_afifo_U24 ( .A1(U_afifo_n54), .A2(U_afifo_f_data2_13_), .B1(
        U_afifo_n178), .B2(m_af_data1_in_13_), .ZN(U_afifo_n49) );
  AOI22_X1 U_afifo_U22 ( .A1(haddr[3]), .A2(U_afifo_n147), .B1(
        U_afifo_f_data2_48_), .B2(U_afifo_n54), .ZN(U_afifo_n15) );
  INV_X1 U_afifo_U21 ( .A(U_afifo_n14), .ZN(U_afifo_m_data_in[47]) );
  AOI22_X1 U_afifo_U20 ( .A1(haddr[2]), .A2(U_afifo_n99), .B1(
        U_afifo_f_data2_47_), .B2(U_afifo_n54), .ZN(U_afifo_n14) );
  INV_X1 U_afifo_U19 ( .A(U_afifo_n13), .ZN(U_afifo_m_data_in[14]) );
  AOI22_X1 U_afifo_U18 ( .A1(haddr[4]), .A2(U_afifo_n98), .B1(
        U_afifo_f_data2_14_), .B2(U_afifo_n54), .ZN(U_afifo_n13) );
  INV_X1 U_afifo_U17 ( .A(U_afifo_n11), .ZN(U_afifo_m_data_in[15]) );
  AOI22_X1 U_afifo_U16 ( .A1(haddr[5]), .A2(U_afifo_n99), .B1(
        U_afifo_f_data2_15_), .B2(U_afifo_n54), .ZN(U_afifo_n11) );
  INV_X1 U_afifo_U15 ( .A(U_afifo_n10), .ZN(U_afifo_m_data_in[18]) );
  AOI22_X1 U_afifo_U14 ( .A1(haddr[8]), .A2(U_afifo_n98), .B1(
        U_afifo_f_data2_18_), .B2(U_afifo_n54), .ZN(U_afifo_n10) );
  INV_X1 U_afifo_U13 ( .A(U_afifo_n9), .ZN(U_afifo_m_data_in[43]) );
  AOI22_X1 U_afifo_U12 ( .A1(hsize[1]), .A2(U_afifo_n93), .B1(
        U_afifo_f_data2_43_), .B2(U_afifo_n54), .ZN(U_afifo_n9) );
  INV_X1 U_afifo_U11 ( .A(U_afifo_n7), .ZN(U_afifo_m_data_in[44]) );
  AOI22_X1 U_afifo_U10 ( .A1(hsize[2]), .A2(U_afifo_n140), .B1(
        U_afifo_f_data2_44_), .B2(U_afifo_n54), .ZN(U_afifo_n7) );
  INV_X1 U_afifo_U9 ( .A(U_afifo_n5), .ZN(U_afifo_m_data_in[0]) );
  AOI22_X1 U_afifo_U8 ( .A1(m_af_data1_in_0_), .A2(U_afifo_n140), .B1(
        U_afifo_f_data2_0_), .B2(U_afifo_n54), .ZN(U_afifo_n5) );
  INV_X1 U_afifo_U7 ( .A(U_afifo_n1), .ZN(U_afifo_m_data_in[4]) );
  AOI22_X2 U_afifo_U6 ( .A1(U_afifo_n54), .A2(U_afifo_f_data2_4_), .B1(
        U_afifo_n93), .B2(m_af_data1_in_4_), .ZN(U_afifo_n1) );
  AND2_X1 U_afifo_U5 ( .A1(U_afifo_n259), .A2(U_afifo_m_data_out_3), .ZN(
        hiu_wrap_burst) );
  INV_X4 U_afifo_U3 ( .A(m_af_push1_n), .ZN(U_afifo_n178) );
  DFFR_X2 U_afifo_f_data2_reg_8_ ( .D(U_afifo_n12), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_8_), .QN(U_afifo_n158) );
  DFFR_X2 U_afifo_f_data2_reg_12_ ( .D(U_afifo_n16), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_12_), .QN(U_afifo_n159) );
  DFFR_X2 U_afifo_f_data2_reg_13_ ( .D(U_afifo_n17), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_13_), .QN(U_afifo_n160) );
  DFFR_X2 U_afifo_f_data2_reg_47_ ( .D(U_afifo_n51), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_47_), .QN(U_afifo_n165) );
  DFFR_X2 U_afifo_f_data2_reg_48_ ( .D(U_afifo_n52), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_48_), .QN(U_afifo_n166) );
  DFFR_X2 U_afifo_f_data2_reg_4_ ( .D(U_afifo_n8), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_4_), .QN(U_afifo_n191) );
  DFFS_X2 U_afifo_f_data2_reg_7_ ( .D(U_afifo_n192), .CK(hclk), .SN(hresetn), 
        .QN(U_afifo_f_data2_7_) );
  DFFR_X1 U_afifo_f_new_req_reg ( .D(U_afifo_n_new_req), .CK(hclk), .RN(
        hresetn), .QN(m_af_new_req) );
  DFFS_X2 U_afifo_f_ready_reg ( .D(U_afifo_n65), .CK(hclk), .SN(hresetn), .QN(
        U_afifo_n151) );
  DFFR_X1 U_afifo_f_clr_pers_reg ( .D(U_afifo_n2), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_clr_pers), .QN(U_afifo_n153) );
  DFFR_X1 U_afifo_f_push2_pending_reg ( .D(U_afifo_n3), .CK(hclk), .RN(hresetn), .Q(U_afifo_f_push2_pending), .QN(U_afifo_n157) );
  DFFS_X2 U_afifo_f_core_ready_reg ( .D(U_afifo_n65), .CK(hclk), .SN(hresetn), 
        .Q(U_afifo_f_core_ready) );
  DFFR_X1 U_afifo_f_data2_reg_0_ ( .D(U_afifo_n4), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_0_) );
  DFFR_X1 U_afifo_f_data2_reg_2_ ( .D(U_afifo_n6), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_2_) );
  DFFR_X1 U_afifo_f_data2_reg_5_ ( .D(U_afifo_n154), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_5_) );
  DFFR_X1 U_afifo_f_data2_reg_6_ ( .D(U_afifo_n155), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_6_) );
  DFFR_X1 U_afifo_f_data2_reg_14_ ( .D(U_afifo_n18), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_14_), .QN(U_afifo_n161) );
  DFFR_X1 U_afifo_f_data2_reg_15_ ( .D(U_afifo_n19), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_15_), .QN(U_afifo_n162) );
  DFFR_X1 U_afifo_f_data2_reg_16_ ( .D(U_afifo_n20), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_16_), .QN(U_afifo_n163) );
  DFFR_X1 U_afifo_f_data2_reg_17_ ( .D(U_afifo_n21), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_17_), .QN(U_afifo_n164) );
  DFFR_X1 U_afifo_f_data2_reg_18_ ( .D(U_afifo_n22), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_18_) );
  DFFR_X1 U_afifo_f_data2_reg_19_ ( .D(U_afifo_n23), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_19_) );
  DFFR_X1 U_afifo_f_data2_reg_20_ ( .D(U_afifo_n24), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_20_) );
  DFFR_X1 U_afifo_f_data2_reg_21_ ( .D(U_afifo_n25), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_21_) );
  DFFR_X1 U_afifo_f_data2_reg_22_ ( .D(U_afifo_n26), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_22_) );
  DFFR_X1 U_afifo_f_data2_reg_23_ ( .D(U_afifo_n27), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_23_) );
  DFFR_X1 U_afifo_f_data2_reg_24_ ( .D(U_afifo_n28), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_24_) );
  DFFR_X1 U_afifo_f_data2_reg_25_ ( .D(U_afifo_n29), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_25_) );
  DFFR_X1 U_afifo_f_data2_reg_26_ ( .D(U_afifo_n30), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_26_) );
  DFFR_X1 U_afifo_f_data2_reg_27_ ( .D(U_afifo_n31), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_27_) );
  DFFR_X1 U_afifo_f_data2_reg_28_ ( .D(U_afifo_n32), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_28_) );
  DFFR_X1 U_afifo_f_data2_reg_29_ ( .D(U_afifo_n33), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_29_) );
  DFFR_X1 U_afifo_f_data2_reg_30_ ( .D(U_afifo_n34), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_30_) );
  DFFR_X1 U_afifo_f_data2_reg_31_ ( .D(U_afifo_n35), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_31_) );
  DFFR_X1 U_afifo_f_data2_reg_32_ ( .D(U_afifo_n36), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_32_) );
  DFFR_X1 U_afifo_f_data2_reg_33_ ( .D(U_afifo_n37), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_33_) );
  DFFR_X1 U_afifo_f_data2_reg_34_ ( .D(U_afifo_n38), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_34_) );
  DFFR_X1 U_afifo_f_data2_reg_35_ ( .D(U_afifo_n39), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_35_) );
  DFFR_X1 U_afifo_f_data2_reg_36_ ( .D(U_afifo_n40), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_36_) );
  DFFR_X1 U_afifo_f_data2_reg_37_ ( .D(U_afifo_n41), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_37_) );
  DFFR_X1 U_afifo_f_data2_reg_38_ ( .D(U_afifo_n42), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_38_) );
  DFFR_X1 U_afifo_f_data2_reg_39_ ( .D(U_afifo_n43), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_39_) );
  DFFR_X1 U_afifo_f_data2_reg_40_ ( .D(U_afifo_n44), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_40_) );
  DFFR_X1 U_afifo_f_data2_reg_41_ ( .D(U_afifo_n45), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_41_) );
  DFFR_X1 U_afifo_f_data2_reg_42_ ( .D(U_afifo_n46), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_42_) );
  DFFR_X1 U_afifo_f_data2_reg_43_ ( .D(U_afifo_n47), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_43_) );
  DFFR_X1 U_afifo_f_data2_reg_44_ ( .D(U_afifo_n48), .CK(hclk), .RN(hresetn), 
        .Q(U_afifo_f_data2_44_) );
  OAI221_X1 U_dfifo_U26 ( .B1(miu_pop_n), .B2(U_dfifo_f_1st_half), .C1(
        U_ctl_n384), .C2(U_dfifo_n2), .A(U_dfifo_m_data_out_1_), .ZN(
        U_dfifo_n3) );
  MUX2_X2 U_dfifo_U25 ( .A(hiu_data[24]), .B(U_dfifo_m_btm_data[8]), .S(
        U_dfifo_n4), .Z(hiu_data[8]) );
  MUX2_X2 U_dfifo_U24 ( .A(hiu_data[16]), .B(U_dfifo_m_btm_data[0]), .S(
        U_dfifo_n4), .Z(hiu_data[0]) );
  MUX2_X2 U_dfifo_U23 ( .A(hiu_data[25]), .B(U_dfifo_m_btm_data[9]), .S(
        U_dfifo_n4), .Z(hiu_data[9]) );
  MUX2_X2 U_dfifo_U22 ( .A(hiu_data[17]), .B(U_dfifo_m_btm_data[1]), .S(
        U_dfifo_n4), .Z(hiu_data[1]) );
  MUX2_X2 U_dfifo_U21 ( .A(hiu_data[26]), .B(U_dfifo_m_btm_data[10]), .S(
        U_dfifo_n4), .Z(hiu_data[10]) );
  MUX2_X2 U_dfifo_U20 ( .A(hiu_data[18]), .B(U_dfifo_m_btm_data[2]), .S(
        U_dfifo_n4), .Z(hiu_data[2]) );
  MUX2_X2 U_dfifo_U19 ( .A(hiu_data[28]), .B(U_dfifo_m_btm_data[12]), .S(
        U_dfifo_n4), .Z(hiu_data[12]) );
  MUX2_X2 U_dfifo_U18 ( .A(hiu_data[20]), .B(U_dfifo_m_btm_data[4]), .S(
        U_dfifo_n4), .Z(hiu_data[4]) );
  MUX2_X2 U_dfifo_U17 ( .A(hiu_data[27]), .B(U_dfifo_m_btm_data[11]), .S(
        U_dfifo_n4), .Z(hiu_data[11]) );
  MUX2_X2 U_dfifo_U16 ( .A(hiu_data[19]), .B(U_dfifo_m_btm_data[3]), .S(
        U_dfifo_n4), .Z(hiu_data[3]) );
  MUX2_X2 U_dfifo_U15 ( .A(hiu_data[29]), .B(U_dfifo_m_btm_data[13]), .S(
        U_dfifo_n4), .Z(hiu_data[13]) );
  MUX2_X2 U_dfifo_U14 ( .A(hiu_data[21]), .B(U_dfifo_m_btm_data[5]), .S(
        U_dfifo_n4), .Z(hiu_data[5]) );
  MUX2_X2 U_dfifo_U13 ( .A(hiu_data[31]), .B(U_dfifo_m_btm_data[15]), .S(
        U_dfifo_n4), .Z(hiu_data[15]) );
  MUX2_X2 U_dfifo_U12 ( .A(hiu_data[23]), .B(U_dfifo_m_btm_data[7]), .S(
        U_dfifo_n4), .Z(hiu_data[7]) );
  MUX2_X2 U_dfifo_U11 ( .A(hiu_data[30]), .B(U_dfifo_m_btm_data[14]), .S(
        U_dfifo_n4), .Z(hiu_data[14]) );
  MUX2_X2 U_dfifo_U10 ( .A(hiu_data[22]), .B(U_dfifo_m_btm_data[6]), .S(
        U_dfifo_n4), .Z(hiu_data[6]) );
  NAND2_X2 U_dfifo_U8 ( .A1(U_dfifo_m_data_out_1_), .A2(U_dfifo_n2), .ZN(
        U_dfifo_n4) );
  AOI21_X2 U_dfifo_U7 ( .B1(U_dfifo_f_1st_half), .B2(U_dfifo_m_data_out_1_), 
        .A(miu_pop_n), .ZN(U_dfifo_n5) );
  AND2_X2 U_dfifo_U6 ( .A1(U_dfifo_n5), .A2(U_dfifo_m_data_out_0_), .ZN(
        m_df_wr_term) );
  AOI21_X2 U_dfifo_U5 ( .B1(U_dfifo_m_afull), .B2(m_df_push_n), .A(
        U_dfifo_m_full), .ZN(m_df_ready) );
  DFFS_X2 U_dfifo_f_1st_half_reg ( .D(U_dfifo_n3), .CK(hclk), .SN(hresetn), 
        .Q(U_dfifo_f_1st_half), .QN(U_dfifo_n2) );
  INV_X4 U_rbuf_U215 ( .A(U_rbuf_n161), .ZN(U_rbuf_n177) );
  AND3_X4 U_rbuf_U214 ( .A1(n48), .A2(m_two_to_one), .A3(U_rbuf_n160), .ZN(
        U_rbuf_n16) );
  INV_X4 U_rbuf_U212 ( .A(U_rbuf_n198), .ZN(U_rbuf_n196) );
  INV_X4 U_rbuf_U211 ( .A(U_rbuf_n143), .ZN(U_rbuf_n119) );
  INV_X4 U_rbuf_U210 ( .A(U_rbuf_n119), .ZN(U_rbuf_n117) );
  NOR2_X2 U_rbuf_U208 ( .A1(U_ctl_n324), .A2(U_rbuf_n17), .ZN(U_rbuf_n148) );
  NOR2_X2 U_rbuf_U207 ( .A1(miu_push_n), .A2(U_rbuf_n148), .ZN(U_rbuf_n154) );
  NAND2_X2 U_rbuf_U206 ( .A1(m_rb_pop_n), .A2(U_rbuf_n154), .ZN(U_rbuf_n151)
         );
  INV_X4 U_rbuf_U205 ( .A(U_rbuf_n151), .ZN(m_rb_overflow) );
  NAND2_X2 U_rbuf_U204 ( .A1(m_double), .A2(U_rbuf_n120), .ZN(U_rbuf_n125) );
  NAND2_X2 U_rbuf_U203 ( .A1(U_rbuf_n125), .A2(n48), .ZN(U_rbuf_n126) );
  NAND2_X2 U_rbuf_U202 ( .A1(U_rbuf_n146), .A2(U_rbuf_n126), .ZN(U_rbuf_n143)
         );
  NAND2_X2 U_rbuf_U201 ( .A1(miu_data[1]), .A2(U_rbuf_n118), .ZN(U_rbuf_n128)
         );
  OAI21_X2 U_rbuf_U200 ( .B1(U_rbuf_n118), .B2(U_rbuf_n19), .A(U_rbuf_n128), 
        .ZN(hrdata[1]) );
  NAND2_X2 U_rbuf_U199 ( .A1(miu_data[9]), .A2(U_rbuf_n118), .ZN(U_rbuf_n136)
         );
  OAI21_X2 U_rbuf_U198 ( .B1(U_rbuf_n117), .B2(U_rbuf_n27), .A(U_rbuf_n136), 
        .ZN(hrdata[9]) );
  NAND2_X2 U_rbuf_U197 ( .A1(miu_data[3]), .A2(U_rbuf_n118), .ZN(U_rbuf_n130)
         );
  OAI21_X2 U_rbuf_U196 ( .B1(U_rbuf_n118), .B2(U_rbuf_n21), .A(U_rbuf_n130), 
        .ZN(hrdata[3]) );
  NAND2_X2 U_rbuf_U195 ( .A1(miu_data[5]), .A2(U_rbuf_n118), .ZN(U_rbuf_n132)
         );
  OAI21_X2 U_rbuf_U194 ( .B1(U_rbuf_n117), .B2(U_rbuf_n23), .A(U_rbuf_n132), 
        .ZN(hrdata[5]) );
  NAND2_X2 U_rbuf_U193 ( .A1(miu_data[7]), .A2(U_rbuf_n118), .ZN(U_rbuf_n134)
         );
  OAI21_X2 U_rbuf_U192 ( .B1(U_rbuf_n117), .B2(U_rbuf_n25), .A(U_rbuf_n134), 
        .ZN(hrdata[7]) );
  NAND2_X2 U_rbuf_U191 ( .A1(m_double), .A2(big_endian), .ZN(U_rbuf_n160) );
  NAND2_X2 U_rbuf_U188 ( .A1(miu_data[29]), .A2(U_rbuf_n6), .ZN(U_rbuf_n39) );
  NAND2_X2 U_rbuf_U187 ( .A1(miu_data[12]), .A2(U_rbuf_n118), .ZN(U_rbuf_n139)
         );
  OAI21_X2 U_rbuf_U186 ( .B1(U_rbuf_n117), .B2(U_rbuf_n30), .A(U_rbuf_n139), 
        .ZN(hrdata[12]) );
  NAND2_X2 U_rbuf_U185 ( .A1(miu_data[8]), .A2(U_rbuf_n118), .ZN(U_rbuf_n135)
         );
  OAI21_X2 U_rbuf_U184 ( .B1(U_rbuf_n117), .B2(U_rbuf_n26), .A(U_rbuf_n135), 
        .ZN(hrdata[8]) );
  NAND2_X2 U_rbuf_U183 ( .A1(miu_data[6]), .A2(U_rbuf_n118), .ZN(U_rbuf_n133)
         );
  OAI21_X2 U_rbuf_U182 ( .B1(U_rbuf_n117), .B2(U_rbuf_n24), .A(U_rbuf_n133), 
        .ZN(hrdata[6]) );
  NAND2_X2 U_rbuf_U181 ( .A1(miu_data[11]), .A2(U_rbuf_n118), .ZN(U_rbuf_n138)
         );
  OAI21_X2 U_rbuf_U180 ( .B1(U_rbuf_n117), .B2(U_rbuf_n29), .A(U_rbuf_n138), 
        .ZN(hrdata[11]) );
  NAND2_X2 U_rbuf_U179 ( .A1(miu_data[15]), .A2(U_rbuf_n118), .ZN(U_rbuf_n142)
         );
  NAND2_X2 U_rbuf_U178 ( .A1(miu_data[4]), .A2(U_rbuf_n118), .ZN(U_rbuf_n131)
         );
  OAI21_X2 U_rbuf_U177 ( .B1(U_rbuf_n117), .B2(U_rbuf_n22), .A(U_rbuf_n131), 
        .ZN(hrdata[4]) );
  NAND2_X2 U_rbuf_U176 ( .A1(miu_data[2]), .A2(U_rbuf_n118), .ZN(U_rbuf_n129)
         );
  OAI21_X2 U_rbuf_U175 ( .B1(U_rbuf_n118), .B2(U_rbuf_n20), .A(U_rbuf_n129), 
        .ZN(hrdata[2]) );
  NAND2_X2 U_rbuf_U174 ( .A1(miu_data[0]), .A2(U_rbuf_n118), .ZN(U_rbuf_n127)
         );
  OAI21_X2 U_rbuf_U173 ( .B1(U_rbuf_n118), .B2(U_rbuf_n18), .A(U_rbuf_n127), 
        .ZN(hrdata[0]) );
  NAND2_X2 U_rbuf_U172 ( .A1(miu_data[13]), .A2(U_rbuf_n118), .ZN(U_rbuf_n140)
         );
  NAND2_X2 U_rbuf_U171 ( .A1(miu_data[14]), .A2(U_rbuf_n118), .ZN(U_rbuf_n141)
         );
  OAI21_X2 U_rbuf_U170 ( .B1(U_rbuf_n117), .B2(U_rbuf_n33), .A(U_rbuf_n141), 
        .ZN(hrdata[14]) );
  NAND2_X2 U_rbuf_U169 ( .A1(miu_data[25]), .A2(U_rbuf_n6), .ZN(U_rbuf_n45) );
  NAND2_X2 U_rbuf_U168 ( .A1(miu_data[9]), .A2(U_rbuf_n16), .ZN(U_rbuf_n44) );
  NAND3_X2 U_rbuf_U167 ( .A1(U_rbuf_n45), .A2(U_rbuf_n44), .A3(U_rbuf_n43), 
        .ZN(hrdata[25]) );
  NAND2_X2 U_rbuf_U166 ( .A1(miu_data[17]), .A2(U_rbuf_n6), .ZN(U_rbuf_n54) );
  NAND2_X2 U_rbuf_U165 ( .A1(miu_data[1]), .A2(U_rbuf_n16), .ZN(U_rbuf_n53) );
  NAND3_X2 U_rbuf_U164 ( .A1(U_rbuf_n54), .A2(U_rbuf_n53), .A3(U_rbuf_n52), 
        .ZN(hrdata[17]) );
  NAND2_X2 U_rbuf_U163 ( .A1(miu_data[19]), .A2(U_rbuf_n6), .ZN(U_rbuf_n51) );
  NAND2_X2 U_rbuf_U162 ( .A1(miu_data[3]), .A2(U_rbuf_n16), .ZN(U_rbuf_n50) );
  NAND3_X2 U_rbuf_U161 ( .A1(U_rbuf_n51), .A2(U_rbuf_n50), .A3(U_rbuf_n49), 
        .ZN(hrdata[19]) );
  NAND2_X2 U_rbuf_U160 ( .A1(miu_data[21]), .A2(U_rbuf_n6), .ZN(U_rbuf_n48) );
  NAND2_X2 U_rbuf_U159 ( .A1(miu_data[5]), .A2(U_rbuf_n16), .ZN(U_rbuf_n47) );
  NAND3_X2 U_rbuf_U158 ( .A1(U_rbuf_n48), .A2(U_rbuf_n47), .A3(U_rbuf_n46), 
        .ZN(hrdata[21]) );
  NAND2_X2 U_rbuf_U157 ( .A1(miu_data[23]), .A2(U_rbuf_n6), .ZN(U_rbuf_n42) );
  NAND2_X2 U_rbuf_U156 ( .A1(miu_data[7]), .A2(U_rbuf_n16), .ZN(U_rbuf_n41) );
  NAND3_X2 U_rbuf_U155 ( .A1(U_rbuf_n42), .A2(U_rbuf_n41), .A3(U_rbuf_n40), 
        .ZN(hrdata[23]) );
  NAND2_X2 U_rbuf_U154 ( .A1(miu_data[10]), .A2(U_rbuf_n118), .ZN(U_rbuf_n137)
         );
  NOR2_X2 U_rbuf_U153 ( .A1(U_rbuf_n154), .A2(U_rbuf_f_rbuf_state_1_), .ZN(
        U_rbuf_n149) );
  NAND2_X2 U_rbuf_U152 ( .A1(U_rbuf_n149), .A2(U_rbuf_f_rbuf_state_0_), .ZN(
        m_rb_ready) );
  NAND2_X2 U_rbuf_U151 ( .A1(miu_data[16]), .A2(U_rbuf_n6), .ZN(U_rbuf_n116)
         );
  NAND2_X2 U_rbuf_U150 ( .A1(miu_data[0]), .A2(U_rbuf_n16), .ZN(U_rbuf_n114)
         );
  NAND3_X2 U_rbuf_U149 ( .A1(U_rbuf_n116), .A2(U_rbuf_n115), .A3(U_rbuf_n114), 
        .ZN(hrdata[16]) );
  NAND2_X2 U_rbuf_U148 ( .A1(miu_data[18]), .A2(U_rbuf_n6), .ZN(U_rbuf_n113)
         );
  NAND2_X2 U_rbuf_U147 ( .A1(miu_data[2]), .A2(U_rbuf_n16), .ZN(U_rbuf_n111)
         );
  NAND3_X2 U_rbuf_U146 ( .A1(U_rbuf_n113), .A2(U_rbuf_n112), .A3(U_rbuf_n111), 
        .ZN(hrdata[18]) );
  NAND2_X2 U_rbuf_U145 ( .A1(miu_data[27]), .A2(U_rbuf_n6), .ZN(U_rbuf_n101)
         );
  NAND2_X2 U_rbuf_U144 ( .A1(miu_data[11]), .A2(U_rbuf_n16), .ZN(U_rbuf_n99)
         );
  NAND3_X2 U_rbuf_U143 ( .A1(U_rbuf_n101), .A2(U_rbuf_n100), .A3(U_rbuf_n99), 
        .ZN(hrdata[27]) );
  NAND2_X2 U_rbuf_U142 ( .A1(miu_data[28]), .A2(U_rbuf_n6), .ZN(U_rbuf_n98) );
  NAND2_X2 U_rbuf_U141 ( .A1(miu_data[12]), .A2(U_rbuf_n16), .ZN(U_rbuf_n96)
         );
  NAND3_X2 U_rbuf_U140 ( .A1(U_rbuf_n98), .A2(U_rbuf_n97), .A3(U_rbuf_n96), 
        .ZN(hrdata[28]) );
  NAND2_X2 U_rbuf_U139 ( .A1(miu_data[24]), .A2(U_rbuf_n6), .ZN(U_rbuf_n104)
         );
  NAND2_X2 U_rbuf_U138 ( .A1(miu_data[8]), .A2(U_rbuf_n16), .ZN(U_rbuf_n102)
         );
  NAND3_X2 U_rbuf_U137 ( .A1(U_rbuf_n104), .A2(U_rbuf_n103), .A3(U_rbuf_n102), 
        .ZN(hrdata[24]) );
  NAND2_X2 U_rbuf_U136 ( .A1(miu_data[31]), .A2(U_rbuf_n6), .ZN(U_rbuf_n92) );
  NAND2_X2 U_rbuf_U135 ( .A1(miu_data[15]), .A2(U_rbuf_n16), .ZN(U_rbuf_n90)
         );
  NAND3_X2 U_rbuf_U134 ( .A1(U_rbuf_n92), .A2(U_rbuf_n91), .A3(U_rbuf_n90), 
        .ZN(hrdata[31]) );
  NAND2_X2 U_rbuf_U133 ( .A1(miu_data[20]), .A2(U_rbuf_n6), .ZN(U_rbuf_n110)
         );
  NAND2_X2 U_rbuf_U132 ( .A1(miu_data[4]), .A2(U_rbuf_n16), .ZN(U_rbuf_n108)
         );
  NAND3_X2 U_rbuf_U131 ( .A1(U_rbuf_n110), .A2(U_rbuf_n109), .A3(U_rbuf_n108), 
        .ZN(hrdata[20]) );
  NAND2_X2 U_rbuf_U130 ( .A1(miu_data[30]), .A2(U_rbuf_n6), .ZN(U_rbuf_n95) );
  NAND2_X2 U_rbuf_U129 ( .A1(miu_data[14]), .A2(U_rbuf_n16), .ZN(U_rbuf_n93)
         );
  NAND3_X2 U_rbuf_U128 ( .A1(U_rbuf_n95), .A2(U_rbuf_n94), .A3(U_rbuf_n93), 
        .ZN(hrdata[30]) );
  NAND2_X2 U_rbuf_U127 ( .A1(miu_data[22]), .A2(U_rbuf_n6), .ZN(U_rbuf_n107)
         );
  NAND2_X2 U_rbuf_U126 ( .A1(miu_data[6]), .A2(U_rbuf_n16), .ZN(U_rbuf_n105)
         );
  NAND3_X2 U_rbuf_U125 ( .A1(U_rbuf_n107), .A2(U_rbuf_n106), .A3(U_rbuf_n105), 
        .ZN(hrdata[22]) );
  NOR4_X2 U_rbuf_U124 ( .A1(m_rb_start), .A2(m_rb_done), .A3(U_ctl_n397), .A4(
        U_rbuf_n152), .ZN(U_rbuf_n87) );
  AOI21_X2 U_rbuf_U123 ( .B1(U_rbuf_n157), .B2(U_rbuf_f_rbuf_state_0_), .A(
        U_rbuf_n156), .ZN(U_rbuf_n158) );
  INV_X4 U_rbuf_U122 ( .A(m_rb_start), .ZN(U_rbuf_n159) );
  OAI211_X2 U_rbuf_U121 ( .C1(m_rb_done), .C2(U_rbuf_n158), .A(U_rbuf_n159), 
        .B(m_rb_ready), .ZN(U_rbuf_n88) );
  NAND2_X1 U_rbuf_U119 ( .A1(m_double), .A2(m_two_to_one), .ZN(U_rbuf_n123) );
  OAI21_X2 U_rbuf_U117 ( .B1(U_rbuf_n181), .B2(U_rbuf_n180), .A(U_rbuf_n162), 
        .ZN(U_rbuf_n55) );
  OAI21_X2 U_rbuf_U116 ( .B1(U_rbuf_n180), .B2(U_rbuf_n192), .A(U_rbuf_n173), 
        .ZN(U_rbuf_n66) );
  AOI22_X2 U_rbuf_U114 ( .A1(miu_data[23]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_7_), .B2(U_rbuf_n177), .ZN(U_rbuf_n169) );
  OAI21_X2 U_rbuf_U113 ( .B1(U_rbuf_n180), .B2(U_rbuf_n188), .A(U_rbuf_n169), 
        .ZN(U_rbuf_n62) );
  OAI21_X2 U_rbuf_U111 ( .B1(U_rbuf_n180), .B2(U_rbuf_n191), .A(U_rbuf_n172), 
        .ZN(U_rbuf_n65) );
  AOI22_X2 U_rbuf_U109 ( .A1(miu_data[19]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_3_), .B2(U_rbuf_n177), .ZN(U_rbuf_n165) );
  OAI21_X2 U_rbuf_U108 ( .B1(U_rbuf_n180), .B2(U_rbuf_n184), .A(U_rbuf_n165), 
        .ZN(U_rbuf_n58) );
  OAI21_X2 U_rbuf_U107 ( .B1(U_rbuf_n180), .B2(U_rbuf_n195), .A(U_rbuf_n176), 
        .ZN(U_rbuf_n69) );
  AOI22_X2 U_rbuf_U106 ( .A1(miu_data[29]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_13_), .B2(U_rbuf_n177), .ZN(U_rbuf_n175) );
  OAI21_X2 U_rbuf_U105 ( .B1(U_rbuf_n180), .B2(U_rbuf_n194), .A(U_rbuf_n175), 
        .ZN(U_rbuf_n68) );
  OAI21_X2 U_rbuf_U104 ( .B1(U_rbuf_n180), .B2(U_rbuf_n189), .A(U_rbuf_n170), 
        .ZN(U_rbuf_n63) );
  OAI21_X2 U_rbuf_U102 ( .B1(U_rbuf_n180), .B2(U_rbuf_n190), .A(U_rbuf_n171), 
        .ZN(U_rbuf_n64) );
  AOI22_X2 U_rbuf_U101 ( .A1(miu_data[31]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_15_), .B2(U_rbuf_n177), .ZN(U_rbuf_n179) );
  OAI21_X2 U_rbuf_U100 ( .B1(U_rbuf_n180), .B2(U_rbuf_n197), .A(U_rbuf_n179), 
        .ZN(U_rbuf_n70) );
  OAI21_X2 U_rbuf_U99 ( .B1(U_rbuf_n180), .B2(U_rbuf_n185), .A(U_rbuf_n166), 
        .ZN(U_rbuf_n59) );
  AOI22_X2 U_rbuf_U98 ( .A1(miu_data[18]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_2_), .B2(U_rbuf_n177), .ZN(U_rbuf_n164) );
  OAI21_X2 U_rbuf_U97 ( .B1(U_rbuf_n180), .B2(U_rbuf_n183), .A(U_rbuf_n164), 
        .ZN(U_rbuf_n57) );
  AOI22_X2 U_rbuf_U95 ( .A1(miu_data[17]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_1_), .B2(U_rbuf_n177), .ZN(U_rbuf_n163) );
  OAI21_X2 U_rbuf_U94 ( .B1(U_rbuf_n180), .B2(U_rbuf_n182), .A(U_rbuf_n163), 
        .ZN(U_rbuf_n56) );
  OAI21_X2 U_rbuf_U92 ( .B1(U_rbuf_n180), .B2(U_rbuf_n186), .A(U_rbuf_n167), 
        .ZN(U_rbuf_n60) );
  AOI22_X2 U_rbuf_U90 ( .A1(miu_data[28]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_12_), .B2(U_rbuf_n177), .ZN(U_rbuf_n174) );
  OAI21_X2 U_rbuf_U89 ( .B1(U_rbuf_n180), .B2(U_rbuf_n193), .A(U_rbuf_n174), 
        .ZN(U_rbuf_n67) );
  AOI22_X2 U_rbuf_U87 ( .A1(miu_data[22]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_6_), .B2(U_rbuf_n177), .ZN(U_rbuf_n168) );
  OAI21_X2 U_rbuf_U86 ( .B1(U_rbuf_n180), .B2(U_rbuf_n187), .A(U_rbuf_n168), 
        .ZN(U_rbuf_n61) );
  NOR2_X2 U_rbuf_U85 ( .A1(U_rbuf_n123), .A2(U_rbuf_n34), .ZN(U_rbuf_n124) );
  AOI22_X2 U_rbuf_U84 ( .A1(U_rbuf_n198), .A2(U_rbuf_n193), .B1(U_rbuf_n30), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n83) );
  AOI22_X2 U_rbuf_U83 ( .A1(U_rbuf_n198), .A2(U_rbuf_n194), .B1(U_rbuf_n31), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n84) );
  AOI22_X2 U_rbuf_U82 ( .A1(U_rbuf_n198), .A2(U_rbuf_n191), .B1(U_rbuf_n28), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n81) );
  AOI22_X2 U_rbuf_U81 ( .A1(U_rbuf_n198), .A2(U_rbuf_n195), .B1(U_rbuf_n33), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n85) );
  AOI22_X2 U_rbuf_U80 ( .A1(U_rbuf_n198), .A2(U_rbuf_n181), .B1(U_rbuf_n18), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n71) );
  AOI22_X2 U_rbuf_U79 ( .A1(U_rbuf_n198), .A2(U_rbuf_n197), .B1(U_rbuf_n32), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n86) );
  AOI22_X2 U_rbuf_U78 ( .A1(U_rbuf_n198), .A2(U_rbuf_n184), .B1(U_rbuf_n21), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n74) );
  AOI22_X2 U_rbuf_U77 ( .A1(U_rbuf_n198), .A2(U_rbuf_n189), .B1(U_rbuf_n26), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n79) );
  AOI22_X2 U_rbuf_U76 ( .A1(U_rbuf_n198), .A2(U_rbuf_n183), .B1(U_rbuf_n20), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n73) );
  AOI22_X2 U_rbuf_U75 ( .A1(U_rbuf_n198), .A2(U_rbuf_n190), .B1(U_rbuf_n27), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n80) );
  AOI22_X2 U_rbuf_U74 ( .A1(U_rbuf_n198), .A2(U_rbuf_n182), .B1(U_rbuf_n19), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n72) );
  AOI22_X2 U_rbuf_U73 ( .A1(U_rbuf_n198), .A2(U_rbuf_n188), .B1(U_rbuf_n25), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n78) );
  AOI22_X2 U_rbuf_U72 ( .A1(U_rbuf_n198), .A2(U_rbuf_n187), .B1(U_rbuf_n24), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n77) );
  AOI22_X2 U_rbuf_U71 ( .A1(U_rbuf_n198), .A2(U_rbuf_n185), .B1(U_rbuf_n22), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n75) );
  AOI22_X2 U_rbuf_U70 ( .A1(U_rbuf_n198), .A2(U_rbuf_n186), .B1(U_rbuf_n23), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n76) );
  AOI22_X2 U_rbuf_U69 ( .A1(U_rbuf_n198), .A2(U_rbuf_n192), .B1(U_rbuf_n29), 
        .B2(U_rbuf_n196), .ZN(U_rbuf_n82) );
  INV_X4 U_rbuf_U68 ( .A(big_endian), .ZN(U_rbuf_n120) );
  NOR2_X2 U_rbuf_U67 ( .A1(miu_push_n), .A2(U_rbuf_n124), .ZN(U_rbuf_n198) );
  NAND2_X1 U_rbuf_U66 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_7_), .ZN(
        U_rbuf_n40) );
  NAND2_X1 U_rbuf_U65 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_5_), .ZN(
        U_rbuf_n46) );
  NAND2_X1 U_rbuf_U64 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_3_), .ZN(
        U_rbuf_n49) );
  NAND2_X1 U_rbuf_U63 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_1_), .ZN(
        U_rbuf_n52) );
  NAND2_X1 U_rbuf_U62 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_9_), .ZN(
        U_rbuf_n43) );
  NAND2_X1 U_rbuf_U61 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_6_), .ZN(
        U_rbuf_n106) );
  NAND2_X1 U_rbuf_U60 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_14_), .ZN(
        U_rbuf_n94) );
  NAND2_X1 U_rbuf_U59 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_4_), .ZN(
        U_rbuf_n109) );
  NAND2_X1 U_rbuf_U58 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_15_), .ZN(
        U_rbuf_n91) );
  NAND2_X1 U_rbuf_U57 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_8_), .ZN(
        U_rbuf_n103) );
  NAND2_X1 U_rbuf_U56 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_12_), .ZN(
        U_rbuf_n97) );
  NAND2_X1 U_rbuf_U55 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_11_), .ZN(
        U_rbuf_n100) );
  NAND2_X1 U_rbuf_U54 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_2_), .ZN(
        U_rbuf_n112) );
  NAND2_X1 U_rbuf_U53 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_0_), .ZN(
        U_rbuf_n115) );
  NAND2_X2 U_rbuf_U52 ( .A1(U_rbuf_n15), .A2(U_rbuf_n142), .ZN(hrdata[15]) );
  NAND3_X2 U_rbuf_U51 ( .A1(U_rbuf_n9), .A2(U_rbuf_n8), .A3(U_rbuf_n7), .ZN(
        hrdata[26]) );
  NAND2_X2 U_rbuf_U50 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_10_), .ZN(
        U_rbuf_n7) );
  NAND2_X2 U_rbuf_U49 ( .A1(miu_data[10]), .A2(U_rbuf_n16), .ZN(U_rbuf_n8) );
  NAND2_X2 U_rbuf_U48 ( .A1(miu_data[26]), .A2(U_rbuf_n6), .ZN(U_rbuf_n9) );
  NAND2_X2 U_rbuf_U47 ( .A1(m_two_to_one), .A2(U_rbuf_n161), .ZN(U_rbuf_n180)
         );
  NOR2_X2 U_rbuf_U46 ( .A1(miu_push_n), .A2(m_two_to_one), .ZN(U_rbuf_n178) );
  XOR2_X1 U_rbuf_U44 ( .A(U_rbuf_f_1st_half), .B(big_endian), .Z(U_rbuf_n34)
         );
  NOR2_X1 U_rbuf_U41 ( .A1(U_ctl_n397), .A2(U_rbuf_f_rbuf_state_1_), .ZN(
        U_rbuf_n155) );
  INV_X1 U_rbuf_U40 ( .A(miu_data[2]), .ZN(U_rbuf_n183) );
  INV_X1 U_rbuf_U39 ( .A(miu_data[11]), .ZN(U_rbuf_n192) );
  INV_X1 U_rbuf_U38 ( .A(miu_data[14]), .ZN(U_rbuf_n195) );
  INV_X1 U_rbuf_U37 ( .A(miu_data[15]), .ZN(U_rbuf_n197) );
  OAI21_X1 U_rbuf_U36 ( .B1(U_rbuf_n155), .B2(m_rb_pop_n), .A(U_rbuf_n154), 
        .ZN(U_rbuf_n157) );
  INV_X1 U_rbuf_U35 ( .A(miu_data[8]), .ZN(U_rbuf_n189) );
  INV_X1 U_rbuf_U34 ( .A(miu_data[4]), .ZN(U_rbuf_n185) );
  INV_X1 U_rbuf_U33 ( .A(miu_data[13]), .ZN(U_rbuf_n194) );
  INV_X1 U_rbuf_U32 ( .A(U_rbuf_n149), .ZN(U_rbuf_n150) );
  OR2_X2 U_rbuf_U31 ( .A1(U_rbuf_n117), .A2(U_rbuf_n32), .ZN(U_rbuf_n15) );
  NOR3_X1 U_rbuf_U30 ( .A1(m_rb_busy), .A2(m_rb_overflow), .A3(U_rbuf_n35), 
        .ZN(U_rbuf_n156) );
  OAI211_X1 U_rbuf_U29 ( .C1(U_rbuf_f_rbuf_state_1_), .C2(
        U_rbuf_f_rbuf_state_0_), .A(U_rbuf_n151), .B(U_rbuf_n150), .ZN(
        U_rbuf_n152) );
  INV_X4 U_rbuf_U28 ( .A(U_rbuf_n146), .ZN(U_rbuf_n6) );
  OAI21_X2 U_rbuf_U27 ( .B1(U_rbuf_n117), .B2(U_rbuf_n28), .A(U_rbuf_n137), 
        .ZN(hrdata[10]) );
  INV_X8 U_rbuf_U26 ( .A(U_rbuf_n119), .ZN(U_rbuf_n118) );
  AOI22_X1 U_rbuf_U25 ( .A1(miu_data[30]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_14_), .B2(U_rbuf_n177), .ZN(U_rbuf_n176) );
  AOI22_X1 U_rbuf_U24 ( .A1(miu_data[27]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_11_), .B2(U_rbuf_n177), .ZN(U_rbuf_n173) );
  AOI22_X1 U_rbuf_U23 ( .A1(miu_data[26]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_10_), .B2(U_rbuf_n177), .ZN(U_rbuf_n172) );
  AOI22_X1 U_rbuf_U22 ( .A1(miu_data[25]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_9_), .B2(U_rbuf_n177), .ZN(U_rbuf_n171) );
  AOI22_X1 U_rbuf_U21 ( .A1(miu_data[24]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_8_), .B2(U_rbuf_n177), .ZN(U_rbuf_n170) );
  AOI22_X1 U_rbuf_U20 ( .A1(miu_data[21]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_5_), .B2(U_rbuf_n177), .ZN(U_rbuf_n167) );
  AOI22_X1 U_rbuf_U19 ( .A1(miu_data[20]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_4_), .B2(U_rbuf_n177), .ZN(U_rbuf_n166) );
  AOI22_X1 U_rbuf_U18 ( .A1(miu_data[16]), .A2(U_rbuf_n178), .B1(
        U_rbuf_f_top_data_0_), .B2(U_rbuf_n177), .ZN(U_rbuf_n162) );
  OAI211_X1 U_rbuf_U17 ( .C1(U_rbuf_n3), .C2(U_rbuf_n17), .A(U_rbuf_n159), .B(
        U_rbuf_n4), .ZN(U_rbuf_n89) );
  NAND2_X1 U_rbuf_U16 ( .A1(U_rbuf_n3), .A2(U_rbuf_n17), .ZN(U_rbuf_n4) );
  NOR2_X1 U_rbuf_U15 ( .A1(miu_push_n), .A2(U_ctl_n96), .ZN(U_rbuf_n3) );
  OR2_X1 U_rbuf_U13 ( .A1(m_two_to_one), .A2(m_rb_sel_buf), .ZN(U_rbuf_n146)
         );
  OAI21_X2 U_rbuf_U12 ( .B1(U_rbuf_n160), .B2(U_ctl_n96), .A(n48), .ZN(
        U_rbuf_n145) );
  AOI21_X2 U_rbuf_U10 ( .B1(miu_data[13]), .B2(U_rbuf_n16), .A(n50), .ZN(
        U_rbuf_n38) );
  NAND2_X2 U_rbuf_U9 ( .A1(U_rbuf_n38), .A2(U_rbuf_n39), .ZN(hrdata[29]) );
  OAI21_X2 U_rbuf_U8 ( .B1(U_rbuf_n117), .B2(U_rbuf_n31), .A(U_rbuf_n140), 
        .ZN(hrdata[13]) );
  DFFR_X2 U_rbuf_f_top_data_reg_0_ ( .D(U_rbuf_n55), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_0_) );
  DFFR_X2 U_rbuf_f_top_data_reg_1_ ( .D(U_rbuf_n56), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_1_) );
  DFFR_X2 U_rbuf_f_top_data_reg_2_ ( .D(U_rbuf_n57), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_2_) );
  DFFR_X2 U_rbuf_f_top_data_reg_3_ ( .D(U_rbuf_n58), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_3_) );
  DFFR_X2 U_rbuf_f_top_data_reg_4_ ( .D(U_rbuf_n59), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_4_) );
  DFFR_X2 U_rbuf_f_top_data_reg_5_ ( .D(U_rbuf_n60), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_5_) );
  DFFR_X2 U_rbuf_f_top_data_reg_6_ ( .D(U_rbuf_n61), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_6_) );
  DFFR_X2 U_rbuf_f_top_data_reg_7_ ( .D(U_rbuf_n62), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_7_) );
  DFFR_X2 U_rbuf_f_top_data_reg_8_ ( .D(U_rbuf_n63), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_8_) );
  DFFR_X2 U_rbuf_f_top_data_reg_9_ ( .D(U_rbuf_n64), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_9_) );
  DFFR_X2 U_rbuf_f_top_data_reg_10_ ( .D(U_rbuf_n65), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_10_) );
  DFFR_X2 U_rbuf_f_top_data_reg_11_ ( .D(U_rbuf_n66), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_11_) );
  DFFR_X2 U_rbuf_f_top_data_reg_12_ ( .D(U_rbuf_n67), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_12_) );
  DFFR_X2 U_rbuf_f_top_data_reg_13_ ( .D(U_rbuf_n68), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_13_) );
  DFFR_X2 U_rbuf_f_top_data_reg_14_ ( .D(U_rbuf_n69), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_14_) );
  DFFR_X2 U_rbuf_f_top_data_reg_15_ ( .D(U_rbuf_n70), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_top_data_15_) );
  DFFR_X2 U_rbuf_f_btm_data_reg_0_ ( .D(U_rbuf_n71), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n18) );
  DFFR_X2 U_rbuf_f_btm_data_reg_1_ ( .D(U_rbuf_n72), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n19) );
  DFFR_X2 U_rbuf_f_btm_data_reg_2_ ( .D(U_rbuf_n73), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n20) );
  DFFR_X2 U_rbuf_f_btm_data_reg_3_ ( .D(U_rbuf_n74), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n21) );
  DFFR_X2 U_rbuf_f_btm_data_reg_4_ ( .D(U_rbuf_n75), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n22) );
  DFFR_X2 U_rbuf_f_btm_data_reg_5_ ( .D(U_rbuf_n76), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n23) );
  DFFR_X2 U_rbuf_f_btm_data_reg_6_ ( .D(U_rbuf_n77), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n24) );
  DFFR_X2 U_rbuf_f_btm_data_reg_7_ ( .D(U_rbuf_n78), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n25) );
  DFFR_X2 U_rbuf_f_btm_data_reg_8_ ( .D(U_rbuf_n79), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n26) );
  DFFR_X2 U_rbuf_f_btm_data_reg_9_ ( .D(U_rbuf_n80), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n27) );
  DFFR_X2 U_rbuf_f_btm_data_reg_10_ ( .D(U_rbuf_n81), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n28) );
  DFFR_X2 U_rbuf_f_btm_data_reg_11_ ( .D(U_rbuf_n82), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n29) );
  DFFR_X2 U_rbuf_f_btm_data_reg_12_ ( .D(U_rbuf_n83), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n30) );
  DFFR_X2 U_rbuf_f_btm_data_reg_13_ ( .D(U_rbuf_n84), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n31) );
  DFFR_X2 U_rbuf_f_btm_data_reg_14_ ( .D(U_rbuf_n85), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n33) );
  DFFR_X2 U_rbuf_f_btm_data_reg_15_ ( .D(U_rbuf_n86), .CK(hclk), .RN(hresetn), 
        .QN(U_rbuf_n32) );
  DFFR_X1 U_rbuf_f_rbuf_state_reg_1_ ( .D(U_rbuf_n87), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_rbuf_state_1_), .QN(U_rbuf_n35) );
  DFFR_X1 U_rbuf_f_rbuf_state_reg_0_ ( .D(U_rbuf_n88), .CK(hclk), .RN(hresetn), 
        .Q(U_rbuf_f_rbuf_state_0_) );
  DFFS_X2 U_rbuf_f_1st_half_reg ( .D(U_rbuf_n89), .CK(hclk), .SN(hresetn), .Q(
        U_rbuf_f_1st_half), .QN(U_rbuf_n17) );
  OAI21_X1 U_ctl_U457 ( .B1(U_rbuf_n120), .B2(U_ctl_n349), .A(m_two_to_one), 
        .ZN(U_ctl_n347) );
  NOR2_X1 U_ctl_U456 ( .A1(htrans[1]), .A2(U_ctl_n421), .ZN(U_ctl_N89) );
  INV_X4 U_ctl_U455 ( .A(U_ctl_n422), .ZN(U_ctl_n326) );
  NAND2_X2 U_ctl_U454 ( .A1(U_ctl_n249), .A2(U_ctl_n319), .ZN(m_af_data1_in_3_) );
  INV_X4 U_ctl_U453 ( .A(hburst[0]), .ZN(U_ctl_n278) );
  INV_X4 U_ctl_U452 ( .A(haddr[5]), .ZN(U_ctl_n276) );
  NAND2_X2 U_ctl_U451 ( .A1(U_ctl_fd_wr_width), .A2(big_endian), .ZN(
        U_ctl_n418) );
  INV_X1 U_ctl_U450 ( .A(hsel_reg), .ZN(U_ctl_n253) );
  AND3_X4 U_ctl_U448 ( .A1(U_ctl_n226), .A2(U_ctl_n229), .A3(haddr[5]), .ZN(
        U_ctl_n318) );
  MUX2_X2 U_ctl_U447 ( .A(hwdata[7]), .B(hwdata[23]), .S(U_ctl_n364), .Z(
        m_df_data_in[25]) );
  MUX2_X2 U_ctl_U446 ( .A(hwdata[0]), .B(hwdata[16]), .S(U_ctl_n364), .Z(
        m_df_data_in[18]) );
  AND4_X4 U_ctl_U445 ( .A1(U_ctl_n284), .A2(hburst[2]), .A3(U_ctl_n283), .A4(
        U_ctl_n282), .ZN(U_ctl_n286) );
  MUX2_X2 U_ctl_U444 ( .A(hwdata[15]), .B(hwdata[31]), .S(U_ctl_n364), .Z(
        m_df_data_in[33]) );
  MUX2_X2 U_ctl_U443 ( .A(hwdata[8]), .B(hwdata[24]), .S(U_ctl_n364), .Z(
        m_df_data_in[26]) );
  OR2_X4 U_ctl_U442 ( .A1(U_ctl_n398), .A2(U_ctl_n397), .ZN(U_ctl_n399) );
  NAND2_X2 U_ctl_U441 ( .A1(htrans[1]), .A2(htrans[0]), .ZN(U_ctl_n298) );
  NOR2_X2 U_ctl_U440 ( .A1(U_ctl_n63), .A2(U_ctl_n346), .ZN(U_ctl_n248) );
  OAI21_X2 U_ctl_U439 ( .B1(U_ctl_n166), .B2(U_ctl_fd_miu_col_width_2_), .A(
        U_ctl_n153), .ZN(U_ctl_n205) );
  NOR2_X2 U_ctl_U438 ( .A1(hburst[1]), .A2(hburst[2]), .ZN(U_ctl_n184) );
  NOR2_X2 U_ctl_U437 ( .A1(haddr[6]), .A2(haddr[7]), .ZN(U_ctl_n325) );
  NAND2_X2 U_ctl_U436 ( .A1(U_ctl_fd_miu_col_width_0_), .A2(
        U_ctl_fd_miu_col_width_2_), .ZN(U_ctl_n201) );
  NOR2_X2 U_ctl_U435 ( .A1(U_ctl_fd_miu_data_width_1_), .A2(
        U_ctl_fd_miu_data_width_0_), .ZN(U_ctl_n202) );
  NAND4_X2 U_ctl_U434 ( .A1(U_ctl_n205), .A2(U_ctl_n244), .A3(U_ctl_n325), 
        .A4(U_ctl_n204), .ZN(U_ctl_n206) );
  INV_X4 U_ctl_U433 ( .A(haddr[2]), .ZN(U_ctl_n288) );
  INV_X4 U_ctl_U432 ( .A(haddr[3]), .ZN(U_ctl_n289) );
  NAND2_X2 U_ctl_U431 ( .A1(U_ctl_n288), .A2(U_ctl_n289), .ZN(U_ctl_n269) );
  NAND2_X2 U_ctl_U430 ( .A1(U_ctl_n267), .A2(U_ctl_n276), .ZN(U_ctl_n329) );
  INV_X4 U_ctl_U429 ( .A(hsize[0]), .ZN(U_ctl_n227) );
  NAND2_X2 U_ctl_U428 ( .A1(U_ctl_n227), .A2(hsize[1]), .ZN(U_ctl_n199) );
  NAND2_X2 U_ctl_U427 ( .A1(U_ctl_n248), .A2(U_ctl_n207), .ZN(U_ctl_n208) );
  NOR2_X2 U_ctl_U426 ( .A1(haddr[7]), .A2(haddr[4]), .ZN(U_ctl_n193) );
  NAND3_X2 U_ctl_U425 ( .A1(U_ctl_n193), .A2(U_ctl_n288), .A3(U_ctl_n276), 
        .ZN(U_ctl_n198) );
  OAI211_X2 U_ctl_U424 ( .C1(U_ctl_fd_miu_col_width_1_), .C2(U_ctl_n154), .A(
        U_ctl_n202), .B(U_ctl_n194), .ZN(U_ctl_n195) );
  NOR2_X2 U_ctl_U423 ( .A1(haddr[3]), .A2(U_ctl_n195), .ZN(U_ctl_n196) );
  NAND2_X2 U_ctl_U422 ( .A1(U_ctl_n196), .A2(U_ctl_n235), .ZN(U_ctl_n197) );
  NOR2_X2 U_ctl_U421 ( .A1(U_ctl_n198), .A2(U_ctl_n197), .ZN(U_ctl_n200) );
  NAND2_X2 U_ctl_U420 ( .A1(U_ctl_n166), .A2(U_ctl_n201), .ZN(U_ctl_n167) );
  NOR2_X2 U_ctl_U419 ( .A1(U_ctl_n338), .A2(U_ctl_fd_hsel_mem), .ZN(U_ctl_n213) );
  NOR2_X2 U_ctl_U418 ( .A1(U_ctl_f_bh_state_1_), .A2(U_ctl_f_bh_state_2_), 
        .ZN(U_ctl_n305) );
  NAND2_X2 U_ctl_U417 ( .A1(U_ctl_n98), .A2(U_ctl_n158), .ZN(U_ctl_n221) );
  AOI21_X2 U_ctl_U416 ( .B1(miu_push_n), .B2(U_ctl_n209), .A(U_ctl_n221), .ZN(
        U_ctl_n211) );
  NOR3_X2 U_ctl_U415 ( .A1(U_ctl_fd_amba_bcnt_0_), .A2(U_ctl_fd_amba_bcnt_1_), 
        .A3(U_ctl_fd_amba_bcnt_2_), .ZN(U_ctl_n336) );
  NOR2_X2 U_ctl_U414 ( .A1(U_ctl_fd_amba_bcnt_3_), .A2(U_ctl_fd_incr), .ZN(
        U_ctl_n210) );
  NAND2_X2 U_ctl_U413 ( .A1(U_ctl_n336), .A2(U_ctl_n210), .ZN(U_ctl_n220) );
  NAND3_X2 U_ctl_U412 ( .A1(hready), .A2(U_ctl_n211), .A3(U_ctl_n220), .ZN(
        U_ctl_n212) );
  NAND2_X2 U_ctl_U411 ( .A1(hready), .A2(U_ctl_fd_rd_ready), .ZN(m_rb_pop_n)
         );
  NOR2_X2 U_ctl_U410 ( .A1(U_ctl_fr_prv_1wrap_tm), .A2(m_af_new_req), .ZN(
        U_ctl_n341) );
  NOR2_X2 U_ctl_U409 ( .A1(m_rb_overflow), .A2(U_ctl_n186), .ZN(U_ctl_n214) );
  NOR3_X2 U_ctl_U408 ( .A1(U_ctl_n339), .A2(U_ctl_fr_wr_bcnt_1_), .A3(
        U_ctl_fr_wr_bcnt_3_), .ZN(U_ctl_n308) );
  INV_X4 U_ctl_U407 ( .A(U_ctl_n304), .ZN(U_ctl_n292) );
  OAI211_X2 U_ctl_U406 ( .C1(U_ctl_n214), .C2(U_ctl_f_bh_state_0_), .A(
        U_ctl_n305), .B(U_ctl_n292), .ZN(U_ctl_n297) );
  AOI21_X2 U_ctl_U405 ( .B1(U_ctl_f_bh_state_1_), .B2(U_ctl_n95), .A(
        U_ctl_f_bh_state_2_), .ZN(U_ctl_n215) );
  AOI21_X2 U_ctl_U404 ( .B1(U_ctl_n297), .B2(U_ctl_n215), .A(m_df_wr_term), 
        .ZN(U_ctl_n218) );
  NAND2_X2 U_ctl_U403 ( .A1(U_ctl_n290), .A2(U_ctl_n216), .ZN(U_ctl_n217) );
  NAND2_X2 U_ctl_U402 ( .A1(U_ctl_n218), .A2(U_ctl_n217), .ZN(U_ctl_n219) );
  INV_X4 U_ctl_U401 ( .A(hwdata[14]), .ZN(U_ctl_n403) );
  INV_X4 U_ctl_U400 ( .A(hwdata[22]), .ZN(U_ctl_n402) );
  NOR2_X2 U_ctl_U399 ( .A1(U_ctl_n402), .A2(U_rbuf_n120), .ZN(U_ctl_n168) );
  NOR2_X2 U_ctl_U398 ( .A1(U_ctl_n169), .A2(U_ctl_n168), .ZN(U_ctl_n170) );
  NOR2_X2 U_ctl_U397 ( .A1(U_ctl_n170), .A2(U_ctl_n126), .ZN(U_ctl_n400) );
  NOR2_X2 U_ctl_U396 ( .A1(U_ctl_n126), .A2(big_endian), .ZN(U_ctl_n335) );
  INV_X4 U_ctl_U395 ( .A(U_ctl_n150), .ZN(U_ctl_n183) );
  NAND2_X2 U_ctl_U394 ( .A1(U_ctl_n253), .A2(U_ctl_n331), .ZN(U_ctl_n264) );
  INV_X4 U_ctl_U393 ( .A(U_ctl_n264), .ZN(U_ctl_n261) );
  AOI21_X2 U_ctl_U392 ( .B1(U_ctl_n276), .B2(U_ctl_f_offset_3_), .A(U_ctl_n159), .ZN(U_ctl_n254) );
  AOI21_X2 U_ctl_U391 ( .B1(U_ctl_n255), .B2(U_ctl_n254), .A(U_ctl_n298), .ZN(
        U_ctl_n258) );
  NAND2_X2 U_ctl_U389 ( .A1(U_ctl_n69), .A2(U_ctl_n258), .ZN(U_ctl_n262) );
  NOR2_X2 U_ctl_U388 ( .A1(U_ctl_n398), .A2(U_ctl_n346), .ZN(U_ctl_n251) );
  NAND2_X2 U_ctl_U387 ( .A1(U_ctl_n251), .A2(U_ctl_n250), .ZN(U_ctl_n252) );
  NAND2_X2 U_ctl_U386 ( .A1(U_ctl_n150), .A2(U_ctl_n252), .ZN(U_ctl_n180) );
  NAND3_X2 U_ctl_U385 ( .A1(U_ctl_n255), .A2(U_ctl_n254), .A3(U_ctl_n300), 
        .ZN(U_ctl_n223) );
  INV_X4 U_ctl_U384 ( .A(U_ctl_n189), .ZN(U_ctl_n249) );
  OAI21_X2 U_ctl_U383 ( .B1(U_ctl_n279), .B2(hburst[1]), .A(U_ctl_n243), .ZN(
        U_ctl_n246) );
  INV_X4 U_ctl_U382 ( .A(U_ctl_n329), .ZN(U_ctl_n245) );
  NOR4_X2 U_ctl_U381 ( .A1(U_ctl_n246), .A2(U_ctl_n245), .A3(U_ctl_n244), .A4(
        U_ctl_n250), .ZN(U_ctl_n247) );
  NAND2_X2 U_ctl_U380 ( .A1(U_ctl_n248), .A2(U_ctl_n247), .ZN(U_ctl_n319) );
  NAND3_X2 U_ctl_U378 ( .A1(U_ctl_n241), .A2(U_ctl_n278), .A3(hburst[1]), .ZN(
        U_ctl_n226) );
  NOR2_X2 U_ctl_U377 ( .A1(U_ctl_n89), .A2(U_ctl_n173), .ZN(m_af_data2_in[7])
         );
  NAND2_X2 U_ctl_U376 ( .A1(U_ctl_n251), .A2(hready), .ZN(U_ctl_n382) );
  INV_X4 U_ctl_U375 ( .A(U_ctl_n382), .ZN(U_ctl_n337) );
  OAI21_X2 U_ctl_U374 ( .B1(U_ctl_n336), .B2(U_ctl_n338), .A(U_ctl_n337), .ZN(
        U_ctl_n392) );
  AOI22_X2 U_ctl_U373 ( .A1(hburst[1]), .A2(U_ctl_n393), .B1(
        U_ctl_fd_amba_bcnt_3_), .B2(U_ctl_n392), .ZN(U_ctl_n394) );
  OAI21_X2 U_ctl_U372 ( .B1(U_ctl_fd_amba_bcnt_3_), .B2(U_ctl_n396), .A(
        U_ctl_n394), .ZN(U_ctl_n116) );
  NAND3_X2 U_ctl_U371 ( .A1(U_ctl_n98), .A2(big_endian), .A3(m_two_to_one), 
        .ZN(U_ctl_n364) );
  INV_X4 U_ctl_U370 ( .A(U_ctl_n262), .ZN(U_ctl_n263) );
  NOR2_X2 U_ctl_U369 ( .A1(U_ctl_n264), .A2(U_ctl_n263), .ZN(U_ctl_n284) );
  AOI21_X2 U_ctl_U368 ( .B1(U_ctl_n329), .B2(U_ctl_n278), .A(U_ctl_n275), .ZN(
        U_ctl_n283) );
  NAND2_X2 U_ctl_U367 ( .A1(U_ctl_n285), .A2(U_ctl_n180), .ZN(U_ctl_n179) );
  NAND3_X2 U_ctl_U366 ( .A1(U_ctl_n284), .A2(U_ctl_n282), .A3(U_ctl_n332), 
        .ZN(U_ctl_n273) );
  AOI211_X2 U_ctl_U365 ( .C1(U_ctl_n269), .C2(U_ctl_n268), .A(hburst[0]), .B(
        U_ctl_n267), .ZN(U_ctl_n271) );
  NOR2_X2 U_ctl_U364 ( .A1(U_ctl_n271), .A2(U_ctl_n270), .ZN(U_ctl_n272) );
  OAI22_X2 U_ctl_U363 ( .A1(U_ctl_n273), .A2(U_ctl_n272), .B1(U_ctl_n280), 
        .B2(U_ctl_n148), .ZN(U_ctl_n281) );
  NAND2_X2 U_ctl_U362 ( .A1(U_ctl_n281), .A2(U_ctl_n50), .ZN(U_ctl_n178) );
  NAND2_X2 U_ctl_U361 ( .A1(U_ctl_n179), .A2(U_ctl_n178), .ZN(m_af_data1_in_7_) );
  NAND2_X2 U_ctl_U360 ( .A1(U_ctl_n285), .A2(U_ctl_n50), .ZN(U_ctl_n182) );
  NAND2_X2 U_ctl_U359 ( .A1(U_ctl_n286), .A2(U_ctl_n180), .ZN(U_ctl_n181) );
  NAND2_X2 U_ctl_U358 ( .A1(U_ctl_n182), .A2(U_ctl_n181), .ZN(m_af_data1_in_8_) );
  NOR3_X2 U_ctl_U357 ( .A1(U_ctl_n382), .A2(htrans[0]), .A3(U_ctl_n332), .ZN(
        U_ctl_n323) );
  OAI21_X2 U_ctl_U355 ( .B1(U_ctl_n338), .B2(U_ctl_n143), .A(U_ctl_n337), .ZN(
        U_ctl_n395) );
  INV_X4 U_ctl_U353 ( .A(U_ctl_n233), .ZN(U_ctl_n228) );
  NOR4_X2 U_ctl_U352 ( .A1(U_ctl_n226), .A2(U_ctl_n228), .A3(hsize[0]), .A4(
        U_ctl_n288), .ZN(m_af_data2_in[12]) );
  INV_X4 U_ctl_U351 ( .A(U_ctl_n226), .ZN(U_ctl_n238) );
  AOI21_X2 U_ctl_U350 ( .B1(U_ctl_n237), .B2(U_ctl_n227), .A(U_ctl_n238), .ZN(
        U_ctl_n232) );
  NOR3_X2 U_ctl_U349 ( .A1(U_ctl_n232), .A2(U_ctl_n228), .A3(U_ctl_n289), .ZN(
        m_af_data2_in[13]) );
  NOR2_X2 U_ctl_U346 ( .A1(U_ctl_n163), .A2(U_ctl_n150), .ZN(m_af_data2_in[4])
         );
  AOI22_X2 U_ctl_U345 ( .A1(U_ctl_n230), .A2(U_ctl_n234), .B1(U_ctl_n238), 
        .B2(U_ctl_n380), .ZN(U_ctl_n231) );
  AOI211_X2 U_ctl_U344 ( .C1(U_ctl_n381), .C2(U_ctl_n234), .A(U_ctl_n233), .B(
        U_ctl_n238), .ZN(U_ctl_n236) );
  NOR2_X2 U_ctl_U343 ( .A1(U_ctl_n236), .A2(U_ctl_n235), .ZN(m_af_data2_in[16]) );
  NAND2_X2 U_ctl_U340 ( .A1(U_ctl_fd_narrow_trans), .A2(U_ctl_fd_haddr_1_), 
        .ZN(U_ctl_n349) );
  AOI21_X2 U_ctl_U339 ( .B1(U_rbuf_n120), .B2(U_ctl_n349), .A(U_ctl_n347), 
        .ZN(U_ctl_n375) );
  AOI21_X2 U_ctl_U338 ( .B1(U_rbuf_n120), .B2(U_ctl_n349), .A(U_ctl_n96), .ZN(
        U_ctl_n348) );
  OAI21_X2 U_ctl_U337 ( .B1(U_rbuf_n120), .B2(U_ctl_n349), .A(U_ctl_n348), 
        .ZN(U_ctl_n374) );
  AOI22_X2 U_ctl_U336 ( .A1(U_ctl_n375), .A2(hwdata[24]), .B1(U_ctl_n374), 
        .B2(hwdata[8]), .ZN(U_ctl_n350) );
  INV_X4 U_ctl_U335 ( .A(U_ctl_n350), .ZN(m_df_data_in[10]) );
  AOI22_X2 U_ctl_U334 ( .A1(U_ctl_n375), .A2(hwdata[31]), .B1(U_ctl_n374), 
        .B2(hwdata[15]), .ZN(U_ctl_n351) );
  INV_X4 U_ctl_U333 ( .A(U_ctl_n351), .ZN(m_df_data_in[17]) );
  NAND3_X2 U_ctl_U332 ( .A1(m_df_ready), .A2(m_af_ready), .A3(m_rb_ready), 
        .ZN(U_ctl_n294) );
  NAND2_X2 U_ctl_U331 ( .A1(U_ctl_n294), .A2(U_ctl_n151), .ZN(hready_resp) );
  AOI22_X2 U_ctl_U330 ( .A1(U_ctl_n375), .A2(hwdata[23]), .B1(U_ctl_n374), 
        .B2(hwdata[7]), .ZN(U_ctl_n376) );
  INV_X4 U_ctl_U329 ( .A(U_ctl_n376), .ZN(m_df_data_in[9]) );
  NAND4_X2 U_ctl_U328 ( .A1(U_ctl_n295), .A2(U_ctl_n297), .A3(U_ctl_n306), 
        .A4(U_ctl_n293), .ZN(hiu_terminate) );
  OAI22_X2 U_ctl_U327 ( .A1(U_ctl_n273), .A2(U_ctl_n266), .B1(U_ctl_n280), 
        .B2(U_ctl_n145), .ZN(U_ctl_n274) );
  NAND2_X2 U_ctl_U326 ( .A1(U_ctl_n274), .A2(U_ctl_n180), .ZN(U_ctl_n175) );
  NAND2_X2 U_ctl_U325 ( .A1(U_ctl_n175), .A2(U_ctl_n174), .ZN(m_af_data1_in_5_) );
  NAND2_X2 U_ctl_U324 ( .A1(U_ctl_n281), .A2(U_ctl_n180), .ZN(U_ctl_n177) );
  NAND2_X2 U_ctl_U323 ( .A1(U_ctl_n274), .A2(U_ctl_n50), .ZN(U_ctl_n176) );
  NAND2_X2 U_ctl_U322 ( .A1(U_ctl_n177), .A2(U_ctl_n176), .ZN(m_af_data1_in_6_) );
  AOI22_X2 U_ctl_U321 ( .A1(U_ctl_n375), .A2(hwdata[16]), .B1(U_ctl_n374), 
        .B2(hwdata[0]), .ZN(U_ctl_n358) );
  INV_X4 U_ctl_U320 ( .A(U_ctl_n358), .ZN(m_df_data_in[2]) );
  INV_X4 U_ctl_U319 ( .A(U_ctl_n364), .ZN(U_ctl_n363) );
  AOI22_X2 U_ctl_U318 ( .A1(U_ctl_n363), .A2(U_ctl_n371), .B1(U_ctl_n402), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[24]) );
  INV_X4 U_ctl_U317 ( .A(U_ctl_n375), .ZN(U_ctl_n373) );
  INV_X4 U_ctl_U316 ( .A(U_ctl_n374), .ZN(U_ctl_n372) );
  OAI22_X2 U_ctl_U315 ( .A1(U_ctl_n373), .A2(U_ctl_n359), .B1(U_ctl_n372), 
        .B2(U_ctl_n360), .ZN(m_df_data_in[14]) );
  OAI22_X2 U_ctl_U314 ( .A1(U_ctl_n373), .A2(U_ctl_n352), .B1(U_ctl_n372), 
        .B2(U_ctl_n353), .ZN(m_df_data_in[11]) );
  OAI22_X2 U_ctl_U313 ( .A1(U_ctl_n373), .A2(U_ctl_n356), .B1(U_ctl_n372), 
        .B2(U_ctl_n357), .ZN(m_df_data_in[13]) );
  OAI22_X2 U_ctl_U312 ( .A1(U_ctl_n373), .A2(U_ctl_n354), .B1(U_ctl_n372), 
        .B2(U_ctl_n355), .ZN(m_df_data_in[12]) );
  OAI22_X2 U_ctl_U311 ( .A1(U_ctl_n323), .A2(U_ctl_n395), .B1(U_ctl_n337), 
        .B2(U_ctl_n143), .ZN(U_ctl_n119) );
  AOI22_X2 U_ctl_U310 ( .A1(U_ctl_n363), .A2(U_ctl_n369), .B1(U_ctl_n370), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[23]) );
  OAI22_X2 U_ctl_U309 ( .A1(U_ctl_n403), .A2(U_ctl_n372), .B1(U_ctl_n373), 
        .B2(U_ctl_n362), .ZN(m_df_data_in[16]) );
  INV_X4 U_ctl_U308 ( .A(hwdata[29]), .ZN(U_ctl_n361) );
  OAI22_X2 U_ctl_U307 ( .A1(U_ctl_n361), .A2(U_ctl_n373), .B1(U_ctl_n222), 
        .B2(U_ctl_n372), .ZN(m_df_data_in[15]) );
  INV_X4 U_ctl_U306 ( .A(hwdata[18]), .ZN(U_ctl_n414) );
  AOI22_X2 U_ctl_U305 ( .A1(U_ctl_n363), .A2(U_ctl_n366), .B1(U_ctl_n414), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[20]) );
  INV_X4 U_ctl_U304 ( .A(hwdata[17]), .ZN(U_ctl_n417) );
  AOI22_X2 U_ctl_U303 ( .A1(U_ctl_n363), .A2(U_ctl_n365), .B1(U_ctl_n417), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[19]) );
  INV_X4 U_ctl_U302 ( .A(hwdata[20]), .ZN(U_ctl_n408) );
  AOI22_X2 U_ctl_U301 ( .A1(U_ctl_n363), .A2(U_ctl_n368), .B1(U_ctl_n408), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[22]) );
  INV_X4 U_ctl_U300 ( .A(hwdata[19]), .ZN(U_ctl_n411) );
  AOI22_X2 U_ctl_U299 ( .A1(U_ctl_n363), .A2(U_ctl_n367), .B1(U_ctl_n411), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[21]) );
  AOI22_X2 U_ctl_U298 ( .A1(m_af_data1_in_2_), .A2(U_ctl_n337), .B1(U_ctl_n421), .B2(U_ctl_fd_rd_ready), .ZN(U_ctl_n391) );
  INV_X4 U_ctl_U297 ( .A(U_ctl_n391), .ZN(U_ctl_n106) );
  OAI22_X2 U_ctl_U296 ( .A1(U_ctl_n402), .A2(U_ctl_n373), .B1(U_ctl_n372), 
        .B2(U_ctl_n371), .ZN(m_df_data_in[8]) );
  INV_X4 U_ctl_U295 ( .A(U_ctl_n286), .ZN(U_ctl_n287) );
  NOR2_X2 U_ctl_U294 ( .A1(U_ctl_n180), .A2(U_ctl_n287), .ZN(m_af_data1_in_9_)
         );
  OAI22_X2 U_ctl_U293 ( .A1(U_ctl_n373), .A2(U_ctl_n411), .B1(U_ctl_n372), 
        .B2(U_ctl_n367), .ZN(m_df_data_in[5]) );
  OAI22_X2 U_ctl_U292 ( .A1(U_ctl_n373), .A2(U_ctl_n414), .B1(U_ctl_n372), 
        .B2(U_ctl_n366), .ZN(m_df_data_in[4]) );
  OAI22_X2 U_ctl_U291 ( .A1(U_ctl_n370), .A2(U_ctl_n373), .B1(U_ctl_n372), 
        .B2(U_ctl_n369), .ZN(m_df_data_in[7]) );
  OAI22_X2 U_ctl_U290 ( .A1(U_ctl_n373), .A2(U_ctl_n408), .B1(U_ctl_n372), 
        .B2(U_ctl_n368), .ZN(m_df_data_in[6]) );
  OAI22_X2 U_ctl_U289 ( .A1(U_ctl_n373), .A2(U_ctl_n417), .B1(U_ctl_n372), 
        .B2(U_ctl_n365), .ZN(m_df_data_in[3]) );
  NAND2_X2 U_ctl_U288 ( .A1(U_ctl_n346), .A2(htrans[0]), .ZN(U_ctl_n397) );
  OAI22_X2 U_ctl_U287 ( .A1(U_ctl_n422), .A2(U_ctl_n400), .B1(
        U_ctl_fd_miu_data_width_1_), .B2(U_ctl_n326), .ZN(U_ctl_n401) );
  INV_X4 U_ctl_U286 ( .A(U_ctl_n401), .ZN(U_ctl_n125) );
  NOR3_X2 U_ctl_U285 ( .A1(U_ctl_n400), .A2(U_ctl_n183), .A3(U_ctl_n378), .ZN(
        m_af_data1_in_11_) );
  AOI22_X2 U_ctl_U284 ( .A1(U_ctl_n180), .A2(U_ctl_n326), .B1(U_ctl_n422), 
        .B2(U_ctl_n324), .ZN(U_ctl_n124) );
  AOI22_X2 U_ctl_U283 ( .A1(U_ctl_n361), .A2(U_ctl_n364), .B1(U_ctl_n222), 
        .B2(U_ctl_n363), .ZN(m_df_data_in[31]) );
  AOI22_X2 U_ctl_U282 ( .A1(hwdata[11]), .A2(U_ctl_n335), .B1(
        U_ctl_f_col_width[2]), .B2(U_ctl_n126), .ZN(U_ctl_n410) );
  OAI21_X2 U_ctl_U281 ( .B1(U_ctl_n418), .B2(U_ctl_n411), .A(U_ctl_n410), .ZN(
        U_ctl_n133) );
  OAI22_X2 U_ctl_U280 ( .A1(U_ctl_n422), .A2(U_ctl_n133), .B1(
        U_ctl_fd_miu_col_width_2_), .B2(U_ctl_n326), .ZN(U_ctl_n412) );
  INV_X4 U_ctl_U279 ( .A(U_ctl_n412), .ZN(U_ctl_n129) );
  AOI22_X2 U_ctl_U278 ( .A1(U_ctl_n363), .A2(U_ctl_n403), .B1(U_ctl_n362), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[32]) );
  AOI22_X2 U_ctl_U277 ( .A1(hwdata[10]), .A2(U_ctl_n335), .B1(
        U_ctl_f_col_width[1]), .B2(U_ctl_n126), .ZN(U_ctl_n413) );
  OAI21_X2 U_ctl_U276 ( .B1(U_ctl_n418), .B2(U_ctl_n414), .A(U_ctl_n413), .ZN(
        U_ctl_n134) );
  OAI22_X2 U_ctl_U275 ( .A1(U_ctl_n422), .A2(U_ctl_n134), .B1(
        U_ctl_fd_miu_col_width_1_), .B2(U_ctl_n326), .ZN(U_ctl_n415) );
  INV_X4 U_ctl_U274 ( .A(U_ctl_n415), .ZN(U_ctl_n130) );
  AOI22_X2 U_ctl_U273 ( .A1(hwdata[12]), .A2(U_ctl_n335), .B1(
        U_ctl_f_col_width[3]), .B2(U_ctl_n126), .ZN(U_ctl_n407) );
  OAI21_X2 U_ctl_U272 ( .B1(U_ctl_n418), .B2(U_ctl_n408), .A(U_ctl_n407), .ZN(
        U_ctl_n132) );
  OAI22_X2 U_ctl_U271 ( .A1(U_ctl_n422), .A2(U_ctl_n132), .B1(
        U_ctl_fd_miu_col_width_3_), .B2(U_ctl_n326), .ZN(U_ctl_n409) );
  INV_X4 U_ctl_U270 ( .A(U_ctl_n409), .ZN(U_ctl_n128) );
  AOI22_X2 U_ctl_U269 ( .A1(hwdata[9]), .A2(U_ctl_n335), .B1(
        U_ctl_f_col_width[0]), .B2(U_ctl_n126), .ZN(U_ctl_n416) );
  OAI21_X2 U_ctl_U268 ( .B1(U_ctl_n418), .B2(U_ctl_n417), .A(U_ctl_n416), .ZN(
        U_ctl_n135) );
  OAI22_X2 U_ctl_U267 ( .A1(U_ctl_n422), .A2(U_ctl_n135), .B1(
        U_ctl_fd_miu_col_width_0_), .B2(U_ctl_n326), .ZN(U_ctl_n419) );
  INV_X4 U_ctl_U266 ( .A(U_ctl_n419), .ZN(U_ctl_n131) );
  OAI22_X2 U_ctl_U265 ( .A1(U_ctl_n326), .A2(U_ctl_n62), .B1(m_af_data1_in_2_), 
        .B2(U_ctl_n399), .ZN(U_ctl_n121) );
  NAND4_X2 U_ctl_U264 ( .A1(hwrite), .A2(U_ctl_n380), .A3(U_ctl_n381), .A4(
        U_ctl_n326), .ZN(U_ctl_n327) );
  NAND2_X2 U_ctl_U263 ( .A1(U_ctl_n171), .A2(U_ctl_f_data_width_0_), .ZN(
        U_ctl_n405) );
  OAI211_X2 U_ctl_U262 ( .C1(U_ctl_n418), .C2(U_ctl_n406), .A(U_ctl_n405), .B(
        U_ctl_n404), .ZN(U_ctl_n127) );
  AOI22_X2 U_ctl_U261 ( .A1(U_ctl_n363), .A2(U_ctl_n355), .B1(U_ctl_n354), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[28]) );
  AOI22_X2 U_ctl_U260 ( .A1(U_ctl_n363), .A2(U_ctl_n353), .B1(U_ctl_n352), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[27]) );
  AOI22_X2 U_ctl_U259 ( .A1(U_ctl_n363), .A2(U_ctl_n357), .B1(U_ctl_n356), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[29]) );
  AOI22_X2 U_ctl_U258 ( .A1(U_ctl_n363), .A2(U_ctl_n360), .B1(U_ctl_n359), 
        .B2(U_ctl_n364), .ZN(m_df_data_in[30]) );
  NOR2_X2 U_ctl_U257 ( .A1(m_af_dummy_req), .A2(U_ctl_n342), .ZN(U_ctl_N236)
         );
  AOI22_X2 U_ctl_U256 ( .A1(U_ctl_n183), .A2(U_ctl_n326), .B1(U_ctl_n422), 
        .B2(U_ctl_n96), .ZN(U_ctl_n122) );
  AOI22_X2 U_ctl_U255 ( .A1(U_ctl_n150), .A2(U_ctl_n326), .B1(U_ctl_n147), 
        .B2(U_ctl_n422), .ZN(U_ctl_n123) );
  OAI22_X2 U_ctl_U254 ( .A1(hwrite), .A2(U_ctl_n399), .B1(U_ctl_n326), .B2(
        U_ctl_n146), .ZN(U_ctl_n120) );
  NOR4_X2 U_ctl_U253 ( .A1(U_ctl_n340), .A2(hiu_burst_size[5]), .A3(
        hiu_burst_size[1]), .A4(U_ctl_n310), .ZN(U_ctl_n309) );
  AOI211_X2 U_ctl_U252 ( .C1(U_ctl_n309), .C2(U_ctl_n384), .A(
        U_ctl_f_hiu_terminate), .B(U_ctl_n386), .ZN(U_ctl_n313) );
  NAND2_X2 U_ctl_U251 ( .A1(U_ctl_C64_DATA2_5), .A2(U_ctl_n313), .ZN(
        U_ctl_n312) );
  NOR3_X2 U_ctl_U250 ( .A1(U_ctl_f_hiu_terminate), .A2(U_ctl_n385), .A3(
        U_ctl_n384), .ZN(U_ctl_n389) );
  NOR3_X2 U_ctl_U249 ( .A1(U_ctl_fr_prv_1wrap), .A2(U_ctl_n144), .A3(
        U_ctl_n386), .ZN(U_ctl_n388) );
  AOI22_X2 U_ctl_U248 ( .A1(U_ctl_fr_wr_bcnt_5_), .A2(U_ctl_n389), .B1(
        U_ctl_n388), .B2(hiu_burst_size[5]), .ZN(U_ctl_n387) );
  NAND3_X2 U_ctl_U247 ( .A1(U_ctl_n312), .A2(U_ctl_n387), .A3(U_ctl_n311), 
        .ZN(U_ctl_n100) );
  OAI22_X2 U_ctl_U246 ( .A1(U_ctl_n422), .A2(haddr[1]), .B1(U_ctl_fd_haddr_1_), 
        .B2(U_ctl_n326), .ZN(U_ctl_n420) );
  INV_X4 U_ctl_U245 ( .A(U_ctl_n420), .ZN(U_ctl_n137) );
  AOI21_X2 U_ctl_U244 ( .B1(U_ctl_n303), .B2(U_ctl_n302), .A(U_ctl_n307), .ZN(
        U_ctl_n_bh_state[2]) );
  AOI21_X2 U_ctl_U243 ( .B1(U_ctl_n142), .B2(U_ctl_n343), .A(U_ctl_n397), .ZN(
        U_ctl_n344) );
  AOI211_X2 U_ctl_U242 ( .C1(U_ctl_n300), .C2(U_ctl_n345), .A(U_ctl_n301), .B(
        U_ctl_n344), .ZN(U_ctl_n296) );
  NOR2_X2 U_ctl_U241 ( .A1(U_ctl_n307), .A2(U_ctl_n296), .ZN(U_ctl_n_sel_buf)
         );
  AOI22_X2 U_ctl_U240 ( .A1(n51), .A2(U_ctl_n326), .B1(U_ctl_n156), .B2(
        U_ctl_n422), .ZN(U_ctl_n141) );
  AOI22_X2 U_ctl_U239 ( .A1(U_ctl_fr_wr_bcnt_0_), .A2(U_ctl_n389), .B1(
        U_ctl_n388), .B2(hiu_burst_size[0]), .ZN(U_ctl_n390) );
  NAND3_X2 U_ctl_U238 ( .A1(U_ctl_n316), .A2(U_ctl_n390), .A3(U_ctl_n315), 
        .ZN(U_ctl_n105) );
  OAI211_X2 U_ctl_U237 ( .C1(U_ctl_n206), .C2(U_ctl_n329), .A(htrans[0]), .B(
        U_ctl_n331), .ZN(U_ctl_n207) );
  NAND2_X2 U_ctl_U236 ( .A1(U_ctl_n165), .A2(htrans[0]), .ZN(U_ctl_n216) );
  INV_X1 U_ctl_U235 ( .A(miu_pop_n), .ZN(U_ctl_n384) );
  NOR2_X1 U_ctl_U234 ( .A1(hiu_rw), .A2(m_af_new_req), .ZN(U_ctl_n385) );
  NAND2_X2 U_ctl_U233 ( .A1(U_ctl_n397), .A2(hready), .ZN(U_ctl_n422) );
  NOR2_X2 U_ctl_U232 ( .A1(U_ctl_n309), .A2(miu_pop_n), .ZN(
        U_ctl_DP_OP_140_125_8947_I2) );
  NAND3_X1 U_ctl_U231 ( .A1(htrans[0]), .A2(U_ctl_n336), .A3(U_ctl_n337), .ZN(
        U_ctl_n396) );
  OAI22_X2 U_ctl_U230 ( .A1(U_ctl_n382), .A2(U_ctl_n331), .B1(U_ctl_n326), 
        .B2(U_ctl_n98), .ZN(U_ctl_n139) );
  NOR2_X1 U_ctl_U229 ( .A1(U_ctl_n187), .A2(U_ctl_n298), .ZN(U_ctl_n257) );
  NAND2_X1 U_ctl_U228 ( .A1(hsize[1]), .A2(hsize[0]), .ZN(U_ctl_n380) );
  AOI221_X1 U_ctl_U227 ( .B1(hsize[0]), .B2(U_ctl_n378), .C1(haddr[0]), .C2(
        U_ctl_n378), .A(hsize[1]), .ZN(U_ctl_n379) );
  INV_X1 U_ctl_U226 ( .A(hsize[1]), .ZN(U_ctl_n230) );
  AOI211_X1 U_ctl_U225 ( .C1(U_ctl_n232), .C2(hsize[1]), .A(hsize[2]), .B(
        U_ctl_n276), .ZN(m_af_data2_in[15]) );
  NAND3_X2 U_ctl_U224 ( .A1(U_ctl_n47), .A2(U_ctl_n244), .A3(U_ctl_n331), .ZN(
        U_ctl_n187) );
  AOI22_X1 U_ctl_U223 ( .A1(U_ctl_n184), .A2(U_ctl_n383), .B1(U_ctl_n422), 
        .B2(U_ctl_n160), .ZN(U_ctl_n140) );
  AOI21_X2 U_ctl_U222 ( .B1(U_ctl_n187), .B2(U_ctl_n213), .A(U_ctl_n212), .ZN(
        U_ctl_n290) );
  INV_X1 U_ctl_U221 ( .A(hburst[2]), .ZN(U_ctl_n241) );
  NAND3_X1 U_ctl_U220 ( .A1(U_ctl_n275), .A2(U_ctl_n278), .A3(hburst[2]), .ZN(
        U_ctl_n229) );
  NAND2_X1 U_ctl_U219 ( .A1(U_ctl_n320), .A2(hburst[2]), .ZN(U_ctl_n268) );
  AOI21_X1 U_ctl_U218 ( .B1(U_ctl_n269), .B2(U_ctl_n278), .A(hburst[2]), .ZN(
        U_ctl_n270) );
  NOR2_X1 U_ctl_U217 ( .A1(hsel_reg), .A2(n8), .ZN(U_ctl_n398) );
  NAND2_X1 U_ctl_U216 ( .A1(haddr[3]), .A2(haddr[2]), .ZN(U_ctl_n265) );
  NAND2_X1 U_ctl_U215 ( .A1(U_ctl_n226), .A2(haddr[4]), .ZN(U_ctl_n317) );
  AOI21_X1 U_ctl_U214 ( .B1(U_ctl_n65), .B2(U_ctl_n258), .A(U_ctl_n257), .ZN(
        U_ctl_n282) );
  INV_X1 U_ctl_U213 ( .A(hsize[2]), .ZN(U_ctl_n381) );
  NOR3_X1 U_ctl_U212 ( .A1(U_ctl_n231), .A2(hsize[2]), .A3(U_ctl_n320), .ZN(
        m_af_data2_in[14]) );
  NAND2_X1 U_ctl_U211 ( .A1(U_ctl_n84), .A2(haddr[3]), .ZN(U_ctl_n75) );
  INV_X4 U_ctl_U209 ( .A(U_ctl_n185), .ZN(U_ctl_n69) );
  NAND2_X2 U_ctl_U208 ( .A1(U_ctl_n67), .A2(U_ctl_n66), .ZN(U_ctl_n185) );
  INV_X4 U_ctl_U207 ( .A(n8), .ZN(U_ctl_n63) );
  NAND2_X2 U_ctl_U206 ( .A1(U_ctl_n61), .A2(U_ctl_f_amba_bsz2[3]), .ZN(
        U_ctl_n60) );
  NOR2_X1 U_ctl_U205 ( .A1(U_ctl_n90), .A2(U_ctl_n223), .ZN(U_ctl_n61) );
  NAND2_X2 U_ctl_U204 ( .A1(U_ctl_n23), .A2(U_ctl_n50), .ZN(U_ctl_n174) );
  OAI22_X2 U_ctl_U203 ( .A1(U_ctl_n330), .A2(m_af_data1_in_0_), .B1(U_ctl_n326), .B2(U_ctl_n126), .ZN(U_ctl_n136) );
  OAI22_X2 U_ctl_U202 ( .A1(m_af_data1_in_0_), .A2(U_ctl_n421), .B1(U_ctl_n326), .B2(U_ctl_n158), .ZN(U_ctl_n138) );
  NAND2_X2 U_ctl_U201 ( .A1(m_af_data1_in_0_), .A2(U_ctl_n208), .ZN(U_ctl_n84)
         );
  NAND3_X2 U_ctl_U200 ( .A1(m_af_data1_in_0_), .A2(n49), .A3(U_ctl_n208), .ZN(
        U_ctl_n85) );
  INV_X1 U_ctl_U199 ( .A(hburst[1]), .ZN(U_ctl_n275) );
  INV_X2 U_ctl_U197 ( .A(haddr[6]), .ZN(U_ctl_n235) );
  INV_X2 U_ctl_U196 ( .A(htrans[1]), .ZN(U_ctl_n346) );
  INV_X2 U_ctl_U195 ( .A(haddr[1]), .ZN(U_ctl_n378) );
  INV_X2 U_ctl_U194 ( .A(hwdata[2]), .ZN(U_ctl_n366) );
  INV_X2 U_ctl_U193 ( .A(hwrite), .ZN(m_af_data1_in_2_) );
  INV_X2 U_ctl_U192 ( .A(hwdata[1]), .ZN(U_ctl_n365) );
  INV_X2 U_ctl_U191 ( .A(hwdata[6]), .ZN(U_ctl_n371) );
  INV_X2 U_ctl_U190 ( .A(hwdata[10]), .ZN(U_ctl_n355) );
  INV_X2 U_ctl_U189 ( .A(hwdata[28]), .ZN(U_ctl_n359) );
  INV_X2 U_ctl_U188 ( .A(hwdata[4]), .ZN(U_ctl_n368) );
  INV_X2 U_ctl_U187 ( .A(hwdata[12]), .ZN(U_ctl_n360) );
  NAND2_X2 U_ctl_U186 ( .A1(hsel_reg), .A2(htrans[1]), .ZN(m_af_data1_in_0_)
         );
  INV_X2 U_ctl_U185 ( .A(hwdata[26]), .ZN(U_ctl_n354) );
  INV_X2 U_ctl_U184 ( .A(hwdata[3]), .ZN(U_ctl_n367) );
  INV_X2 U_ctl_U183 ( .A(hwdata[11]), .ZN(U_ctl_n357) );
  INV_X2 U_ctl_U182 ( .A(hwdata[27]), .ZN(U_ctl_n356) );
  INV_X2 U_ctl_U181 ( .A(hwdata[25]), .ZN(U_ctl_n352) );
  INV_X2 U_ctl_U180 ( .A(hwdata[9]), .ZN(U_ctl_n353) );
  INV_X2 U_ctl_U179 ( .A(hwdata[30]), .ZN(U_ctl_n362) );
  INV_X2 U_ctl_U178 ( .A(hwdata[5]), .ZN(U_ctl_n369) );
  INV_X2 U_ctl_U177 ( .A(hwdata[21]), .ZN(U_ctl_n370) );
  INV_X2 U_ctl_U176 ( .A(hwdata[13]), .ZN(U_ctl_n222) );
  NAND2_X1 U_ctl_U175 ( .A1(hwdata[21]), .A2(U_ctl_n402), .ZN(U_ctl_n406) );
  INV_X4 U_ctl_U174 ( .A(U_ctl_n184), .ZN(U_ctl_n332) );
  INV_X1 U_ctl_U173 ( .A(U_ctl_n325), .ZN(U_ctl_n328) );
  OR3_X2 U_ctl_U172 ( .A1(U_ctl_fr_wr_bcnt_2_), .A2(U_ctl_fr_wr_bcnt_4_), .A3(
        U_ctl_fr_wr_bcnt_5_), .ZN(U_ctl_n339) );
  NAND3_X1 U_ctl_U171 ( .A1(U_ctl_f_bh_state_0_), .A2(U_ctl_f_bh_state_1_), 
        .A3(U_ctl_n142), .ZN(U_ctl_n343) );
  NOR2_X2 U_ctl_U170 ( .A1(U_ctl_fd_wr_width), .A2(U_ctl_f_data_width_0_), 
        .ZN(U_ctl_n55) );
  OR3_X2 U_ctl_U169 ( .A1(U_ctl_n144), .A2(U_ctl_f_burst_done), .A3(
        U_ctl_f_burst_done2), .ZN(U_ctl_n293) );
  NOR2_X2 U_ctl_U168 ( .A1(hsize[1]), .A2(hsize[2]), .ZN(U_ctl_n233) );
  NAND2_X1 U_ctl_U167 ( .A1(U_ctl_n229), .A2(hsize[0]), .ZN(U_ctl_n234) );
  INV_X2 U_ctl_U166 ( .A(U_ctl_n397), .ZN(m_rb_busy) );
  INV_X2 U_ctl_U165 ( .A(U_ctl_n229), .ZN(U_ctl_n237) );
  INV_X1 U_ctl_U164 ( .A(hready), .ZN(U_ctl_n421) );
  INV_X1 U_ctl_U163 ( .A(U_ctl_n269), .ZN(U_ctl_n242) );
  AOI21_X1 U_ctl_U162 ( .B1(U_ctl_n332), .B2(U_ctl_n288), .A(hburst[0]), .ZN(
        U_ctl_n260) );
  NOR2_X1 U_ctl_U161 ( .A1(U_ctl_n403), .A2(big_endian), .ZN(U_ctl_n169) );
  NAND3_X1 U_ctl_U160 ( .A1(U_ctl_n269), .A2(U_ctl_n278), .A3(U_ctl_n265), 
        .ZN(U_ctl_n266) );
  NAND2_X2 U_ctl_U159 ( .A1(U_ctl_n332), .A2(U_ctl_n278), .ZN(U_ctl_n244) );
  NOR2_X2 U_ctl_U158 ( .A1(U_ctl_n269), .A2(haddr[4]), .ZN(U_ctl_n267) );
  OAI21_X1 U_ctl_U157 ( .B1(U_ctl_n201), .B2(U_ctl_fd_miu_col_width_3_), .A(
        U_ctl_fd_miu_col_width_1_), .ZN(U_ctl_n203) );
  INV_X2 U_ctl_U156 ( .A(U_ctl_n343), .ZN(U_ctl_n345) );
  NAND2_X1 U_ctl_U155 ( .A1(U_ctl_f_bh_state_2_), .A2(m_rb_busy), .ZN(
        U_ctl_n302) );
  INV_X2 U_ctl_U154 ( .A(U_ctl_n267), .ZN(U_ctl_n279) );
  AOI21_X1 U_ctl_U153 ( .B1(U_ctl_n242), .B2(U_ctl_n241), .A(htrans[0]), .ZN(
        U_ctl_n243) );
  NOR2_X1 U_ctl_U151 ( .A1(hburst[0]), .A2(U_ctl_n422), .ZN(U_ctl_n383) );
  NAND3_X1 U_ctl_U150 ( .A1(hwdata[13]), .A2(U_ctl_n335), .A3(U_ctl_n403), 
        .ZN(U_ctl_n404) );
  INV_X2 U_ctl_U149 ( .A(U_ctl_n335), .ZN(U_ctl_n54) );
  INV_X1 U_ctl_U148 ( .A(U_ctl_n317), .ZN(U_ctl_n87) );
  AND2_X2 U_ctl_U147 ( .A1(U_ctl_n203), .A2(U_ctl_n202), .ZN(U_ctl_n204) );
  NOR2_X2 U_ctl_U146 ( .A1(U_ctl_n199), .A2(hsize[2]), .ZN(U_ctl_n331) );
  NOR2_X2 U_ctl_U145 ( .A1(hwdata[13]), .A2(U_ctl_n54), .ZN(U_ctl_n56) );
  NAND3_X1 U_ctl_U144 ( .A1(U_ctl_n329), .A2(U_ctl_n278), .A3(U_ctl_n276), 
        .ZN(U_ctl_n277) );
  OR4_X2 U_ctl_U143 ( .A1(U_ctl_n379), .A2(U_ctl_n329), .A3(U_ctl_n328), .A4(
        U_ctl_n327), .ZN(U_ctl_n330) );
  INV_X2 U_ctl_U142 ( .A(U_ctl_n331), .ZN(U_ctl_n250) );
  NAND2_X1 U_ctl_U141 ( .A1(U_ctl_n170), .A2(U_ctl_fd_wr_width), .ZN(
        U_ctl_n171) );
  NOR2_X2 U_ctl_U140 ( .A1(U_ctl_n56), .A2(U_ctl_n55), .ZN(U_ctl_n58) );
  OR4_X2 U_ctl_U139 ( .A1(hiu_burst_size[0]), .A2(hiu_burst_size[4]), .A3(
        hiu_burst_size[2]), .A4(hiu_burst_size[3]), .ZN(U_ctl_n340) );
  INV_X2 U_ctl_U138 ( .A(U_ctl_n385), .ZN(U_ctl_n386) );
  NAND2_X2 U_ctl_U137 ( .A1(U_ctl_n58), .A2(U_ctl_n57), .ZN(U_ctl_n150) );
  INV_X4 U_ctl_U136 ( .A(U_ctl_n180), .ZN(U_ctl_n50) );
  NAND2_X1 U_ctl_U135 ( .A1(hwrite), .A2(U_ctl_n337), .ZN(U_ctl_n299) );
  INV_X2 U_ctl_U133 ( .A(hiu_wrap_burst), .ZN(U_ctl_n342) );
  AND2_X2 U_ctl_U132 ( .A1(U_ctl_n165), .A2(htrans[0]), .ZN(U_ctl_n94) );
  INV_X2 U_ctl_U131 ( .A(U_ctl_n70), .ZN(U_ctl_n393) );
  NAND2_X1 U_ctl_U130 ( .A1(U_ctl_n314), .A2(U_ctl_N288), .ZN(U_ctl_n311) );
  OAI21_X1 U_ctl_U129 ( .B1(U_ctl_n84), .B2(U_ctl_n159), .A(U_ctl_n319), .ZN(
        U_ctl_n111) );
  NAND2_X1 U_ctl_U128 ( .A1(U_ctl_n314), .A2(U_ctl_n97), .ZN(U_ctl_n315) );
  OAI21_X2 U_ctl_U126 ( .B1(n8), .B2(U_ctl_n155), .A(U_ctl_n94), .ZN(m_rb_done) );
  OAI21_X1 U_ctl_U125 ( .B1(U_ctl_n84), .B2(U_ctl_n83), .A(U_ctl_n82), .ZN(
        U_ctl_n107) );
  OAI21_X1 U_ctl_U124 ( .B1(U_ctl_n84), .B2(U_ctl_n74), .A(U_ctl_n73), .ZN(
        U_ctl_n115) );
  OAI21_X1 U_ctl_U123 ( .B1(U_ctl_n84), .B2(U_ctl_n77), .A(U_ctl_n82), .ZN(
        U_ctl_n112) );
  OAI21_X1 U_ctl_U122 ( .B1(U_ctl_n84), .B2(U_ctl_n81), .A(U_ctl_n75), .ZN(
        U_ctl_n108) );
  OAI21_X1 U_ctl_U121 ( .B1(U_ctl_n84), .B2(U_ctl_n76), .A(U_ctl_n75), .ZN(
        U_ctl_n113) );
  OAI21_X1 U_ctl_U120 ( .B1(U_ctl_n84), .B2(U_ctl_n79), .A(U_ctl_n78), .ZN(
        U_ctl_n110) );
  AOI21_X2 U_ctl_U119 ( .B1(U_ctl_n291), .B2(U_ctl_n290), .A(m_df_wr_term), 
        .ZN(U_ctl_n295) );
  INV_X1 U_ctl_U118 ( .A(U_ctl_n257), .ZN(U_ctl_n256) );
  NAND2_X1 U_ctl_U116 ( .A1(U_ctl_C64_DATA2_0), .A2(U_ctl_n313), .ZN(
        U_ctl_n316) );
  INV_X2 U_ctl_U115 ( .A(U_ctl_n295), .ZN(U_ctl_n307) );
  INV_X2 U_ctl_U114 ( .A(U_ctl_n219), .ZN(U_ctl_n66) );
  AND2_X2 U_ctl_U113 ( .A1(hiu_terminate), .A2(U_ctl_N236), .ZN(U_ctl_N237) );
  OAI21_X1 U_ctl_U112 ( .B1(U_ctl_n301), .B2(U_ctl_n345), .A(U_ctl_n300), .ZN(
        U_ctl_n303) );
  NOR2_X2 U_ctl_U111 ( .A1(U_ctl_n164), .A2(U_ctl_n259), .ZN(U_ctl_n90) );
  NOR2_X2 U_ctl_U110 ( .A1(U_ctl_n69), .A2(U_ctl_n65), .ZN(U_ctl_n172) );
  OAI21_X2 U_ctl_U108 ( .B1(U_ctl_n61), .B2(U_ctl_n91), .A(U_ctl_n60), .ZN(
        U_ctl_n92) );
  NOR2_X2 U_ctl_U107 ( .A1(U_ctl_n172), .A2(U_ctl_n223), .ZN(U_ctl_n189) );
  NOR2_X2 U_ctl_U105 ( .A1(U_ctl_n150), .A2(U_ctl_n92), .ZN(U_ctl_n173) );
  NOR2_X2 U_ctl_U104 ( .A1(U_ctl_n189), .A2(U_ctl_n87), .ZN(U_ctl_n88) );
  NAND2_X2 U_ctl_U103 ( .A1(U_ctl_n85), .A2(hready), .ZN(m_af_push1_n) );
  NOR2_X2 U_ctl_U101 ( .A1(m_af_push1_n), .A2(hwrite), .ZN(m_rb_start) );
  NOR2_X2 U_ctl_U100 ( .A1(U_ctl_n86), .A2(U_ctl_n88), .ZN(U_ctl_n225) );
  INV_X2 U_ctl_U99 ( .A(haddr[4]), .ZN(U_ctl_n320) );
  INV_X2 U_ctl_U98 ( .A(htrans[0]), .ZN(U_ctl_n338) );
  INV_X2 U_ctl_U97 ( .A(U_ctl_n298), .ZN(U_ctl_n300) );
  NAND2_X2 U_ctl_U96 ( .A1(U_ctl_fd_miu_col_width_3_), .A2(
        U_ctl_fd_miu_col_width_1_), .ZN(U_ctl_n194) );
  NAND2_X2 U_ctl_U94 ( .A1(n8), .A2(U_ctl_fd_wr_bz), .ZN(U_ctl_n64) );
  NAND3_X1 U_ctl_U93 ( .A1(U_ctl_n305), .A2(U_ctl_fd_rd_bz), .A3(
        U_ctl_f_bh_state_0_), .ZN(U_ctl_n209) );
  INV_X4 U_ctl_U92 ( .A(U_ctl_n64), .ZN(U_ctl_n65) );
  INV_X1 U_ctl_U91 ( .A(U_ctl_n318), .ZN(U_ctl_n91) );
  NOR2_X2 U_ctl_U90 ( .A1(U_ctl_n63), .A2(U_ctl_n62), .ZN(U_ctl_n259) );
  OR2_X2 U_ctl_U89 ( .A1(hwdata[21]), .A2(U_ctl_n418), .ZN(U_ctl_n57) );
  INV_X4 U_ctl_U88 ( .A(U_ctl_n341), .ZN(U_ctl_n186) );
  NAND2_X1 U_ctl_U87 ( .A1(U_ctl_n308), .A2(U_ctl_n97), .ZN(U_ctl_n310) );
  NAND2_X2 U_ctl_U85 ( .A1(U_ctl_n94), .A2(n8), .ZN(U_ctl_n291) );
  NAND2_X1 U_ctl_U84 ( .A1(U_ctl_n84), .A2(haddr[5]), .ZN(U_ctl_n73) );
  NAND2_X1 U_ctl_U83 ( .A1(U_ctl_n84), .A2(haddr[2]), .ZN(U_ctl_n82) );
  NAND2_X1 U_ctl_U82 ( .A1(U_ctl_n84), .A2(U_ctl_n318), .ZN(U_ctl_n78) );
  INV_X2 U_ctl_U81 ( .A(U_ctl_n290), .ZN(U_ctl_n190) );
  INV_X1 U_ctl_U79 ( .A(U_ctl_n306), .ZN(U_ctl_n301) );
  NOR2_X2 U_ctl_U78 ( .A1(U_ctl_n68), .A2(U_ctl_n219), .ZN(U_ctl_n164) );
  NAND2_X1 U_ctl_U77 ( .A1(U_ctl_n61), .A2(U_ctl_f_amba_bsz2[1]), .ZN(
        U_ctl_n59) );
  OAI21_X1 U_ctl_U76 ( .B1(U_ctl_n61), .B2(U_ctl_n289), .A(U_ctl_n59), .ZN(
        U_ctl_n224) );
  AND2_X1 U_ctl_U75 ( .A1(U_ctl_n189), .A2(U_ctl_n188), .ZN(U_ctl_n86) );
  AND2_X4 U_ctl_U74 ( .A1(U_ctl_n167), .A2(U_ctl_n200), .ZN(U_ctl_n47) );
  NAND2_X1 U_ctl_U73 ( .A1(U_ctl_n45), .A2(U_ctl_n44), .ZN(U_ctl_n104) );
  NAND2_X1 U_ctl_U72 ( .A1(U_ctl_n314), .A2(U_ctl_N284), .ZN(U_ctl_n45) );
  AOI222_X1 U_ctl_U71 ( .A1(U_ctl_fr_wr_bcnt_1_), .A2(U_ctl_n389), .B1(
        hiu_burst_size[1]), .B2(U_ctl_n388), .C1(U_ctl_n313), .C2(U_ctl_n43), 
        .ZN(U_ctl_n44) );
  XOR2_X1 U_ctl_U70 ( .A(U_ctl_DP_OP_140_125_8947_n14), .B(
        U_ctl_DP_OP_140_125_8947_n9), .Z(U_ctl_n43) );
  NOR2_X1 U_ctl_U69 ( .A1(U_ctl_n307), .A2(U_ctl_n42), .ZN(U_ctl_n_bh_state[0]) );
  AOI21_X1 U_ctl_U68 ( .B1(U_ctl_f_bh_state_0_), .B2(U_ctl_n344), .A(U_ctl_n41), .ZN(U_ctl_n42) );
  OAI22_X1 U_ctl_U67 ( .A1(U_ctl_n306), .A2(U_ctl_n397), .B1(m_rb_overflow), 
        .B2(U_ctl_n40), .ZN(U_ctl_n41) );
  NAND3_X1 U_ctl_U66 ( .A1(U_ctl_n305), .A2(U_ctl_n304), .A3(U_ctl_n39), .ZN(
        U_ctl_n40) );
  OAI22_X1 U_ctl_U65 ( .A1(U_ctl_n342), .A2(U_ctl_n95), .B1(miu_burst_done), 
        .B2(U_ctl_n38), .ZN(U_ctl_n39) );
  NOR2_X1 U_ctl_U64 ( .A1(U_ctl_f_bh_state_0_), .A2(U_ctl_n341), .ZN(U_ctl_n38) );
  AOI21_X1 U_ctl_U63 ( .B1(U_ctl_n84), .B2(U_ctl_n317), .A(U_ctl_n37), .ZN(
        U_ctl_n109) );
  NOR2_X1 U_ctl_U62 ( .A1(U_ctl_n84), .A2(U_ctl_n80), .ZN(U_ctl_n37) );
  OAI211_X1 U_ctl_U61 ( .C1(U_ctl_n148), .C2(U_ctl_n36), .A(U_ctl_n70), .B(
        U_ctl_n396), .ZN(U_ctl_n117) );
  AOI21_X1 U_ctl_U60 ( .B1(U_ctl_fd_amba_bcnt_1_), .B2(htrans[0]), .A(
        U_ctl_n395), .ZN(U_ctl_n36) );
  AOI21_X1 U_ctl_U59 ( .B1(U_ctl_n183), .B2(U_ctl_n400), .A(U_ctl_n289), .ZN(
        m_af_data1_in_13_) );
  XOR2_X1 U_ctl_U58 ( .A(U_ctl_fr_wr_bcnt_5_), .B(U_ctl_n35), .Z(U_ctl_N288)
         );
  NOR2_X1 U_ctl_U57 ( .A1(U_ctl_fr_wr_bcnt_4_), .A2(
        U_ctl_DP_OP_140_125_8947_n22), .ZN(U_ctl_n35) );
  OAI21_X1 U_ctl_U56 ( .B1(U_ctl_n280), .B2(U_ctl_n161), .A(U_ctl_n34), .ZN(
        U_ctl_n285) );
  NAND4_X1 U_ctl_U55 ( .A1(U_ctl_n282), .A2(hburst[2]), .A3(U_ctl_n284), .A4(
        U_ctl_n33), .ZN(U_ctl_n34) );
  OAI221_X1 U_ctl_U54 ( .B1(hburst[1]), .B2(U_ctl_n278), .C1(U_ctl_n275), .C2(
        U_ctl_n277), .A(U_ctl_n32), .ZN(U_ctl_n33) );
  OR2_X1 U_ctl_U53 ( .A1(U_ctl_n283), .A2(U_ctl_n279), .ZN(U_ctl_n32) );
  NAND2_X1 U_ctl_U51 ( .A1(U_ctl_n28), .A2(U_ctl_n30), .ZN(U_ctl_n103) );
  AOI222_X1 U_ctl_U50 ( .A1(U_ctl_fr_wr_bcnt_2_), .A2(U_ctl_n389), .B1(
        hiu_burst_size[2]), .B2(U_ctl_n388), .C1(U_ctl_n313), .C2(U_ctl_n29), 
        .ZN(U_ctl_n30) );
  XOR2_X1 U_ctl_U49 ( .A(U_ctl_DP_OP_140_125_8947_n7), .B(
        U_ctl_DP_OP_140_125_8947_n13), .Z(U_ctl_n29) );
  NAND2_X1 U_ctl_U48 ( .A1(U_ctl_n314), .A2(U_ctl_N285), .ZN(U_ctl_n28) );
  AOI221_X1 U_ctl_U47 ( .B1(U_ctl_n297), .B2(U_ctl_n26), .C1(U_ctl_n300), .C2(
        U_ctl_n26), .A(U_ctl_n307), .ZN(U_ctl_n_bh_state[1]) );
  OAI21_X1 U_ctl_U45 ( .B1(U_ctl_n301), .B2(U_ctl_f_bh_state_1_), .A(m_rb_busy), .ZN(U_ctl_n26) );
  AOI21_X1 U_ctl_U44 ( .B1(U_ctl_n84), .B2(U_ctl_n320), .A(U_ctl_n25), .ZN(
        U_ctl_n114) );
  NOR2_X1 U_ctl_U43 ( .A1(U_ctl_n84), .A2(U_ctl_f_offset_2_), .ZN(U_ctl_n25)
         );
  INV_X1 U_ctl_U42 ( .A(U_ctl_n24), .ZN(m_af_data2_in[6]) );
  AOI22_X1 U_ctl_U41 ( .A1(U_ctl_n150), .A2(U_ctl_n224), .B1(U_ctl_n183), .B2(
        U_ctl_n225), .ZN(U_ctl_n24) );
  NAND3_X1 U_ctl_U40 ( .A1(U_ctl_n337), .A2(hburst[2]), .A3(U_ctl_n338), .ZN(
        U_ctl_n70) );
  INV_X1 U_ctl_U39 ( .A(U_ctl_n23), .ZN(U_ctl_n53) );
  OAI211_X1 U_ctl_U38 ( .C1(U_ctl_n280), .C2(U_ctl_n143), .A(U_ctl_n261), .B(
        U_ctl_n22), .ZN(U_ctl_n23) );
  NAND3_X1 U_ctl_U37 ( .A1(U_ctl_n262), .A2(U_ctl_n260), .A3(U_ctl_n282), .ZN(
        U_ctl_n22) );
  NAND2_X1 U_ctl_U36 ( .A1(U_ctl_n19), .A2(U_ctl_n21), .ZN(U_ctl_n102) );
  AOI222_X1 U_ctl_U35 ( .A1(U_ctl_fr_wr_bcnt_3_), .A2(U_ctl_n389), .B1(
        hiu_burst_size[3]), .B2(U_ctl_n388), .C1(U_ctl_n313), .C2(U_ctl_n20), 
        .ZN(U_ctl_n21) );
  XOR2_X1 U_ctl_U34 ( .A(U_ctl_DP_OP_140_125_8947_n5), .B(
        U_ctl_DP_OP_140_125_8947_n12), .Z(U_ctl_n20) );
  NAND2_X1 U_ctl_U33 ( .A1(U_ctl_n314), .A2(U_ctl_N286), .ZN(U_ctl_n19) );
  OAI21_X1 U_ctl_U32 ( .B1(U_ctl_n163), .B2(U_ctl_n183), .A(U_ctl_n18), .ZN(
        m_af_data2_in[5]) );
  NAND2_X1 U_ctl_U31 ( .A1(U_ctl_n224), .A2(U_ctl_n183), .ZN(U_ctl_n18) );
  NAND3_X1 U_ctl_U29 ( .A1(U_ctl_fd_miu_col_width_3_), .A2(U_ctl_n99), .A3(
        U_ctl_n16), .ZN(U_ctl_n166) );
  INV_X1 U_ctl_U28 ( .A(haddr[8]), .ZN(U_ctl_n16) );
  NAND2_X1 U_ctl_U27 ( .A1(U_ctl_n13), .A2(U_ctl_n15), .ZN(U_ctl_n101) );
  AOI222_X1 U_ctl_U26 ( .A1(U_ctl_fr_wr_bcnt_4_), .A2(U_ctl_n389), .B1(
        hiu_burst_size[4]), .B2(U_ctl_n388), .C1(U_ctl_n313), .C2(U_ctl_n14), 
        .ZN(U_ctl_n15) );
  XOR2_X1 U_ctl_U25 ( .A(U_ctl_DP_OP_140_125_8947_n3), .B(
        U_ctl_DP_OP_140_125_8947_n11), .Z(U_ctl_n14) );
  NAND2_X1 U_ctl_U24 ( .A1(U_ctl_n314), .A2(U_ctl_N287), .ZN(U_ctl_n13) );
  NOR2_X2 U_ctl_U23 ( .A1(U_ctl_n50), .A2(U_ctl_n53), .ZN(m_af_data1_in_4_) );
  NOR2_X1 U_ctl_U22 ( .A1(U_ctl_n225), .A2(U_ctl_n183), .ZN(U_ctl_n89) );
  NOR2_X1 U_ctl_U20 ( .A1(U_ctl_n11), .A2(U_ctl_n221), .ZN(m_df_data_in[0]) );
  AOI22_X1 U_ctl_U19 ( .A1(m_rb_busy), .A2(U_ctl_fd_non_single), .B1(m_rb_done), .B2(U_ctl_n220), .ZN(U_ctl_n11) );
  NAND2_X1 U_ctl_U18 ( .A1(U_ctl_n10), .A2(U_ctl_n7), .ZN(U_ctl_n255) );
  NAND3_X1 U_ctl_U17 ( .A1(U_ctl_n8), .A2(U_ctl_n9), .A3(U_ctl_n269), .ZN(
        U_ctl_n10) );
  AOI22_X1 U_ctl_U16 ( .A1(U_ctl_f_offset_2_), .A2(U_ctl_n320), .B1(
        U_ctl_f_offset_1_), .B2(U_ctl_n265), .ZN(U_ctl_n9) );
  OAI21_X1 U_ctl_U15 ( .B1(U_ctl_n289), .B2(U_ctl_f_offset_1_), .A(
        U_ctl_f_offset_0_), .ZN(U_ctl_n8) );
  AOI22_X1 U_ctl_U14 ( .A1(haddr[4]), .A2(U_ctl_n157), .B1(haddr[5]), .B2(
        U_ctl_n74), .ZN(U_ctl_n7) );
  NOR2_X1 U_ctl_U13 ( .A1(miu_pop_n), .A2(U_ctl_n6), .ZN(U_ctl_n314) );
  NAND3_X1 U_ctl_U12 ( .A1(U_ctl_n144), .A2(U_ctl_n386), .A3(U_ctl_n310), .ZN(
        U_ctl_n6) );
  NAND4_X2 U_ctl_U11 ( .A1(U_ctl_n261), .A2(U_ctl_n258), .A3(n51), .A4(
        U_ctl_n5), .ZN(U_ctl_n280) );
  NAND3_X2 U_ctl_U10 ( .A1(U_ctl_n185), .A2(U_ctl_n64), .A3(U_ctl_n256), .ZN(
        U_ctl_n5) );
  NAND3_X1 U_ctl_U8 ( .A1(U_ctl_n3), .A2(m_rb_overflow), .A3(U_ctl_n305), .ZN(
        U_ctl_n306) );
  NAND2_X1 U_ctl_U7 ( .A1(U_ctl_n292), .A2(U_ctl_f_bh_state_0_), .ZN(U_ctl_n3)
         );
  NAND4_X1 U_ctl_U6 ( .A1(U_ctl_n167), .A2(U_ctl_n331), .A3(U_ctl_n244), .A4(
        U_ctl_n200), .ZN(U_ctl_n165) );
  DFFR_X2 U_ctl_f_hiu_terminate_reg ( .D(hiu_terminate), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_f_hiu_terminate), .QN(U_ctl_n144) );
  DFFR_X2 U_ctl_fr_wr_bcnt_reg_0_ ( .D(U_ctl_n105), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fr_wr_bcnt_0_), .QN(U_ctl_n97) );
  DFFR_X2 U_ctl_f_offset_reg_2_ ( .D(U_ctl_n114), .CK(hclk), .RN(hresetn), .Q(
        U_ctl_f_offset_2_), .QN(U_ctl_n157) );
  DFFR_X2 U_ctl_fd_miu_col_width_reg_2_ ( .D(U_ctl_n129), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_fd_miu_col_width_2_), .QN(U_ctl_n154) );
  DFFR_X2 U_ctl_fd_miu_col_width_reg_0_ ( .D(U_ctl_n131), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_fd_miu_col_width_0_), .QN(U_ctl_n99) );
  DFFR_X2 U_ctl_fd_miu_col_width_reg_1_ ( .D(U_ctl_n130), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_fd_miu_col_width_1_), .QN(U_ctl_n153) );
  DFFR_X2 U_ctl_fd_miu_data_width_reg_0_ ( .D(U_ctl_n123), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_fd_miu_data_width_0_), .QN(U_ctl_n147) );
  DFFR_X2 U_ctl_fd_amba_bcnt_reg_2_ ( .D(U_ctl_n117), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fd_amba_bcnt_2_), .QN(U_ctl_n148) );
  DFFR_X2 U_ctl_o_two_to_one_reg ( .D(U_ctl_n122), .CK(hclk), .RN(hresetn), 
        .Q(m_two_to_one), .QN(U_ctl_n96) );
  DFFR_X2 U_ctl_fd_wr_width_reg ( .D(U_ctl_n136), .CK(hclk), .RN(hresetn), .Q(
        U_ctl_fd_wr_width), .QN(U_ctl_n126) );
  DFFR_X2 U_ctl_fd_amba_bcnt_reg_0_ ( .D(U_ctl_n119), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fd_amba_bcnt_0_), .QN(U_ctl_n143) );
  DFFR_X2 U_ctl_fd_non_single_reg ( .D(U_ctl_n140), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fd_non_single), .QN(U_ctl_n160) );
  DFFR_X2 U_ctl_fd_narrow_trans_reg ( .D(U_ctl_n139), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fd_narrow_trans), .QN(U_ctl_n98) );
  DFFR_X2 U_ctl_fd_rd_bz_reg ( .D(U_ctl_n120), .CK(hclk), .RN(hresetn), .Q(
        U_ctl_fd_rd_bz), .QN(U_ctl_n146) );
  DFFR_X2 U_ctl_fd_incr_reg ( .D(U_ctl_n141), .CK(hclk), .RN(hresetn), .Q(
        U_ctl_fd_incr), .QN(U_ctl_n156) );
  DFFR_X2 U_ctl_fd_wr_bz_reg ( .D(U_ctl_n121), .CK(hclk), .RN(hresetn), .Q(
        U_ctl_fd_wr_bz), .QN(U_ctl_n62) );
  DFFR_X2 U_ctl_f_offset_reg_3_ ( .D(U_ctl_n115), .CK(hclk), .RN(hresetn), .Q(
        U_ctl_f_offset_3_), .QN(U_ctl_n74) );
  DFFR_X2 U_ctl_fd_amba_bcnt_reg_3_ ( .D(U_ctl_n116), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fd_amba_bcnt_3_), .QN(U_ctl_n161) );
  DFFR_X2 U_ctl_fd_double_reg ( .D(U_ctl_n124), .CK(hclk), .RN(hresetn), .Q(
        m_double), .QN(U_ctl_n324) );
  DFFR_X2 U_ctl_fd_amba_bcnt_reg_1_ ( .D(U_ctl_n118), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fd_amba_bcnt_1_), .QN(U_ctl_n145) );
  DFFR_X2 U_ctl_f_amba_bsz2_reg_0_ ( .D(U_ctl_n107), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_f_amba_bsz2[0]), .QN(U_ctl_n83) );
  DFFR_X2 U_ctl_f_offset_reg_0_ ( .D(U_ctl_n112), .CK(hclk), .RN(hresetn), .Q(
        U_ctl_f_offset_0_), .QN(U_ctl_n77) );
  DFFR_X2 U_ctl_f_amba_bsz2_reg_1_ ( .D(U_ctl_n108), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_f_amba_bsz2[1]), .QN(U_ctl_n81) );
  DFFR_X2 U_ctl_f_offset_reg_1_ ( .D(U_ctl_n113), .CK(hclk), .RN(hresetn), .Q(
        U_ctl_f_offset_1_), .QN(U_ctl_n76) );
  DFFR_X2 U_ctl_f_amba_bsz2_reg_3_ ( .D(U_ctl_n110), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_f_amba_bsz2[3]), .QN(U_ctl_n79) );
  DFFR_X2 U_ctl_fd_miu_col_width_reg_3_ ( .D(U_ctl_n128), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_fd_miu_col_width_3_) );
  DFFR_X2 U_ctl_fr_prv_1wrap_reg ( .D(U_ctl_N236), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fr_prv_1wrap) );
  DFFR_X2 U_ctl_f_col_width_reg_2_ ( .D(U_ctl_n133), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_f_col_width[2]) );
  DFFR_X2 U_ctl_fd_miu_data_width_reg_1_ ( .D(U_ctl_n125), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_fd_miu_data_width_1_) );
  DFFR_X2 U_ctl_fd_haddr_reg_1_ ( .D(U_ctl_n137), .CK(hclk), .RN(hresetn), .Q(
        U_ctl_fd_haddr_1_) );
  DFFR_X2 U_ctl_f_burst_done2_reg ( .D(U_ctl_f_burst_done), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_f_burst_done2) );
  DFFR_X2 U_ctl_f_amba_bsz2_reg_2_ ( .D(U_ctl_n109), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_n80), .QN(U_ctl_n188) );
  DFFR_X2 U_ctl_f_wrap_burst_reg ( .D(U_ctl_n111), .CK(hclk), .RN(hresetn), 
        .QN(U_ctl_n159) );
  DFFR_X2 U_ctl_fd_reg_access_reg ( .D(U_ctl_n138), .CK(hclk), .RN(hresetn), 
        .QN(U_ctl_n158) );
  INV_X2 U_ctl_DP_OP_140_125_8947_U31 ( .A(U_ctl_DP_OP_140_125_8947_n20), .ZN(
        U_ctl_DP_OP_140_125_8947_n30) );
  XNOR2_X1 U_ctl_DP_OP_140_125_8947_U38 ( .A(U_ctl_DP_OP_140_125_8947_n24), 
        .B(U_ctl_fr_wr_bcnt_2_), .ZN(U_ctl_N285) );
  XOR2_X1 U_ctl_DP_OP_140_125_8947_U2 ( .A(hiu_burst_size[5]), .B(
        U_ctl_DP_OP_140_125_8947_n35), .Z(U_ctl_DP_OP_140_125_8947_n1) );
  XOR2_X1 U_ctl_DP_OP_140_125_8947_U19 ( .A(hiu_burst_size[0]), .B(
        U_ctl_DP_OP_140_125_8947_n30), .Z(U_ctl_C64_DATA2_0) );
  INV_X2 U_ctl_DP_OP_140_125_8947_U21 ( .A(U_ctl_DP_OP_140_125_8947_n15), .ZN(
        U_ctl_DP_OP_140_125_8947_n35) );
  OR2_X2 U_ctl_DP_OP_140_125_8947_U37 ( .A1(U_ctl_DP_OP_140_125_8947_n23), 
        .A2(U_ctl_fr_wr_bcnt_3_), .ZN(U_ctl_DP_OP_140_125_8947_n22) );
  XNOR2_X1 U_ctl_DP_OP_140_125_8947_U36 ( .A(U_ctl_DP_OP_140_125_8947_n23), 
        .B(U_ctl_fr_wr_bcnt_3_), .ZN(U_ctl_N286) );
  OR2_X2 U_ctl_DP_OP_140_125_8947_U39 ( .A1(U_ctl_DP_OP_140_125_8947_n24), 
        .A2(U_ctl_fr_wr_bcnt_2_), .ZN(U_ctl_DP_OP_140_125_8947_n23) );
  OR2_X2 U_ctl_DP_OP_140_125_8947_U41 ( .A1(U_ctl_fr_wr_bcnt_0_), .A2(
        U_ctl_fr_wr_bcnt_1_), .ZN(U_ctl_DP_OP_140_125_8947_n24) );
  AOI22_X1 U_ctl_DP_OP_140_125_8947_U24 ( .A1(U_ctl_N287), .A2(
        U_ctl_DP_OP_140_125_8947_I2), .B1(miu_pop_n), .B2(U_ctl_fr_wr_bcnt_4_), 
        .ZN(U_ctl_DP_OP_140_125_8947_n16) );
  AOI22_X1 U_ctl_DP_OP_140_125_8947_U26 ( .A1(U_ctl_N286), .A2(
        U_ctl_DP_OP_140_125_8947_I2), .B1(miu_pop_n), .B2(U_ctl_fr_wr_bcnt_3_), 
        .ZN(U_ctl_DP_OP_140_125_8947_n17) );
  AOI22_X1 U_ctl_DP_OP_140_125_8947_U28 ( .A1(U_ctl_N285), .A2(
        U_ctl_DP_OP_140_125_8947_I2), .B1(miu_pop_n), .B2(U_ctl_fr_wr_bcnt_2_), 
        .ZN(U_ctl_DP_OP_140_125_8947_n18) );
  AOI22_X1 U_ctl_DP_OP_140_125_8947_U32 ( .A1(U_ctl_n97), .A2(
        U_ctl_DP_OP_140_125_8947_I2), .B1(miu_pop_n), .B2(U_ctl_fr_wr_bcnt_0_), 
        .ZN(U_ctl_DP_OP_140_125_8947_n20) );
  AOI22_X1 U_ctl_DP_OP_140_125_8947_U30 ( .A1(U_ctl_N284), .A2(
        U_ctl_DP_OP_140_125_8947_I2), .B1(miu_pop_n), .B2(U_ctl_fr_wr_bcnt_1_), 
        .ZN(U_ctl_DP_OP_140_125_8947_n19) );
  AOI22_X1 U_ctl_DP_OP_140_125_8947_U22 ( .A1(U_ctl_N288), .A2(
        U_ctl_DP_OP_140_125_8947_I2), .B1(miu_pop_n), .B2(U_ctl_fr_wr_bcnt_5_), 
        .ZN(U_ctl_DP_OP_140_125_8947_n15) );
  INV_X4 U_ctl_DP_OP_140_125_8947_U4 ( .A(U_ctl_DP_OP_140_125_8947_n2), .ZN(
        U_ctl_DP_OP_140_125_8947_n10) );
  AOI22_X2 U_ctl_DP_OP_140_125_8947_U5 ( .A1(U_ctl_DP_OP_140_125_8947_n11), 
        .A2(U_ctl_DP_OP_140_125_8947_n3), .B1(U_ctl_DP_OP_140_125_8947_n34), 
        .B2(hiu_burst_size[4]), .ZN(U_ctl_DP_OP_140_125_8947_n2) );
  INV_X4 U_ctl_DP_OP_140_125_8947_U23 ( .A(U_ctl_DP_OP_140_125_8947_n16), .ZN(
        U_ctl_DP_OP_140_125_8947_n34) );
  INV_X4 U_ctl_DP_OP_140_125_8947_U8 ( .A(U_ctl_DP_OP_140_125_8947_n4), .ZN(
        U_ctl_DP_OP_140_125_8947_n11) );
  AOI22_X2 U_ctl_DP_OP_140_125_8947_U9 ( .A1(U_ctl_DP_OP_140_125_8947_n12), 
        .A2(U_ctl_DP_OP_140_125_8947_n5), .B1(U_ctl_DP_OP_140_125_8947_n33), 
        .B2(hiu_burst_size[3]), .ZN(U_ctl_DP_OP_140_125_8947_n4) );
  INV_X4 U_ctl_DP_OP_140_125_8947_U25 ( .A(U_ctl_DP_OP_140_125_8947_n17), .ZN(
        U_ctl_DP_OP_140_125_8947_n33) );
  INV_X4 U_ctl_DP_OP_140_125_8947_U12 ( .A(U_ctl_DP_OP_140_125_8947_n6), .ZN(
        U_ctl_DP_OP_140_125_8947_n12) );
  AOI22_X2 U_ctl_DP_OP_140_125_8947_U13 ( .A1(U_ctl_DP_OP_140_125_8947_n13), 
        .A2(U_ctl_DP_OP_140_125_8947_n7), .B1(U_ctl_DP_OP_140_125_8947_n32), 
        .B2(hiu_burst_size[2]), .ZN(U_ctl_DP_OP_140_125_8947_n6) );
  INV_X4 U_ctl_DP_OP_140_125_8947_U27 ( .A(U_ctl_DP_OP_140_125_8947_n18), .ZN(
        U_ctl_DP_OP_140_125_8947_n32) );
  INV_X4 U_ctl_DP_OP_140_125_8947_U16 ( .A(U_ctl_DP_OP_140_125_8947_n8), .ZN(
        U_ctl_DP_OP_140_125_8947_n13) );
  AOI22_X2 U_ctl_DP_OP_140_125_8947_U17 ( .A1(U_ctl_DP_OP_140_125_8947_n9), 
        .A2(U_ctl_DP_OP_140_125_8947_n14), .B1(U_ctl_DP_OP_140_125_8947_n31), 
        .B2(hiu_burst_size[1]), .ZN(U_ctl_DP_OP_140_125_8947_n8) );
  INV_X4 U_ctl_DP_OP_140_125_8947_U29 ( .A(U_ctl_DP_OP_140_125_8947_n19), .ZN(
        U_ctl_DP_OP_140_125_8947_n31) );
  DFFS_X2 U_ctl_fd_hsel_mem_reg ( .D(U_ctl_n63), .CK(hclk), .SN(hresetn), .Q(
        U_ctl_n155), .QN(U_ctl_fd_hsel_mem) );
  XOR2_X2 U_ctl_DP_OP_140_125_8947_U1 ( .A(U_ctl_DP_OP_140_125_8947_n1), .B(
        U_ctl_DP_OP_140_125_8947_n10), .Z(U_ctl_C64_DATA2_5) );
  XOR2_X2 U_ctl_DP_OP_140_125_8947_U6 ( .A(hiu_burst_size[4]), .B(
        U_ctl_DP_OP_140_125_8947_n34), .Z(U_ctl_DP_OP_140_125_8947_n3) );
  XOR2_X2 U_ctl_DP_OP_140_125_8947_U10 ( .A(hiu_burst_size[3]), .B(
        U_ctl_DP_OP_140_125_8947_n33), .Z(U_ctl_DP_OP_140_125_8947_n5) );
  XOR2_X2 U_ctl_DP_OP_140_125_8947_U14 ( .A(hiu_burst_size[2]), .B(
        U_ctl_DP_OP_140_125_8947_n32), .Z(U_ctl_DP_OP_140_125_8947_n7) );
  XOR2_X2 U_ctl_DP_OP_140_125_8947_U18 ( .A(hiu_burst_size[1]), .B(
        U_ctl_DP_OP_140_125_8947_n31), .Z(U_ctl_DP_OP_140_125_8947_n9) );
  AND2_X4 U_ctl_DP_OP_140_125_8947_U20 ( .A1(U_ctl_DP_OP_140_125_8947_n30), 
        .A2(hiu_burst_size[0]), .ZN(U_ctl_DP_OP_140_125_8947_n14) );
  XNOR2_X2 U_ctl_DP_OP_140_125_8947_U34 ( .A(U_ctl_DP_OP_140_125_8947_n22), 
        .B(U_ctl_fr_wr_bcnt_4_), .ZN(U_ctl_N287) );
  XNOR2_X2 U_ctl_DP_OP_140_125_8947_U40 ( .A(U_ctl_fr_wr_bcnt_0_), .B(
        U_ctl_fr_wr_bcnt_1_), .ZN(U_ctl_N284) );
  DFFR_X1 U_ctl_f_sel_buf_reg ( .D(U_ctl_n_sel_buf), .CK(hclk), .RN(hresetn), 
        .Q(m_rb_sel_buf), .QN(n48) );
  DFFR_X1 U_ctl_f_bh_state_reg_1_ ( .D(U_ctl_n_bh_state[1]), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_f_bh_state_1_) );
  DFFR_X1 U_ctl_fr_prv_1wrap_tm_reg ( .D(U_ctl_N237), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fr_prv_1wrap_tm) );
  DFFR_X1 U_ctl_f_bh_state_reg_2_ ( .D(U_ctl_n_bh_state[2]), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_f_bh_state_2_), .QN(U_ctl_n142) );
  DFFR_X1 U_ctl_f_bh_state_reg_0_ ( .D(U_ctl_n_bh_state[0]), .CK(hclk), .RN(
        hresetn), .Q(U_ctl_f_bh_state_0_), .QN(U_ctl_n95) );
  DFFR_X1 U_ctl_fr_wr_bcnt_reg_5_ ( .D(U_ctl_n100), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fr_wr_bcnt_5_) );
  DFFR_X1 U_ctl_fr_wr_bcnt_reg_4_ ( .D(U_ctl_n101), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fr_wr_bcnt_4_) );
  DFFR_X1 U_ctl_fr_wr_bcnt_reg_3_ ( .D(U_ctl_n102), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fr_wr_bcnt_3_) );
  DFFR_X1 U_ctl_fr_wr_bcnt_reg_2_ ( .D(U_ctl_n103), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fr_wr_bcnt_2_) );
  DFFR_X1 U_ctl_fr_wr_bcnt_reg_1_ ( .D(U_ctl_n104), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_fr_wr_bcnt_1_) );
  DFFR_X1 U_ctl_f_burst_done_reg ( .D(miu_burst_done), .CK(hclk), .RN(hresetn), 
        .Q(U_ctl_f_burst_done) );
  DFFS_X2 U_ctl_fd_rd_ready_reg ( .D(U_ctl_n106), .CK(hclk), .SN(hresetn), .Q(
        U_ctl_fd_rd_ready) );
  DFFS_X2 U_ctl_fd_df_push_n_reg ( .D(U_ctl_n299), .CK(hclk), .SN(hresetn), 
        .QN(m_df_push_n) );
  DFFS_X2 U_ctl_fd_zero_wait_ok_reg ( .D(U_ctl_N89), .CK(hclk), .SN(hresetn), 
        .QN(U_ctl_n151) );
  DFFS_X2 U_ctl_f_data_width_reg_0_ ( .D(U_ctl_n127), .CK(hclk), .SN(hresetn), 
        .Q(U_ctl_f_data_width_0_) );
  DFFS_X2 U_ctl_f_col_width_reg_3_ ( .D(U_ctl_n132), .CK(hclk), .SN(hresetn), 
        .Q(U_ctl_f_col_width[3]) );
  DFFS_X2 U_ctl_f_col_width_reg_1_ ( .D(U_ctl_n134), .CK(hclk), .SN(hresetn), 
        .Q(U_ctl_f_col_width[1]) );
  DFFS_X2 U_ctl_f_col_width_reg_0_ ( .D(U_ctl_n135), .CK(hclk), .SN(hresetn), 
        .Q(U_ctl_f_col_width[0]) );
  MUX2_X2 U_afifo_U_acore_U191 ( .A(U_afifo_U_acore_f_obuf_41_), .B(
        U_afifo_U_acore_f_ibuf_41_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[31])
         );
  MUX2_X2 U_afifo_U_acore_U190 ( .A(U_afifo_U_acore_f_obuf_40_), .B(
        U_afifo_U_acore_f_ibuf_40_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[30])
         );
  MUX2_X2 U_afifo_U_acore_U189 ( .A(U_afifo_U_acore_f_obuf_39_), .B(
        U_afifo_U_acore_f_ibuf_39_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[29])
         );
  MUX2_X2 U_afifo_U_acore_U188 ( .A(U_afifo_U_acore_f_obuf_38_), .B(
        U_afifo_U_acore_f_ibuf_38_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[28])
         );
  MUX2_X2 U_afifo_U_acore_U187 ( .A(U_afifo_U_acore_f_obuf_37_), .B(
        U_afifo_U_acore_f_ibuf_37_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[27])
         );
  MUX2_X2 U_afifo_U_acore_U186 ( .A(U_afifo_U_acore_f_obuf_36_), .B(
        U_afifo_U_acore_f_ibuf_36_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[26])
         );
  MUX2_X2 U_afifo_U_acore_U185 ( .A(U_afifo_U_acore_f_obuf_35_), .B(
        U_afifo_U_acore_f_ibuf_35_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[25])
         );
  MUX2_X2 U_afifo_U_acore_U184 ( .A(U_afifo_U_acore_f_obuf_34_), .B(
        U_afifo_U_acore_f_ibuf_34_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[24])
         );
  MUX2_X2 U_afifo_U_acore_U183 ( .A(U_afifo_U_acore_f_obuf_33_), .B(
        U_afifo_U_acore_f_ibuf_33_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[23])
         );
  MUX2_X2 U_afifo_U_acore_U182 ( .A(U_afifo_U_acore_f_obuf_32_), .B(
        U_afifo_U_acore_f_ibuf_32_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[22])
         );
  MUX2_X2 U_afifo_U_acore_U181 ( .A(U_afifo_U_acore_f_obuf_31_), .B(
        U_afifo_U_acore_f_ibuf_31_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[21])
         );
  MUX2_X2 U_afifo_U_acore_U180 ( .A(U_afifo_U_acore_f_obuf_30_), .B(
        U_afifo_U_acore_f_ibuf_30_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[20])
         );
  MUX2_X2 U_afifo_U_acore_U179 ( .A(U_afifo_U_acore_f_obuf_18_), .B(
        U_afifo_U_acore_f_ibuf_18_), .S(U_afifo_U_acore_n1), .Z(hiu_addr[8])
         );
  MUX2_X2 U_afifo_U_acore_U178 ( .A(U_afifo_U_acore_f_obuf_2_), .B(
        U_afifo_U_acore_f_ibuf_2_), .S(U_afifo_U_acore_n1), .Z(hiu_rw) );
  INV_X4 U_afifo_U_acore_U177 ( .A(U_afifo_m_pop_n), .ZN(U_afifo_U_acore_n45)
         );
  OAI22_X1 U_afifo_U_acore_U176 ( .A1(U_afifo_U_acore_n168), .A2(
        U_afifo_U_acore_n35), .B1(U_afifo_m_pop_n), .B2(U_afifo_U_acore_n170), 
        .ZN(U_afifo_U_acore_n_obuf_empty) );
  INV_X4 U_afifo_U_acore_U175 ( .A(U_afifo_U_acore_n211), .ZN(
        U_afifo_U_acore_n42) );
  OAI21_X2 U_afifo_U_acore_U174 ( .B1(U_afifo_U_acore_n100), .B2(
        U_afifo_U_acore_n35), .A(U_afifo_U_acore_n60), .ZN(hiu_addr[16]) );
  OAI21_X2 U_afifo_U_acore_U173 ( .B1(U_afifo_U_acore_n156), .B2(
        U_afifo_U_acore_n37), .A(U_afifo_U_acore_n56), .ZN(hiu_addr[12]) );
  OAI21_X2 U_afifo_U_acore_U172 ( .B1(U_afifo_U_acore_n153), .B2(
        U_afifo_U_acore_n37), .A(U_afifo_U_acore_n57), .ZN(hiu_addr[13]) );
  OAI21_X2 U_afifo_U_acore_U171 ( .B1(U_afifo_U_acore_n160), .B2(
        U_afifo_U_acore_n35), .A(U_afifo_U_acore_n54), .ZN(hiu_addr[10]) );
  NOR2_X2 U_afifo_U_acore_U170 ( .A1(U_afifo_U_acore_n45), .A2(
        U_afifo_U_acore_n44), .ZN(U_afifo_U_acore_n49) );
  OAI211_X2 U_afifo_U_acore_U169 ( .C1(U_afifo_m_pop_n), .C2(
        U_afifo_U_acore_n64), .A(U_afifo_U_acore_n169), .B(U_afifo_U_acore_n11), .ZN(U_afifo_U_acore_n165) );
  OAI21_X1 U_afifo_U_acore_U168 ( .B1(U_afifo_U_acore_n166), .B2(
        U_afifo_U_acore_n11), .A(U_afifo_U_acore_f_afull), .ZN(
        U_afifo_U_acore_n65) );
  OAI21_X2 U_afifo_U_acore_U167 ( .B1(U_afifo_U_acore_n102), .B2(
        U_afifo_U_acore_n37), .A(U_afifo_U_acore_n59), .ZN(hiu_addr[15]) );
  NAND2_X2 U_afifo_U_acore_U166 ( .A1(U_afifo_U_acore_n2), .A2(
        U_afifo_U_acore_n1), .ZN(U_afifo_U_acore_n169) );
  OAI21_X2 U_afifo_U_acore_U165 ( .B1(U_afifo_U_acore_n162), .B2(
        U_afifo_U_acore_n35), .A(U_afifo_U_acore_n53), .ZN(hiu_addr[9]) );
  NOR2_X2 U_afifo_U_acore_U164 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_f_push_req_n), .ZN(U_afifo_U_acore_n46) );
  INV_X8 U_afifo_U_acore_U163 ( .A(U_afifo_U_acore_n34), .ZN(
        U_afifo_U_acore_n43) );
  INV_X4 U_afifo_U_acore_U162 ( .A(U_afifo_U_acore_n38), .ZN(
        U_afifo_U_acore_n36) );
  NAND2_X2 U_afifo_U_acore_U161 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_26_), .ZN(U_afifo_U_acore_n60) );
  NAND2_X2 U_afifo_U_acore_U160 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_25_), .ZN(U_afifo_U_acore_n59) );
  NAND2_X2 U_afifo_U_acore_U159 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_27_), .ZN(U_afifo_U_acore_n61) );
  OAI21_X2 U_afifo_U_acore_U158 ( .B1(U_afifo_U_acore_n98), .B2(
        U_afifo_U_acore_n35), .A(U_afifo_U_acore_n61), .ZN(hiu_addr[17]) );
  NAND2_X2 U_afifo_U_acore_U157 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_28_), .ZN(U_afifo_U_acore_n62) );
  OAI21_X2 U_afifo_U_acore_U156 ( .B1(U_afifo_U_acore_n96), .B2(
        U_afifo_U_acore_n35), .A(U_afifo_U_acore_n62), .ZN(hiu_addr[18]) );
  OAI21_X2 U_afifo_U_acore_U155 ( .B1(U_afifo_U_acore_n94), .B2(
        U_afifo_U_acore_n43), .A(U_afifo_U_acore_n63), .ZN(hiu_addr[19]) );
  NAND2_X2 U_afifo_U_acore_U154 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_22_), .ZN(U_afifo_U_acore_n56) );
  NAND2_X2 U_afifo_U_acore_U153 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_23_), .ZN(U_afifo_U_acore_n57) );
  NAND2_X2 U_afifo_U_acore_U152 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_21_), .ZN(U_afifo_U_acore_n55) );
  NAND2_X2 U_afifo_U_acore_U151 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_24_), .ZN(U_afifo_U_acore_n58) );
  NOR2_X2 U_afifo_U_acore_U150 ( .A1(U_afifo_U_acore_n11), .A2(
        U_afifo_U_acore_n169), .ZN(U_afifo_m_empty) );
  INV_X4 U_afifo_U_acore_U149 ( .A(U_afifo_U_acore_n2), .ZN(
        U_afifo_U_acore_n64) );
  NAND2_X2 U_afifo_U_acore_U148 ( .A1(U_afifo_U_acore_n64), .A2(
        U_afifo_U_acore_n11), .ZN(U_afifo_U_acore_n66) );
  NAND2_X2 U_afifo_U_acore_U147 ( .A1(U_afifo_U_acore_n66), .A2(
        U_afifo_U_acore_n12), .ZN(U_afifo_m_afull) );
  NAND2_X2 U_afifo_U_acore_U146 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_20_), .ZN(U_afifo_U_acore_n54) );
  NAND2_X2 U_afifo_U_acore_U145 ( .A1(U_afifo_U_acore_n37), .A2(
        U_afifo_U_acore_f_obuf_19_), .ZN(U_afifo_U_acore_n53) );
  NOR2_X2 U_afifo_U_acore_U144 ( .A1(U_afifo_U_acore_n64), .A2(
        U_afifo_U_acore_n46), .ZN(U_afifo_m_aempty) );
  AOI22_X2 U_afifo_U_acore_U143 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_18_), .B1(U_afifo_U_acore_m_sf_data_out[18]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n164) );
  AOI22_X2 U_afifo_U_acore_U142 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_28_), .B1(U_afifo_U_acore_m_sf_data_out[28]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n95) );
  AOI22_X2 U_afifo_U_acore_U141 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_27_), .B1(U_afifo_U_acore_m_sf_data_out[27]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n97) );
  AOI22_X2 U_afifo_U_acore_U140 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_25_), .B1(U_afifo_U_acore_m_sf_data_out[25]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n101) );
  AOI22_X2 U_afifo_U_acore_U139 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_29_), .B1(U_afifo_U_acore_m_sf_data_out[29]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n93) );
  AOI22_X2 U_afifo_U_acore_U138 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_26_), .B1(U_afifo_U_acore_m_sf_data_out[26]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n99) );
  AOI22_X2 U_afifo_U_acore_U137 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_24_), .B1(U_afifo_U_acore_m_sf_data_out[24]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n103) );
  AOI22_X2 U_afifo_U_acore_U136 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_23_), .B1(U_afifo_U_acore_m_sf_data_out[23]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n143) );
  AOI22_X2 U_afifo_U_acore_U135 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_22_), .B1(U_afifo_U_acore_m_sf_data_out[22]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n155) );
  AOI22_X2 U_afifo_U_acore_U134 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_20_), .B1(U_afifo_U_acore_m_sf_data_out[20]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n159) );
  AOI22_X2 U_afifo_U_acore_U133 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_19_), .B1(U_afifo_U_acore_m_sf_data_out[19]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n161) );
  AOI22_X2 U_afifo_U_acore_U132 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_21_), .B1(U_afifo_U_acore_m_sf_data_out[21]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n157) );
  AOI22_X2 U_afifo_U_acore_U131 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_37_), .B1(U_afifo_U_acore_m_sf_data_out[37]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n75) );
  AOI22_X2 U_afifo_U_acore_U130 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_36_), .B1(U_afifo_U_acore_m_sf_data_out[36]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n77) );
  AOI22_X2 U_afifo_U_acore_U129 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_38_), .B1(U_afifo_U_acore_m_sf_data_out[38]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n73) );
  AOI22_X2 U_afifo_U_acore_U128 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_39_), .B1(U_afifo_U_acore_m_sf_data_out[39]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n71) );
  AOI22_X2 U_afifo_U_acore_U127 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_17_), .B1(U_afifo_U_acore_m_sf_data_out[17]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n196) );
  AOI22_X2 U_afifo_U_acore_U126 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_16_), .B1(U_afifo_U_acore_m_sf_data_out[16]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n198) );
  AOI22_X2 U_afifo_U_acore_U125 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_15_), .B1(U_afifo_U_acore_m_sf_data_out[15]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n200) );
  AOI22_X2 U_afifo_U_acore_U124 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_14_), .B1(U_afifo_U_acore_m_sf_data_out[14]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n202) );
  AOI22_X2 U_afifo_U_acore_U123 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_0_), .B1(U_afifo_U_acore_m_sf_data_out[0]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n209) );
  AOI22_X2 U_afifo_U_acore_U122 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_13_), .B1(U_afifo_U_acore_m_sf_data_out[13]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n204) );
  AOI22_X2 U_afifo_U_acore_U121 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_12_), .B1(U_afifo_U_acore_m_sf_data_out[12]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n206) );
  AOI22_X2 U_afifo_U_acore_U120 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_43_), .B1(U_afifo_U_acore_m_sf_data_out[43]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n191) );
  AOI22_X2 U_afifo_U_acore_U119 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_11_), .B1(U_afifo_U_acore_m_sf_data_out[11]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n208) );
  AOI22_X2 U_afifo_U_acore_U118 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_46_), .B1(U_afifo_U_acore_m_sf_data_out[46]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n187) );
  AOI22_X2 U_afifo_U_acore_U117 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_47_), .B1(U_afifo_U_acore_m_sf_data_out[47]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n185) );
  AOI22_X2 U_afifo_U_acore_U116 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_42_), .B1(U_afifo_U_acore_m_sf_data_out[42]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n193) );
  AOI22_X2 U_afifo_U_acore_U115 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_3_), .B1(U_afifo_U_acore_m_sf_data_out[3]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n195) );
  AOI22_X2 U_afifo_U_acore_U114 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_5_), .B1(U_afifo_U_acore_m_sf_data_out[5]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n178) );
  AOI22_X2 U_afifo_U_acore_U113 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_44_), .B1(U_afifo_U_acore_m_sf_data_out[44]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n189) );
  AOI22_X2 U_afifo_U_acore_U112 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_4_), .B1(U_afifo_U_acore_m_sf_data_out[4]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n180) );
  AOI22_X2 U_afifo_U_acore_U111 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_9_), .B1(U_afifo_U_acore_m_sf_data_out[9]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n171) );
  AOI22_X2 U_afifo_U_acore_U110 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_45_), .B1(U_afifo_U_acore_m_sf_data_out[45]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n188) );
  AOI22_X2 U_afifo_U_acore_U109 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_48_), .B1(U_afifo_U_acore_m_sf_data_out[48]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n183) );
  AOI22_X2 U_afifo_U_acore_U108 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_7_), .B1(U_afifo_U_acore_m_sf_data_out[7]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n174) );
  AOI22_X2 U_afifo_U_acore_U107 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_49_), .B1(U_afifo_U_acore_m_sf_data_out[49]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n182) );
  AOI22_X2 U_afifo_U_acore_U106 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_6_), .B1(U_afifo_U_acore_m_sf_data_out[6]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n176) );
  AOI22_X2 U_afifo_U_acore_U105 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_8_), .B1(U_afifo_U_acore_m_sf_data_out[8]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n172) );
  AOI22_X2 U_afifo_U_acore_U104 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_41_), .B1(U_afifo_U_acore_m_sf_data_out[41]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n67) );
  AOI22_X2 U_afifo_U_acore_U103 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_40_), .B1(U_afifo_U_acore_m_sf_data_out[40]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n69) );
  AOI22_X2 U_afifo_U_acore_U102 ( .A1(U_afifo_U_acore_n39), .A2(
        U_afifo_U_acore_f_obuf_2_), .B1(U_afifo_U_acore_m_sf_data_out[2]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n91) );
  OAI211_X1 U_afifo_U_acore_U101 ( .C1(U_afifo_U_acore_n45), .C2(
        U_afifo_U_acore_n66), .A(U_afifo_U_acore_n65), .B(
        U_afifo_U_acore_m_sf_full), .ZN(U_afifo_U_acore_n_afull) );
  INV_X8 U_afifo_U_acore_U100 ( .A(U_afifo_U_acore_n36), .ZN(
        U_afifo_U_acore_n37) );
  INV_X4 U_afifo_U_acore_U99 ( .A(U_afifo_U_acore_n166), .ZN(
        U_afifo_U_acore_n163) );
  OAI21_X2 U_afifo_U_acore_U96 ( .B1(U_afifo_U_acore_n1), .B2(
        U_afifo_U_acore_n7), .A(U_afifo_U_acore_n51), .ZN(hiu_burst_size[3])
         );
  INV_X4 U_afifo_U_acore_U95 ( .A(U_afifo_U_acore_n36), .ZN(
        U_afifo_U_acore_n35) );
  NOR2_X2 U_afifo_U_acore_U94 ( .A1(U_afifo_U_acore_n49), .A2(
        U_afifo_U_acore_n48), .ZN(U_afifo_U_acore_n168) );
  NAND2_X2 U_afifo_U_acore_U93 ( .A1(U_afifo_U_acore_n168), .A2(
        U_afifo_U_acore_n2), .ZN(U_afifo_U_acore_n211) );
  INV_X32 U_afifo_U_acore_U92 ( .A(U_afifo_U_acore_n43), .ZN(
        U_afifo_U_acore_n1) );
  OAI21_X1 U_afifo_U_acore_U91 ( .B1(U_afifo_U_acore_f_push_req_n), .B2(
        U_afifo_U_acore_n12), .A(U_afifo_U_acore_m_sf_full), .ZN(
        U_afifo_m_full) );
  NAND2_X1 U_afifo_U_acore_U90 ( .A1(U_afifo_U_acore_n2), .A2(
        U_afifo_U_acore_f_push_req_n), .ZN(U_afifo_U_acore_n170) );
  OR2_X2 U_afifo_U_acore_U89 ( .A1(U_afifo_U_acore_n175), .A2(
        U_afifo_U_acore_n35), .ZN(U_afifo_U_acore_n51) );
  NOR2_X1 U_afifo_U_acore_U86 ( .A1(U_afifo_U_acore_f_push_req_n), .A2(
        U_afifo_U_acore_n169), .ZN(U_afifo_U_acore_n44) );
  NOR2_X1 U_afifo_U_acore_U85 ( .A1(U_afifo_m_pop_n), .A2(U_afifo_U_acore_n47), 
        .ZN(U_afifo_U_acore_n48) );
  NAND2_X2 U_afifo_U_acore_U84 ( .A1(U_afifo_U_acore_n64), .A2(
        U_afifo_U_acore_n45), .ZN(U_afifo_U_acore_n166) );
  INV_X4 U_afifo_U_acore_U83 ( .A(U_afifo_U_acore_n168), .ZN(
        U_afifo_U_acore_n39) );
  INV_X4 U_afifo_U_acore_U82 ( .A(U_afifo_U_acore_n168), .ZN(
        U_afifo_U_acore_n40) );
  INV_X4 U_afifo_U_acore_U81 ( .A(U_afifo_U_acore_n42), .ZN(
        U_afifo_U_acore_n41) );
  OAI21_X1 U_afifo_U_acore_U80 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n190), .A(U_afifo_U_acore_n189), .ZN(
        U_afifo_U_acore_n116) );
  OAI21_X1 U_afifo_U_acore_U79 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n207), .A(U_afifo_U_acore_n206), .ZN(
        U_afifo_U_acore_n151) );
  OAI21_X1 U_afifo_U_acore_U78 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n199), .A(U_afifo_U_acore_n198), .ZN(
        U_afifo_U_acore_n147) );
  OAI21_X1 U_afifo_U_acore_U77 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n192), .A(U_afifo_U_acore_n191), .ZN(
        U_afifo_U_acore_n117) );
  OAI21_X1 U_afifo_U_acore_U76 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n210), .A(U_afifo_U_acore_n209), .ZN(
        U_afifo_U_acore_n154) );
  OAI21_X1 U_afifo_U_acore_U75 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n181), .A(U_afifo_U_acore_n180), .ZN(
        U_afifo_U_acore_n110) );
  OAI21_X1 U_afifo_U_acore_U74 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n203), .A(U_afifo_U_acore_n202), .ZN(
        U_afifo_U_acore_n149) );
  OAI21_X1 U_afifo_U_acore_U73 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n31), .A(U_afifo_U_acore_n208), .ZN(
        U_afifo_U_acore_n152) );
  OAI21_X1 U_afifo_U_acore_U72 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n179), .A(U_afifo_U_acore_n178), .ZN(
        U_afifo_U_acore_n109) );
  OAI21_X1 U_afifo_U_acore_U71 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n205), .A(U_afifo_U_acore_n204), .ZN(
        U_afifo_U_acore_n150) );
  OAI21_X1 U_afifo_U_acore_U70 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n201), .A(U_afifo_U_acore_n200), .ZN(
        U_afifo_U_acore_n148) );
  OAI21_X1 U_afifo_U_acore_U69 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n30), .A(U_afifo_U_acore_n188), .ZN(
        U_afifo_U_acore_n115) );
  OAI21_X1 U_afifo_U_acore_U68 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n175), .A(U_afifo_U_acore_n174), .ZN(
        U_afifo_U_acore_n107) );
  OAI21_X1 U_afifo_U_acore_U67 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n29), .A(U_afifo_U_acore_n187), .ZN(
        U_afifo_U_acore_n114) );
  OAI21_X1 U_afifo_U_acore_U66 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n28), .A(U_afifo_U_acore_n182), .ZN(
        U_afifo_U_acore_n111) );
  OAI21_X1 U_afifo_U_acore_U65 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n197), .A(U_afifo_U_acore_n196), .ZN(
        U_afifo_U_acore_n146) );
  OAI21_X1 U_afifo_U_acore_U64 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n177), .A(U_afifo_U_acore_n176), .ZN(
        U_afifo_U_acore_n108) );
  OAI21_X1 U_afifo_U_acore_U63 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n33), .A(U_afifo_U_acore_n195), .ZN(
        U_afifo_U_acore_n121) );
  OAI21_X1 U_afifo_U_acore_U62 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n184), .A(U_afifo_U_acore_n183), .ZN(
        U_afifo_U_acore_n112) );
  OAI21_X1 U_afifo_U_acore_U61 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n194), .A(U_afifo_U_acore_n193), .ZN(
        U_afifo_U_acore_n118) );
  OAI21_X1 U_afifo_U_acore_U60 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n70), .A(U_afifo_U_acore_n69), .ZN(
        U_afifo_U_acore_n120) );
  OAI21_X1 U_afifo_U_acore_U59 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n186), .A(U_afifo_U_acore_n185), .ZN(
        U_afifo_U_acore_n113) );
  OAI21_X1 U_afifo_U_acore_U58 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n173), .A(U_afifo_U_acore_n172), .ZN(
        U_afifo_U_acore_n106) );
  OAI21_X1 U_afifo_U_acore_U57 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n32), .A(U_afifo_U_acore_n171), .ZN(
        U_afifo_U_acore_n105) );
  OAI21_X1 U_afifo_U_acore_U56 ( .B1(U_afifo_U_acore_n68), .B2(
        U_afifo_U_acore_n41), .A(U_afifo_U_acore_n67), .ZN(
        U_afifo_U_acore_n119) );
  OAI21_X1 U_afifo_U_acore_U55 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n92), .A(U_afifo_U_acore_n91), .ZN(
        U_afifo_U_acore_n132) );
  OAI21_X1 U_afifo_U_acore_U54 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n98), .A(U_afifo_U_acore_n97), .ZN(
        U_afifo_U_acore_n135) );
  OAI21_X1 U_afifo_U_acore_U53 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n96), .A(U_afifo_U_acore_n95), .ZN(
        U_afifo_U_acore_n134) );
  OAI21_X1 U_afifo_U_acore_U52 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n100), .A(U_afifo_U_acore_n99), .ZN(
        U_afifo_U_acore_n136) );
  OAI21_X1 U_afifo_U_acore_U51 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n94), .A(U_afifo_U_acore_n93), .ZN(
        U_afifo_U_acore_n133) );
  OAI21_X1 U_afifo_U_acore_U50 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n102), .A(U_afifo_U_acore_n101), .ZN(
        U_afifo_U_acore_n137) );
  OAI21_X1 U_afifo_U_acore_U49 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n167), .A(U_afifo_U_acore_n164), .ZN(
        U_afifo_U_acore_n145) );
  OAI21_X1 U_afifo_U_acore_U48 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n104), .A(U_afifo_U_acore_n103), .ZN(
        U_afifo_U_acore_n138) );
  OAI21_X1 U_afifo_U_acore_U47 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n162), .A(U_afifo_U_acore_n161), .ZN(
        U_afifo_U_acore_n144) );
  OAI21_X1 U_afifo_U_acore_U46 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n160), .A(U_afifo_U_acore_n159), .ZN(
        U_afifo_U_acore_n142) );
  OAI21_X1 U_afifo_U_acore_U45 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n153), .A(U_afifo_U_acore_n143), .ZN(
        U_afifo_U_acore_n139) );
  OAI21_X1 U_afifo_U_acore_U44 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n158), .A(U_afifo_U_acore_n157), .ZN(
        U_afifo_U_acore_n141) );
  OAI21_X1 U_afifo_U_acore_U43 ( .B1(U_afifo_U_acore_n211), .B2(
        U_afifo_U_acore_n156), .A(U_afifo_U_acore_n155), .ZN(
        U_afifo_U_acore_n140) );
  OAI21_X1 U_afifo_U_acore_U42 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n90), .A(U_afifo_U_acore_n89), .ZN(
        U_afifo_U_acore_n131) );
  OAI21_X1 U_afifo_U_acore_U41 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n88), .A(U_afifo_U_acore_n87), .ZN(
        U_afifo_U_acore_n130) );
  OAI21_X1 U_afifo_U_acore_U40 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n82), .A(U_afifo_U_acore_n81), .ZN(
        U_afifo_U_acore_n127) );
  OAI21_X1 U_afifo_U_acore_U39 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n86), .A(U_afifo_U_acore_n85), .ZN(
        U_afifo_U_acore_n129) );
  OAI21_X1 U_afifo_U_acore_U38 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n80), .A(U_afifo_U_acore_n79), .ZN(
        U_afifo_U_acore_n126) );
  OAI21_X1 U_afifo_U_acore_U37 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n84), .A(U_afifo_U_acore_n83), .ZN(
        U_afifo_U_acore_n128) );
  NAND2_X1 U_afifo_U_acore_U36 ( .A1(U_afifo_U_acore_n35), .A2(
        U_afifo_U_acore_f_obuf_29_), .ZN(U_afifo_U_acore_n63) );
  INV_X2 U_afifo_U_acore_U35 ( .A(U_afifo_m_aempty), .ZN(U_afifo_U_acore_n47)
         );
  AOI22_X1 U_afifo_U_acore_U34 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_31_), .B1(U_afifo_U_acore_m_sf_data_out[31]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n87) );
  AOI22_X1 U_afifo_U_acore_U33 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_32_), .B1(U_afifo_U_acore_m_sf_data_out[32]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n85) );
  AOI22_X1 U_afifo_U_acore_U32 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_33_), .B1(U_afifo_U_acore_m_sf_data_out[33]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n83) );
  AOI22_X1 U_afifo_U_acore_U31 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_34_), .B1(U_afifo_U_acore_m_sf_data_out[34]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n81) );
  AOI22_X1 U_afifo_U_acore_U30 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_35_), .B1(U_afifo_U_acore_m_sf_data_out[35]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n79) );
  AOI22_X1 U_afifo_U_acore_U29 ( .A1(U_afifo_U_acore_n40), .A2(
        U_afifo_U_acore_f_obuf_30_), .B1(U_afifo_U_acore_m_sf_data_out[30]), 
        .B2(U_afifo_U_acore_n163), .ZN(U_afifo_U_acore_n89) );
  OAI21_X2 U_afifo_U_acore_U28 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n78), .A(U_afifo_U_acore_n77), .ZN(
        U_afifo_U_acore_n125) );
  OAI21_X2 U_afifo_U_acore_U27 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n74), .A(U_afifo_U_acore_n73), .ZN(
        U_afifo_U_acore_n123) );
  OAI21_X2 U_afifo_U_acore_U26 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n76), .A(U_afifo_U_acore_n75), .ZN(
        U_afifo_U_acore_n124) );
  OAI21_X2 U_afifo_U_acore_U25 ( .B1(U_afifo_U_acore_n41), .B2(
        U_afifo_U_acore_n72), .A(U_afifo_U_acore_n71), .ZN(
        U_afifo_U_acore_n122) );
  OAI22_X1 U_afifo_U_acore_U24 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n19), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n197), .ZN(hiu_addr[7]) );
  OAI22_X1 U_afifo_U_acore_U23 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n15), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n207), .ZN(hiu_addr[2]) );
  OAI22_X1 U_afifo_U_acore_U22 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n21), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n30), .ZN(hiu_haddr[0]) );
  OAI22_X1 U_afifo_U_acore_U21 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n18), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n199), .ZN(hiu_addr[6]) );
  OAI22_X1 U_afifo_U_acore_U20 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n22), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n29), .ZN(hiu_haddr[1]) );
  OAI22_X1 U_afifo_U_acore_U19 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n17), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n201), .ZN(hiu_addr[5]) );
  OAI22_X1 U_afifo_U_acore_U18 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n14), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n31), .ZN(hiu_addr[1]) );
  OAI22_X1 U_afifo_U_acore_U17 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n10), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n28), .ZN(U_afifo_m_data_out_49) );
  OAI22_X1 U_afifo_U_acore_U16 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n26), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n192), .ZN(hiu_hsize[1]) );
  OAI22_X1 U_afifo_U_acore_U15 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n27), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n190), .ZN(hiu_hsize[2]) );
  OAI22_X1 U_afifo_U_acore_U14 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n25), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n33), .ZN(U_afifo_m_data_out_3) );
  OAI22_X1 U_afifo_U_acore_U13 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n3), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n210), .ZN(U_afifo_m_data_out_0_) );
  OAI22_X1 U_afifo_U_acore_U12 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n20), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n194), .ZN(hiu_hsize[0]) );
  OAI22_X1 U_afifo_U_acore_U11 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n9), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n203), .ZN(hiu_addr[4]) );
  OAI22_X1 U_afifo_U_acore_U10 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n16), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n205), .ZN(hiu_addr[3]) );
  OAI22_X2 U_afifo_U_acore_U9 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n5), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n179), .ZN(hiu_burst_size[1]) );
  OAI22_X1 U_afifo_U_acore_U8 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n6), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n177), .ZN(hiu_burst_size[2]) );
  OAI22_X1 U_afifo_U_acore_U7 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n23), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n186), .ZN(hiu_haddr[2]) );
  OAI22_X1 U_afifo_U_acore_U6 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n13), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n173), .ZN(hiu_burst_size[4]) );
  OAI22_X1 U_afifo_U_acore_U5 ( .A1(U_afifo_U_acore_n1), .A2(
        U_afifo_U_acore_n24), .B1(U_afifo_U_acore_n35), .B2(
        U_afifo_U_acore_n184), .ZN(hiu_haddr[3]) );
  OAI21_X2 U_afifo_U_acore_U4 ( .B1(U_afifo_U_acore_n104), .B2(
        U_afifo_U_acore_n37), .A(U_afifo_U_acore_n58), .ZN(hiu_addr[14]) );
  OAI21_X2 U_afifo_U_acore_U3 ( .B1(U_afifo_U_acore_n158), .B2(
        U_afifo_U_acore_n37), .A(U_afifo_U_acore_n55), .ZN(hiu_addr[11]) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_5_ ( .D(U_afifo_m_data_in[5]), .CK(hclk), 
        .RN(hresetn), .QN(U_afifo_U_acore_n179) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_6_ ( .D(U_afifo_m_data_in[6]), .CK(hclk), 
        .RN(hresetn), .QN(U_afifo_U_acore_n177) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_7_ ( .D(U_afifo_m_data_in[7]), .CK(hclk), 
        .RN(hresetn), .QN(U_afifo_U_acore_n175) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_8_ ( .D(U_afifo_m_data_in[8]), .CK(hclk), 
        .RN(hresetn), .QN(U_afifo_U_acore_n173) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_44_ ( .D(U_afifo_m_data_in[44]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n190) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_0_ ( .D(U_afifo_m_data_in[0]), .CK(hclk), 
        .RN(hresetn), .QN(U_afifo_U_acore_n210) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_43_ ( .D(U_afifo_m_data_in[43]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n192) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_18_ ( .D(U_afifo_m_data_in[18]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_18_), .QN(U_afifo_U_acore_n167) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_15_ ( .D(U_afifo_m_data_in[15]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n201) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_14_ ( .D(U_afifo_m_data_in[14]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n203) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_47_ ( .D(U_afifo_m_data_in[47]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n186) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_48_ ( .D(U_afifo_m_data_in[48]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n184) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_2_ ( .D(U_afifo_m_data_in[2]), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_2_), .QN(U_afifo_U_acore_n92)
         );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_19_ ( .D(U_afifo_m_data_in[19]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n162) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_20_ ( .D(U_afifo_m_data_in[20]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n160) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_21_ ( .D(U_afifo_m_data_in[21]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n158) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_22_ ( .D(U_afifo_m_data_in[22]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n156) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_23_ ( .D(U_afifo_m_data_in[23]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n153) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_24_ ( .D(U_afifo_m_data_in[24]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n104) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_25_ ( .D(U_afifo_m_data_in[25]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n102) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_26_ ( .D(U_afifo_m_data_in[26]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n100) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_27_ ( .D(U_afifo_m_data_in[27]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n98) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_28_ ( .D(U_afifo_m_data_in[28]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n96) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_29_ ( .D(U_afifo_m_data_in[29]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n94) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_30_ ( .D(U_afifo_m_data_in[30]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_30_), .QN(U_afifo_U_acore_n90) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_31_ ( .D(U_afifo_m_data_in[31]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_31_), .QN(U_afifo_U_acore_n88) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_32_ ( .D(U_afifo_m_data_in[32]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_32_), .QN(U_afifo_U_acore_n86) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_33_ ( .D(U_afifo_m_data_in[33]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_33_), .QN(U_afifo_U_acore_n84) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_34_ ( .D(U_afifo_m_data_in[34]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_34_), .QN(U_afifo_U_acore_n82) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_35_ ( .D(U_afifo_m_data_in[35]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_35_), .QN(U_afifo_U_acore_n80) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_36_ ( .D(U_afifo_m_data_in[36]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_36_), .QN(U_afifo_U_acore_n78) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_37_ ( .D(U_afifo_m_data_in[37]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_37_), .QN(U_afifo_U_acore_n76) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_38_ ( .D(U_afifo_m_data_in[38]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_38_), .QN(U_afifo_U_acore_n74) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_39_ ( .D(U_afifo_m_data_in[39]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_39_), .QN(U_afifo_U_acore_n72) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_40_ ( .D(U_afifo_m_data_in[40]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_40_), .QN(U_afifo_U_acore_n70) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_41_ ( .D(U_afifo_m_data_in[41]), .CK(hclk), .RN(hresetn), .Q(U_afifo_U_acore_f_ibuf_41_), .QN(U_afifo_U_acore_n68) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_42_ ( .D(U_afifo_m_data_in[42]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n194) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_17_ ( .D(U_afifo_m_data_in[17]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n197) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_13_ ( .D(U_afifo_m_data_in[13]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n205) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_16_ ( .D(U_afifo_m_data_in[16]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n199) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_12_ ( .D(U_afifo_m_data_in[12]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n207) );
  DFFR_X2 U_afifo_U_acore_f_ibuf_reg_4_ ( .D(U_afifo_m_data_in[4]), .CK(hclk), 
        .RN(hresetn), .QN(U_afifo_U_acore_n181) );
  DFFR_X1 U_afifo_U_acore_f_afull_reg ( .D(U_afifo_U_acore_n_afull), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_afull), .QN(U_afifo_U_acore_n12) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_9_ ( .D(U_afifo_U_acore_n105), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_9_), .QN(U_afifo_U_acore_n8)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_8_ ( .D(U_afifo_U_acore_n106), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_8_), .QN(U_afifo_U_acore_n13)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_7_ ( .D(U_afifo_U_acore_n107), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_7_), .QN(U_afifo_U_acore_n7)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_6_ ( .D(U_afifo_U_acore_n108), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_6_), .QN(U_afifo_U_acore_n6)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_5_ ( .D(U_afifo_U_acore_n109), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_5_), .QN(U_afifo_U_acore_n5)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_4_ ( .D(U_afifo_U_acore_n110), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_4_), .QN(U_afifo_U_acore_n4)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_49_ ( .D(U_afifo_U_acore_n111), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_49_), .QN(U_afifo_U_acore_n10)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_48_ ( .D(U_afifo_U_acore_n112), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_48_), .QN(U_afifo_U_acore_n24)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_47_ ( .D(U_afifo_U_acore_n113), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_47_), .QN(U_afifo_U_acore_n23)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_46_ ( .D(U_afifo_U_acore_n114), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_46_), .QN(U_afifo_U_acore_n22)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_45_ ( .D(U_afifo_U_acore_n115), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_45_), .QN(U_afifo_U_acore_n21)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_44_ ( .D(U_afifo_U_acore_n116), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_44_), .QN(U_afifo_U_acore_n27)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_43_ ( .D(U_afifo_U_acore_n117), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_43_), .QN(U_afifo_U_acore_n26)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_42_ ( .D(U_afifo_U_acore_n118), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_42_), .QN(U_afifo_U_acore_n20)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_41_ ( .D(U_afifo_U_acore_n119), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_41_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_40_ ( .D(U_afifo_U_acore_n120), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_40_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_3_ ( .D(U_afifo_U_acore_n121), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_3_), .QN(U_afifo_U_acore_n25)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_39_ ( .D(U_afifo_U_acore_n122), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_39_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_38_ ( .D(U_afifo_U_acore_n123), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_38_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_37_ ( .D(U_afifo_U_acore_n124), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_37_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_36_ ( .D(U_afifo_U_acore_n125), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_36_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_35_ ( .D(U_afifo_U_acore_n126), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_35_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_34_ ( .D(U_afifo_U_acore_n127), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_34_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_33_ ( .D(U_afifo_U_acore_n128), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_33_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_32_ ( .D(U_afifo_U_acore_n129), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_32_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_31_ ( .D(U_afifo_U_acore_n130), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_31_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_30_ ( .D(U_afifo_U_acore_n131), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_30_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_2_ ( .D(U_afifo_U_acore_n132), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_2_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_29_ ( .D(U_afifo_U_acore_n133), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_29_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_28_ ( .D(U_afifo_U_acore_n134), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_28_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_27_ ( .D(U_afifo_U_acore_n135), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_27_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_26_ ( .D(U_afifo_U_acore_n136), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_26_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_25_ ( .D(U_afifo_U_acore_n137), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_25_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_24_ ( .D(U_afifo_U_acore_n138), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_24_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_23_ ( .D(U_afifo_U_acore_n139), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_23_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_22_ ( .D(U_afifo_U_acore_n140), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_22_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_21_ ( .D(U_afifo_U_acore_n141), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_21_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_20_ ( .D(U_afifo_U_acore_n142), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_20_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_19_ ( .D(U_afifo_U_acore_n144), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_19_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_18_ ( .D(U_afifo_U_acore_n145), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_18_) );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_17_ ( .D(U_afifo_U_acore_n146), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_17_), .QN(U_afifo_U_acore_n19)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_16_ ( .D(U_afifo_U_acore_n147), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_16_), .QN(U_afifo_U_acore_n18)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_15_ ( .D(U_afifo_U_acore_n148), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_15_), .QN(U_afifo_U_acore_n17)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_14_ ( .D(U_afifo_U_acore_n149), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_14_), .QN(U_afifo_U_acore_n9)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_13_ ( .D(U_afifo_U_acore_n150), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_13_), .QN(U_afifo_U_acore_n16)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_12_ ( .D(U_afifo_U_acore_n151), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_12_), .QN(U_afifo_U_acore_n15)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_11_ ( .D(U_afifo_U_acore_n152), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_11_), .QN(U_afifo_U_acore_n14)
         );
  DFFR_X1 U_afifo_U_acore_f_obuf_reg_0_ ( .D(U_afifo_U_acore_n154), .CK(hclk), 
        .RN(hresetn), .Q(U_afifo_U_acore_f_obuf_0_), .QN(U_afifo_U_acore_n3)
         );
  DFFS_X2 U_afifo_U_acore_f_obuf_empty_reg ( .D(U_afifo_U_acore_n_obuf_empty), 
        .CK(hclk), .SN(hresetn), .Q(U_afifo_U_acore_n34), .QN(
        U_afifo_U_acore_n38) );
  DFFS_X2 U_afifo_U_acore_f_push_req_n_reg ( .D(U_afifo_n55), .CK(hclk), .SN(
        hresetn), .Q(U_afifo_U_acore_f_push_req_n), .QN(U_afifo_U_acore_n11)
         );
  DFFR_X1 U_afifo_U_acore_f_ibuf_reg_3_ ( .D(U_afifo_m_data_in[3]), .CK(hclk), 
        .RN(hresetn), .QN(U_afifo_U_acore_n33) );
  DFFR_X1 U_afifo_U_acore_f_ibuf_reg_9_ ( .D(U_afifo_m_data_in[9]), .CK(hclk), 
        .RN(hresetn), .QN(U_afifo_U_acore_n32) );
  DFFR_X1 U_afifo_U_acore_f_ibuf_reg_11_ ( .D(U_afifo_m_data_in[11]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n31) );
  DFFR_X1 U_afifo_U_acore_f_ibuf_reg_45_ ( .D(U_afifo_m_data_in[45]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n30) );
  DFFR_X1 U_afifo_U_acore_f_ibuf_reg_46_ ( .D(U_afifo_m_data_in[46]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n29) );
  DFFR_X1 U_afifo_U_acore_f_ibuf_reg_49_ ( .D(U_afifo_m_data_in[49]), .CK(hclk), .RN(hresetn), .QN(U_afifo_U_acore_n28) );
  AOI22_X1 U_dfifo_U_dcore_U224 ( .A1(U_dfifo_U_dcore_f_buf_data_0_), .A2(
        U_dfifo_U_dcore_n126), .B1(U_dfifo_m_data_out_0_), .B2(
        U_dfifo_U_dcore_n125), .ZN(U_dfifo_U_dcore_n129) );
  AOI22_X1 U_dfifo_U_dcore_U223 ( .A1(U_dfifo_U_dcore_f_buf_data_1_), .A2(
        U_dfifo_U_dcore_n126), .B1(U_dfifo_m_data_out_1_), .B2(
        U_dfifo_U_dcore_n125), .ZN(U_dfifo_U_dcore_n124) );
  AOI22_X1 U_dfifo_U_dcore_U222 ( .A1(U_dfifo_U_dcore_f_buf_data_33_), .A2(
        U_dfifo_U_dcore_n126), .B1(hiu_data[31]), .B2(U_dfifo_U_dcore_n125), 
        .ZN(U_dfifo_U_dcore_n122) );
  AOI22_X1 U_dfifo_U_dcore_U221 ( .A1(U_dfifo_U_dcore_f_buf_data_32_), .A2(
        U_dfifo_U_dcore_n126), .B1(hiu_data[30]), .B2(U_dfifo_U_dcore_n125), 
        .ZN(U_dfifo_U_dcore_n120) );
  AOI22_X1 U_dfifo_U_dcore_U220 ( .A1(U_dfifo_U_dcore_f_buf_data_31_), .A2(
        U_dfifo_U_dcore_n126), .B1(hiu_data[29]), .B2(U_dfifo_U_dcore_n125), 
        .ZN(U_dfifo_U_dcore_n118) );
  AOI22_X1 U_dfifo_U_dcore_U219 ( .A1(U_dfifo_U_dcore_f_buf_data_30_), .A2(
        U_dfifo_U_dcore_n126), .B1(hiu_data[28]), .B2(U_dfifo_U_dcore_n125), 
        .ZN(U_dfifo_U_dcore_n116) );
  AOI22_X1 U_dfifo_U_dcore_U218 ( .A1(U_dfifo_U_dcore_f_buf_data_29_), .A2(
        U_dfifo_U_dcore_n126), .B1(hiu_data[27]), .B2(U_dfifo_U_dcore_n125), 
        .ZN(U_dfifo_U_dcore_n114) );
  AOI22_X1 U_dfifo_U_dcore_U217 ( .A1(U_dfifo_U_dcore_f_buf_data_28_), .A2(
        U_dfifo_U_dcore_n126), .B1(hiu_data[26]), .B2(U_dfifo_U_dcore_n125), 
        .ZN(U_dfifo_U_dcore_n112) );
  AOI22_X1 U_dfifo_U_dcore_U216 ( .A1(U_dfifo_U_dcore_f_buf_data_27_), .A2(
        U_dfifo_U_dcore_n126), .B1(hiu_data[25]), .B2(U_dfifo_U_dcore_n125), 
        .ZN(U_dfifo_U_dcore_n110) );
  AOI22_X1 U_dfifo_U_dcore_U215 ( .A1(U_dfifo_U_dcore_f_buf_data_26_), .A2(
        U_dfifo_U_dcore_n126), .B1(hiu_data[24]), .B2(U_dfifo_U_dcore_n125), 
        .ZN(U_dfifo_U_dcore_n108) );
  NAND2_X2 U_dfifo_U_dcore_U213 ( .A1(U_dfifo_U_dcore_n28), .A2(
        U_dfifo_U_dcore_n125), .ZN(U_dfifo_U_dcore_n106) );
  NOR2_X4 U_dfifo_U_dcore_U212 ( .A1(U_dfifo_m_empty), .A2(
        U_dfifo_U_dcore_n209), .ZN(U_dfifo_U_dcore_n127) );
  AND2_X4 U_dfifo_U_dcore_U211 ( .A1(m_df_push_n), .A2(U_dfifo_U_dcore_n27), 
        .ZN(U_dfifo_U_dcore_n2) );
  NOR4_X4 U_dfifo_U_dcore_U210 ( .A1(U_dfifo_m_empty), .A2(U_dfifo_m_aempty), 
        .A3(U_dfifo_U_dcore_n26), .A4(U_dfifo_U_dcore_n25), .ZN(
        U_dfifo_U_dcore_n126) );
  INV_X4 U_dfifo_U_dcore_U209 ( .A(U_dfifo_U_dcore_m_sf_empty), .ZN(
        U_dfifo_U_dcore_n25) );
  NOR2_X2 U_dfifo_U_dcore_U208 ( .A1(U_dfifo_U_dcore_f_buf_has_data), .A2(
        U_dfifo_U_dcore_n25), .ZN(U_dfifo_m_aempty) );
  AOI21_X2 U_dfifo_U_dcore_U207 ( .B1(U_dfifo_m_empty), .B2(m_df_push_n), .A(
        U_dfifo_n5), .ZN(U_dfifo_U_dcore_n125) );
  NAND2_X1 U_dfifo_U_dcore_U206 ( .A1(U_dfifo_m_empty), .A2(m_two_to_one), 
        .ZN(U_dfifo_U_dcore_n55) );
  NAND2_X2 U_dfifo_U_dcore_U205 ( .A1(U_dfifo_U_dcore_n125), .A2(
        U_dfifo_U_dcore_n55), .ZN(U_dfifo_U_dcore_n88) );
  AOI21_X2 U_dfifo_U_dcore_U204 ( .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[25]), .A(U_dfifo_U_dcore_n57), .ZN(
        U_dfifo_U_dcore_n59) );
  AOI21_X2 U_dfifo_U_dcore_U203 ( .B1(U_dfifo_n5), .B2(U_dfifo_m_aempty), .A(
        U_dfifo_m_empty), .ZN(U_dfifo_U_dcore_n27) );
  NOR2_X4 U_dfifo_U_dcore_U202 ( .A1(U_dfifo_U_dcore_n125), .A2(
        U_dfifo_U_dcore_n27), .ZN(U_dfifo_U_dcore_n3) );
  OAI211_X2 U_dfifo_U_dcore_U201 ( .C1(U_dfifo_U_dcore_n14), .C2(
        U_dfifo_U_dcore_n88), .A(U_dfifo_U_dcore_n59), .B(U_dfifo_U_dcore_n58), 
        .ZN(U_dfifo_U_dcore_n142) );
  AOI21_X2 U_dfifo_U_dcore_U200 ( .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[18]), .A(U_dfifo_U_dcore_n85), .ZN(
        U_dfifo_U_dcore_n87) );
  OAI211_X2 U_dfifo_U_dcore_U199 ( .C1(U_dfifo_U_dcore_n13), .C2(
        U_dfifo_U_dcore_n88), .A(U_dfifo_U_dcore_n87), .B(U_dfifo_U_dcore_n86), 
        .ZN(U_dfifo_U_dcore_n149) );
  NOR2_X2 U_dfifo_U_dcore_U198 ( .A1(U_dfifo_m_empty), .A2(U_dfifo_n5), .ZN(
        U_dfifo_U_dcore_n103) );
  OAI211_X2 U_dfifo_U_dcore_U197 ( .C1(U_dfifo_U_dcore_n106), .C2(
        U_dfifo_U_dcore_n5), .A(U_dfifo_U_dcore_n90), .B(U_dfifo_U_dcore_n89), 
        .ZN(U_dfifo_U_dcore_n150) );
  OAI211_X2 U_dfifo_U_dcore_U196 ( .C1(U_dfifo_U_dcore_n106), .C2(
        U_dfifo_U_dcore_n11), .A(U_dfifo_U_dcore_n105), .B(
        U_dfifo_U_dcore_n104), .ZN(U_dfifo_U_dcore_n157) );
  NAND2_X2 U_dfifo_U_dcore_U195 ( .A1(U_dfifo_U_dcore_m_sf_afull), .A2(
        U_dfifo_U_dcore_f_buf_has_data), .ZN(U_dfifo_U_dcore_n21) );
  AOI22_X2 U_dfifo_U_dcore_U194 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_9_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[9]), .ZN(U_dfifo_U_dcore_n53) );
  NAND4_X2 U_dfifo_U_dcore_U193 ( .A1(U_dfifo_U_dcore_n54), .A2(
        U_dfifo_U_dcore_n53), .A3(U_dfifo_U_dcore_n52), .A4(
        U_dfifo_U_dcore_n56), .ZN(U_dfifo_U_dcore_n141) );
  AOI22_X2 U_dfifo_U_dcore_U192 ( .A1(U_dfifo_U_dcore_f_buf_data_2_), .A2(
        U_dfifo_U_dcore_n126), .B1(m_df_data_in[2]), .B2(U_dfifo_U_dcore_n3), 
        .ZN(U_dfifo_U_dcore_n30) );
  NAND4_X2 U_dfifo_U_dcore_U191 ( .A1(U_dfifo_U_dcore_n31), .A2(
        U_dfifo_U_dcore_n30), .A3(U_dfifo_U_dcore_n29), .A4(
        U_dfifo_U_dcore_n84), .ZN(U_dfifo_U_dcore_n134) );
  AOI21_X2 U_dfifo_U_dcore_U190 ( .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[24]), .A(U_dfifo_U_dcore_n61), .ZN(
        U_dfifo_U_dcore_n63) );
  OAI211_X2 U_dfifo_U_dcore_U189 ( .C1(U_dfifo_U_dcore_n15), .C2(
        U_dfifo_U_dcore_n88), .A(U_dfifo_U_dcore_n63), .B(U_dfifo_U_dcore_n62), 
        .ZN(U_dfifo_U_dcore_n143) );
  OAI211_X2 U_dfifo_U_dcore_U188 ( .C1(U_dfifo_U_dcore_n106), .C2(
        U_dfifo_U_dcore_n8), .A(U_dfifo_U_dcore_n98), .B(U_dfifo_U_dcore_n97), 
        .ZN(U_dfifo_U_dcore_n154) );
  OAI211_X2 U_dfifo_U_dcore_U187 ( .C1(U_dfifo_U_dcore_n106), .C2(
        U_dfifo_U_dcore_n6), .A(U_dfifo_U_dcore_n92), .B(U_dfifo_U_dcore_n91), 
        .ZN(U_dfifo_U_dcore_n151) );
  OAI211_X2 U_dfifo_U_dcore_U186 ( .C1(U_dfifo_U_dcore_n106), .C2(
        U_dfifo_U_dcore_n7), .A(U_dfifo_U_dcore_n96), .B(U_dfifo_U_dcore_n95), 
        .ZN(U_dfifo_U_dcore_n153) );
  OAI211_X2 U_dfifo_U_dcore_U185 ( .C1(U_dfifo_U_dcore_n106), .C2(
        U_dfifo_U_dcore_n12), .A(U_dfifo_U_dcore_n94), .B(U_dfifo_U_dcore_n93), 
        .ZN(U_dfifo_U_dcore_n152) );
  AOI22_X2 U_dfifo_U_dcore_U184 ( .A1(U_dfifo_U_dcore_n3), .A2(
        m_df_data_in[33]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[33]), .ZN(U_dfifo_U_dcore_n121) );
  NAND2_X2 U_dfifo_U_dcore_U183 ( .A1(U_dfifo_U_dcore_n122), .A2(
        U_dfifo_U_dcore_n121), .ZN(U_dfifo_U_dcore_n165) );
  AOI22_X2 U_dfifo_U_dcore_U182 ( .A1(U_dfifo_U_dcore_n3), .A2(
        m_df_data_in[26]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[26]), .ZN(U_dfifo_U_dcore_n107) );
  NAND2_X2 U_dfifo_U_dcore_U181 ( .A1(U_dfifo_U_dcore_n108), .A2(
        U_dfifo_U_dcore_n107), .ZN(U_dfifo_U_dcore_n158) );
  AOI21_X2 U_dfifo_U_dcore_U180 ( .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[23]), .A(U_dfifo_U_dcore_n65), .ZN(
        U_dfifo_U_dcore_n67) );
  OAI211_X2 U_dfifo_U_dcore_U179 ( .C1(U_dfifo_U_dcore_n16), .C2(
        U_dfifo_U_dcore_n88), .A(U_dfifo_U_dcore_n67), .B(U_dfifo_U_dcore_n66), 
        .ZN(U_dfifo_U_dcore_n144) );
  OAI211_X2 U_dfifo_U_dcore_U178 ( .C1(U_dfifo_U_dcore_n106), .C2(
        U_dfifo_U_dcore_n10), .A(U_dfifo_U_dcore_n102), .B(
        U_dfifo_U_dcore_n101), .ZN(U_dfifo_U_dcore_n156) );
  OAI211_X2 U_dfifo_U_dcore_U177 ( .C1(U_dfifo_U_dcore_n106), .C2(
        U_dfifo_U_dcore_n9), .A(U_dfifo_U_dcore_n100), .B(U_dfifo_U_dcore_n99), 
        .ZN(U_dfifo_U_dcore_n155) );
  OAI22_X2 U_dfifo_U_dcore_U176 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[33]), .B1(U_dfifo_U_dcore_f_buf_data_33_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n234) );
  INV_X4 U_dfifo_U_dcore_U175 ( .A(U_dfifo_U_dcore_n234), .ZN(
        U_dfifo_U_dcore_n201) );
  OAI22_X2 U_dfifo_U_dcore_U174 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[26]), .B1(U_dfifo_U_dcore_f_buf_data_26_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n227) );
  INV_X4 U_dfifo_U_dcore_U173 ( .A(U_dfifo_U_dcore_n227), .ZN(
        U_dfifo_U_dcore_n194) );
  OAI22_X2 U_dfifo_U_dcore_U172 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[18]), .B1(U_dfifo_U_dcore_f_buf_data_18_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n219) );
  INV_X4 U_dfifo_U_dcore_U171 ( .A(U_dfifo_U_dcore_n219), .ZN(
        U_dfifo_U_dcore_n186) );
  OAI22_X2 U_dfifo_U_dcore_U170 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[25]), .B1(U_dfifo_U_dcore_f_buf_data_25_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n226) );
  INV_X4 U_dfifo_U_dcore_U169 ( .A(U_dfifo_U_dcore_n226), .ZN(
        U_dfifo_U_dcore_n193) );
  AOI21_X2 U_dfifo_U_dcore_U168 ( .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[20]), .A(U_dfifo_U_dcore_n77), .ZN(
        U_dfifo_U_dcore_n79) );
  OAI211_X2 U_dfifo_U_dcore_U167 ( .C1(U_dfifo_U_dcore_n19), .C2(
        U_dfifo_U_dcore_n88), .A(U_dfifo_U_dcore_n79), .B(U_dfifo_U_dcore_n78), 
        .ZN(U_dfifo_U_dcore_n147) );
  AOI21_X2 U_dfifo_U_dcore_U166 ( .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[19]), .A(U_dfifo_U_dcore_n81), .ZN(
        U_dfifo_U_dcore_n83) );
  OAI211_X2 U_dfifo_U_dcore_U165 ( .C1(U_dfifo_U_dcore_n20), .C2(
        U_dfifo_U_dcore_n88), .A(U_dfifo_U_dcore_n83), .B(U_dfifo_U_dcore_n82), 
        .ZN(U_dfifo_U_dcore_n148) );
  AOI21_X2 U_dfifo_U_dcore_U164 ( .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[22]), .A(U_dfifo_U_dcore_n69), .ZN(
        U_dfifo_U_dcore_n71) );
  OAI211_X2 U_dfifo_U_dcore_U163 ( .C1(U_dfifo_U_dcore_n17), .C2(
        U_dfifo_U_dcore_n88), .A(U_dfifo_U_dcore_n71), .B(U_dfifo_U_dcore_n70), 
        .ZN(U_dfifo_U_dcore_n145) );
  AOI21_X2 U_dfifo_U_dcore_U162 ( .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[21]), .A(U_dfifo_U_dcore_n73), .ZN(
        U_dfifo_U_dcore_n75) );
  OAI211_X2 U_dfifo_U_dcore_U161 ( .C1(U_dfifo_U_dcore_n18), .C2(
        U_dfifo_U_dcore_n88), .A(U_dfifo_U_dcore_n75), .B(U_dfifo_U_dcore_n74), 
        .ZN(U_dfifo_U_dcore_n146) );
  NAND4_X2 U_dfifo_U_dcore_U160 ( .A1(U_dfifo_U_dcore_n49), .A2(
        U_dfifo_U_dcore_n48), .A3(U_dfifo_U_dcore_n47), .A4(
        U_dfifo_U_dcore_n60), .ZN(U_dfifo_U_dcore_n140) );
  OAI221_X2 U_dfifo_U_dcore_U159 ( .B1(U_dfifo_n5), .B2(U_dfifo_U_dcore_n24), 
        .C1(U_dfifo_U_dcore_n26), .C2(U_dfifo_U_dcore_n25), .A(
        U_dfifo_U_dcore_f_buf_has_data), .ZN(U_dfifo_U_dcore_n208) );
  NAND4_X2 U_dfifo_U_dcore_U158 ( .A1(U_dfifo_U_dcore_n40), .A2(
        U_dfifo_U_dcore_n39), .A3(U_dfifo_U_dcore_n38), .A4(
        U_dfifo_U_dcore_n72), .ZN(U_dfifo_U_dcore_n137) );
  NAND4_X2 U_dfifo_U_dcore_U157 ( .A1(U_dfifo_U_dcore_n37), .A2(
        U_dfifo_U_dcore_n36), .A3(U_dfifo_U_dcore_n35), .A4(
        U_dfifo_U_dcore_n76), .ZN(U_dfifo_U_dcore_n136) );
  NAND4_X2 U_dfifo_U_dcore_U156 ( .A1(U_dfifo_U_dcore_n46), .A2(
        U_dfifo_U_dcore_n45), .A3(U_dfifo_U_dcore_n44), .A4(
        U_dfifo_U_dcore_n64), .ZN(U_dfifo_U_dcore_n139) );
  NAND4_X2 U_dfifo_U_dcore_U155 ( .A1(U_dfifo_U_dcore_n43), .A2(
        U_dfifo_U_dcore_n42), .A3(U_dfifo_U_dcore_n41), .A4(
        U_dfifo_U_dcore_n68), .ZN(U_dfifo_U_dcore_n138) );
  NAND4_X2 U_dfifo_U_dcore_U154 ( .A1(U_dfifo_U_dcore_n34), .A2(
        U_dfifo_U_dcore_n33), .A3(U_dfifo_U_dcore_n32), .A4(
        U_dfifo_U_dcore_n80), .ZN(U_dfifo_U_dcore_n135) );
  OAI22_X2 U_dfifo_U_dcore_U153 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[2]), .B1(U_dfifo_U_dcore_f_buf_data_2_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n132) );
  INV_X4 U_dfifo_U_dcore_U152 ( .A(U_dfifo_U_dcore_n132), .ZN(
        U_dfifo_U_dcore_n170) );
  OAI22_X2 U_dfifo_U_dcore_U151 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[17]), .B1(U_dfifo_U_dcore_f_buf_data_17_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n218) );
  INV_X4 U_dfifo_U_dcore_U150 ( .A(U_dfifo_U_dcore_n218), .ZN(
        U_dfifo_U_dcore_n185) );
  OAI22_X2 U_dfifo_U_dcore_U149 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[9]), .B1(U_dfifo_U_dcore_f_buf_data_9_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n210) );
  INV_X4 U_dfifo_U_dcore_U148 ( .A(U_dfifo_U_dcore_n210), .ZN(
        U_dfifo_U_dcore_n177) );
  OAI22_X2 U_dfifo_U_dcore_U147 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[10]), .B1(U_dfifo_U_dcore_f_buf_data_10_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n211) );
  INV_X4 U_dfifo_U_dcore_U146 ( .A(U_dfifo_U_dcore_n211), .ZN(
        U_dfifo_U_dcore_n178) );
  AOI22_X2 U_dfifo_U_dcore_U145 ( .A1(U_dfifo_U_dcore_n3), .A2(
        m_df_data_in[31]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[31]), .ZN(U_dfifo_U_dcore_n117) );
  NAND2_X2 U_dfifo_U_dcore_U144 ( .A1(U_dfifo_U_dcore_n118), .A2(
        U_dfifo_U_dcore_n117), .ZN(U_dfifo_U_dcore_n163) );
  AOI22_X2 U_dfifo_U_dcore_U143 ( .A1(U_dfifo_U_dcore_n3), .A2(
        m_df_data_in[32]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[32]), .ZN(U_dfifo_U_dcore_n119) );
  NAND2_X2 U_dfifo_U_dcore_U142 ( .A1(U_dfifo_U_dcore_n120), .A2(
        U_dfifo_U_dcore_n119), .ZN(U_dfifo_U_dcore_n164) );
  AOI22_X2 U_dfifo_U_dcore_U141 ( .A1(U_dfifo_U_dcore_n3), .A2(m_df_data_in[0]), .B1(U_dfifo_U_dcore_n127), .B2(U_dfifo_U_dcore_m_sf_data_out[0]), .ZN(
        U_dfifo_U_dcore_n128) );
  NAND2_X2 U_dfifo_U_dcore_U140 ( .A1(U_dfifo_U_dcore_n129), .A2(
        U_dfifo_U_dcore_n128), .ZN(U_dfifo_U_dcore_n167) );
  OAI22_X2 U_dfifo_U_dcore_U139 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[24]), .B1(U_dfifo_U_dcore_f_buf_data_24_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n225) );
  INV_X4 U_dfifo_U_dcore_U138 ( .A(U_dfifo_U_dcore_n225), .ZN(
        U_dfifo_U_dcore_n192) );
  OAI22_X2 U_dfifo_U_dcore_U137 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[31]), .B1(U_dfifo_U_dcore_f_buf_data_31_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n232) );
  INV_X4 U_dfifo_U_dcore_U136 ( .A(U_dfifo_U_dcore_n232), .ZN(
        U_dfifo_U_dcore_n199) );
  OAI22_X2 U_dfifo_U_dcore_U135 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[32]), .B1(U_dfifo_U_dcore_f_buf_data_32_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n233) );
  INV_X4 U_dfifo_U_dcore_U134 ( .A(U_dfifo_U_dcore_n233), .ZN(
        U_dfifo_U_dcore_n200) );
  AOI22_X2 U_dfifo_U_dcore_U133 ( .A1(U_dfifo_U_dcore_n3), .A2(
        m_df_data_in[28]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[28]), .ZN(U_dfifo_U_dcore_n111) );
  NAND2_X2 U_dfifo_U_dcore_U132 ( .A1(U_dfifo_U_dcore_n112), .A2(
        U_dfifo_U_dcore_n111), .ZN(U_dfifo_U_dcore_n160) );
  AOI22_X2 U_dfifo_U_dcore_U131 ( .A1(U_dfifo_U_dcore_n3), .A2(
        m_df_data_in[27]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[27]), .ZN(U_dfifo_U_dcore_n109) );
  NAND2_X2 U_dfifo_U_dcore_U130 ( .A1(U_dfifo_U_dcore_n110), .A2(
        U_dfifo_U_dcore_n109), .ZN(U_dfifo_U_dcore_n159) );
  AOI22_X2 U_dfifo_U_dcore_U129 ( .A1(U_dfifo_U_dcore_n3), .A2(
        m_df_data_in[29]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[29]), .ZN(U_dfifo_U_dcore_n113) );
  NAND2_X2 U_dfifo_U_dcore_U128 ( .A1(U_dfifo_U_dcore_n114), .A2(
        U_dfifo_U_dcore_n113), .ZN(U_dfifo_U_dcore_n161) );
  AOI22_X2 U_dfifo_U_dcore_U127 ( .A1(U_dfifo_U_dcore_n3), .A2(
        m_df_data_in[30]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[30]), .ZN(U_dfifo_U_dcore_n115) );
  NAND2_X2 U_dfifo_U_dcore_U126 ( .A1(U_dfifo_U_dcore_n116), .A2(
        U_dfifo_U_dcore_n115), .ZN(U_dfifo_U_dcore_n162) );
  OAI22_X2 U_dfifo_U_dcore_U125 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[15]), .B1(U_dfifo_U_dcore_f_buf_data_15_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n216) );
  INV_X4 U_dfifo_U_dcore_U124 ( .A(U_dfifo_U_dcore_n216), .ZN(
        U_dfifo_U_dcore_n183) );
  OAI22_X2 U_dfifo_U_dcore_U123 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[16]), .B1(U_dfifo_U_dcore_f_buf_data_16_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n217) );
  INV_X4 U_dfifo_U_dcore_U122 ( .A(U_dfifo_U_dcore_n217), .ZN(
        U_dfifo_U_dcore_n184) );
  OAI22_X2 U_dfifo_U_dcore_U121 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[8]), .B1(U_dfifo_U_dcore_f_buf_data_8_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n207) );
  INV_X4 U_dfifo_U_dcore_U120 ( .A(U_dfifo_U_dcore_n207), .ZN(
        U_dfifo_U_dcore_n176) );
  OAI22_X2 U_dfifo_U_dcore_U119 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[11]), .B1(U_dfifo_U_dcore_f_buf_data_11_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n212) );
  INV_X4 U_dfifo_U_dcore_U118 ( .A(U_dfifo_U_dcore_n212), .ZN(
        U_dfifo_U_dcore_n179) );
  OAI22_X2 U_dfifo_U_dcore_U117 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[13]), .B1(U_dfifo_U_dcore_f_buf_data_13_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n214) );
  INV_X4 U_dfifo_U_dcore_U116 ( .A(U_dfifo_U_dcore_n214), .ZN(
        U_dfifo_U_dcore_n181) );
  OAI22_X2 U_dfifo_U_dcore_U115 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[12]), .B1(U_dfifo_U_dcore_f_buf_data_12_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n213) );
  INV_X4 U_dfifo_U_dcore_U114 ( .A(U_dfifo_U_dcore_n213), .ZN(
        U_dfifo_U_dcore_n180) );
  OAI22_X2 U_dfifo_U_dcore_U113 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[14]), .B1(U_dfifo_U_dcore_f_buf_data_14_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n215) );
  INV_X4 U_dfifo_U_dcore_U112 ( .A(U_dfifo_U_dcore_n215), .ZN(
        U_dfifo_U_dcore_n182) );
  OAI22_X2 U_dfifo_U_dcore_U111 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[23]), .B1(U_dfifo_U_dcore_f_buf_data_23_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n224) );
  INV_X4 U_dfifo_U_dcore_U110 ( .A(U_dfifo_U_dcore_n224), .ZN(
        U_dfifo_U_dcore_n191) );
  OAI22_X2 U_dfifo_U_dcore_U109 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[19]), .B1(U_dfifo_U_dcore_f_buf_data_19_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n220) );
  INV_X4 U_dfifo_U_dcore_U108 ( .A(U_dfifo_U_dcore_n220), .ZN(
        U_dfifo_U_dcore_n187) );
  OAI22_X2 U_dfifo_U_dcore_U107 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[20]), .B1(U_dfifo_U_dcore_f_buf_data_20_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n221) );
  INV_X4 U_dfifo_U_dcore_U106 ( .A(U_dfifo_U_dcore_n221), .ZN(
        U_dfifo_U_dcore_n188) );
  OAI22_X2 U_dfifo_U_dcore_U105 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[21]), .B1(U_dfifo_U_dcore_f_buf_data_21_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n222) );
  INV_X4 U_dfifo_U_dcore_U104 ( .A(U_dfifo_U_dcore_n222), .ZN(
        U_dfifo_U_dcore_n189) );
  OAI22_X2 U_dfifo_U_dcore_U103 ( .A1(U_dfifo_U_dcore_n1), .A2(
        m_df_data_in[22]), .B1(U_dfifo_U_dcore_f_buf_data_22_), .B2(
        U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n223) );
  INV_X4 U_dfifo_U_dcore_U102 ( .A(U_dfifo_U_dcore_n223), .ZN(
        U_dfifo_U_dcore_n190) );
  OAI22_X2 U_dfifo_U_dcore_U101 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[0]), .B1(U_dfifo_U_dcore_f_buf_data_0_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n130) );
  INV_X4 U_dfifo_U_dcore_U100 ( .A(U_dfifo_U_dcore_n130), .ZN(
        U_dfifo_U_dcore_n168) );
  OAI22_X2 U_dfifo_U_dcore_U99 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[7]), 
        .B1(U_dfifo_U_dcore_f_buf_data_7_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n206) );
  INV_X4 U_dfifo_U_dcore_U98 ( .A(U_dfifo_U_dcore_n206), .ZN(
        U_dfifo_U_dcore_n175) );
  OAI22_X2 U_dfifo_U_dcore_U97 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[6]), 
        .B1(U_dfifo_U_dcore_f_buf_data_6_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n205) );
  INV_X4 U_dfifo_U_dcore_U96 ( .A(U_dfifo_U_dcore_n205), .ZN(
        U_dfifo_U_dcore_n174) );
  OAI22_X2 U_dfifo_U_dcore_U95 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[3]), 
        .B1(U_dfifo_U_dcore_f_buf_data_3_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n133) );
  INV_X4 U_dfifo_U_dcore_U94 ( .A(U_dfifo_U_dcore_n133), .ZN(
        U_dfifo_U_dcore_n171) );
  OAI22_X2 U_dfifo_U_dcore_U93 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[4]), 
        .B1(U_dfifo_U_dcore_f_buf_data_4_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n202) );
  INV_X4 U_dfifo_U_dcore_U92 ( .A(U_dfifo_U_dcore_n202), .ZN(
        U_dfifo_U_dcore_n172) );
  OAI22_X2 U_dfifo_U_dcore_U91 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[5]), 
        .B1(U_dfifo_U_dcore_f_buf_data_5_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n204) );
  INV_X4 U_dfifo_U_dcore_U90 ( .A(U_dfifo_U_dcore_n204), .ZN(
        U_dfifo_U_dcore_n173) );
  OAI22_X2 U_dfifo_U_dcore_U89 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[27]), .B1(U_dfifo_U_dcore_f_buf_data_27_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n228) );
  INV_X4 U_dfifo_U_dcore_U88 ( .A(U_dfifo_U_dcore_n228), .ZN(
        U_dfifo_U_dcore_n195) );
  OAI22_X2 U_dfifo_U_dcore_U87 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[29]), .B1(U_dfifo_U_dcore_f_buf_data_29_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n230) );
  INV_X4 U_dfifo_U_dcore_U86 ( .A(U_dfifo_U_dcore_n230), .ZN(
        U_dfifo_U_dcore_n197) );
  OAI22_X2 U_dfifo_U_dcore_U85 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[28]), .B1(U_dfifo_U_dcore_f_buf_data_28_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n229) );
  INV_X4 U_dfifo_U_dcore_U84 ( .A(U_dfifo_U_dcore_n229), .ZN(
        U_dfifo_U_dcore_n196) );
  OAI22_X2 U_dfifo_U_dcore_U83 ( .A1(U_dfifo_U_dcore_n1), .A2(m_df_data_in[30]), .B1(U_dfifo_U_dcore_f_buf_data_30_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n231) );
  INV_X4 U_dfifo_U_dcore_U82 ( .A(U_dfifo_U_dcore_n231), .ZN(
        U_dfifo_U_dcore_n198) );
  NAND2_X2 U_dfifo_U_dcore_U81 ( .A1(U_dfifo_U_dcore_n124), .A2(
        U_dfifo_U_dcore_n123), .ZN(U_dfifo_U_dcore_n166) );
  OAI22_X2 U_dfifo_U_dcore_U80 ( .A1(U_dfifo_U_dcore_n1), .A2(m_double), .B1(
        U_dfifo_U_dcore_f_buf_data_1_), .B2(U_dfifo_U_dcore_n2), .ZN(
        U_dfifo_U_dcore_n131) );
  INV_X4 U_dfifo_U_dcore_U79 ( .A(U_dfifo_U_dcore_n131), .ZN(
        U_dfifo_U_dcore_n169) );
  OAI21_X1 U_dfifo_U_dcore_U78 ( .B1(U_dfifo_n5), .B2(U_dfifo_U_dcore_n23), 
        .A(U_dfifo_U_dcore_n1), .ZN(U_dfifo_U_dcore_n203) );
  AOI22_X2 U_dfifo_U_dcore_U77 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_8_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[8]), .ZN(U_dfifo_U_dcore_n48) );
  AOI22_X2 U_dfifo_U_dcore_U76 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_5_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[5]), .ZN(U_dfifo_U_dcore_n39) );
  AOI22_X2 U_dfifo_U_dcore_U75 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_4_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[4]), .ZN(U_dfifo_U_dcore_n36) );
  AOI22_X2 U_dfifo_U_dcore_U74 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_7_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[7]), .ZN(U_dfifo_U_dcore_n45) );
  AOI22_X2 U_dfifo_U_dcore_U73 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_6_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[6]), .ZN(U_dfifo_U_dcore_n42) );
  AOI22_X2 U_dfifo_U_dcore_U72 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_3_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[3]), .ZN(U_dfifo_U_dcore_n33) );
  AOI22_X2 U_dfifo_U_dcore_U71 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_10_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[10]), .ZN(U_dfifo_U_dcore_n89) );
  AOI22_X2 U_dfifo_U_dcore_U70 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_17_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[17]), .ZN(U_dfifo_U_dcore_n104) );
  NOR3_X1 U_dfifo_U_dcore_U69 ( .A1(U_dfifo_n5), .A2(m_df_push_n), .A3(
        U_dfifo_U_dcore_n55), .ZN(U_dfifo_U_dcore_n51) );
  AOI22_X2 U_dfifo_U_dcore_U68 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_25_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[25]), .ZN(U_dfifo_U_dcore_n58) );
  AOI22_X2 U_dfifo_U_dcore_U67 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_18_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[18]), .ZN(U_dfifo_U_dcore_n86) );
  AOI22_X2 U_dfifo_U_dcore_U66 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_24_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[24]), .ZN(U_dfifo_U_dcore_n62) );
  AOI22_X2 U_dfifo_U_dcore_U65 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_14_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[14]), .ZN(U_dfifo_U_dcore_n97) );
  AOI22_X2 U_dfifo_U_dcore_U64 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_11_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[11]), .ZN(U_dfifo_U_dcore_n91) );
  AOI22_X2 U_dfifo_U_dcore_U63 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_13_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[13]), .ZN(U_dfifo_U_dcore_n95) );
  AOI22_X2 U_dfifo_U_dcore_U62 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_12_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[12]), .ZN(U_dfifo_U_dcore_n93) );
  AOI22_X2 U_dfifo_U_dcore_U61 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_23_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[23]), .ZN(U_dfifo_U_dcore_n66) );
  AOI22_X2 U_dfifo_U_dcore_U60 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_16_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[16]), .ZN(U_dfifo_U_dcore_n101) );
  AOI22_X2 U_dfifo_U_dcore_U59 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_15_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[15]), .ZN(U_dfifo_U_dcore_n99) );
  AOI22_X2 U_dfifo_U_dcore_U58 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_20_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[20]), .ZN(U_dfifo_U_dcore_n78) );
  AOI22_X2 U_dfifo_U_dcore_U57 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_19_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[19]), .ZN(U_dfifo_U_dcore_n82) );
  AOI22_X2 U_dfifo_U_dcore_U56 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_22_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[22]), .ZN(U_dfifo_U_dcore_n70) );
  AOI22_X2 U_dfifo_U_dcore_U55 ( .A1(U_dfifo_U_dcore_n126), .A2(
        U_dfifo_U_dcore_f_buf_data_21_), .B1(U_dfifo_U_dcore_n3), .B2(
        m_df_data_in[21]), .ZN(U_dfifo_U_dcore_n74) );
  AOI22_X2 U_dfifo_U_dcore_U54 ( .A1(U_dfifo_U_dcore_n3), .A2(m_double), .B1(
        U_dfifo_U_dcore_n127), .B2(U_dfifo_U_dcore_m_sf_data_out[1]), .ZN(
        U_dfifo_U_dcore_n123) );
  NAND2_X2 U_dfifo_U_dcore_U53 ( .A1(U_dfifo_n5), .A2(U_dfifo_U_dcore_n25), 
        .ZN(U_dfifo_U_dcore_n209) );
  NOR2_X1 U_dfifo_U_dcore_U52 ( .A1(m_two_to_one), .A2(U_dfifo_U_dcore_n106), 
        .ZN(U_dfifo_U_dcore_n50) );
  NAND2_X1 U_dfifo_U_dcore_U51 ( .A1(U_dfifo_U_dcore_m_sf_full), .A2(
        U_dfifo_U_dcore_n4), .ZN(U_dfifo_U_dcore_n22) );
  INV_X2 U_dfifo_U_dcore_U50 ( .A(U_dfifo_U_dcore_m_sf_full), .ZN(
        U_dfifo_U_dcore_n24) );
  INV_X2 U_dfifo_U_dcore_U49 ( .A(U_dfifo_n5), .ZN(U_dfifo_U_dcore_n26) );
  NAND2_X1 U_dfifo_U_dcore_U48 ( .A1(U_dfifo_U_dcore_n51), .A2(hiu_data[26]), 
        .ZN(U_dfifo_U_dcore_n76) );
  NOR2_X1 U_dfifo_U_dcore_U47 ( .A1(m_df_push_n), .A2(U_dfifo_U_dcore_n27), 
        .ZN(U_dfifo_U_dcore_n_empty) );
  NAND2_X1 U_dfifo_U_dcore_U46 ( .A1(U_dfifo_U_dcore_n51), .A2(hiu_data[31]), 
        .ZN(U_dfifo_U_dcore_n56) );
  NAND2_X1 U_dfifo_U_dcore_U45 ( .A1(U_dfifo_U_dcore_n51), .A2(hiu_data[25]), 
        .ZN(U_dfifo_U_dcore_n80) );
  NAND2_X1 U_dfifo_U_dcore_U44 ( .A1(U_dfifo_U_dcore_n51), .A2(hiu_data[30]), 
        .ZN(U_dfifo_U_dcore_n60) );
  NAND2_X1 U_dfifo_U_dcore_U43 ( .A1(U_dfifo_U_dcore_n51), .A2(hiu_data[29]), 
        .ZN(U_dfifo_U_dcore_n64) );
  NAND2_X1 U_dfifo_U_dcore_U42 ( .A1(U_dfifo_U_dcore_n51), .A2(hiu_data[27]), 
        .ZN(U_dfifo_U_dcore_n72) );
  NAND2_X1 U_dfifo_U_dcore_U41 ( .A1(U_dfifo_U_dcore_n51), .A2(hiu_data[28]), 
        .ZN(U_dfifo_U_dcore_n68) );
  NAND2_X1 U_dfifo_U_dcore_U40 ( .A1(hiu_data[24]), .A2(U_dfifo_U_dcore_n51), 
        .ZN(U_dfifo_U_dcore_n84) );
  INV_X2 U_dfifo_U_dcore_U39 ( .A(U_dfifo_U_dcore_n56), .ZN(
        U_dfifo_U_dcore_n57) );
  AOI22_X1 U_dfifo_U_dcore_U38 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[1]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[3]), .ZN(U_dfifo_U_dcore_n34) );
  INV_X2 U_dfifo_U_dcore_U37 ( .A(U_dfifo_U_dcore_n72), .ZN(
        U_dfifo_U_dcore_n73) );
  AOI22_X1 U_dfifo_U_dcore_U36 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[0]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[2]), .ZN(U_dfifo_U_dcore_n31) );
  INV_X2 U_dfifo_U_dcore_U35 ( .A(U_dfifo_U_dcore_n68), .ZN(
        U_dfifo_U_dcore_n69) );
  AOI22_X1 U_dfifo_U_dcore_U34 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[9]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[11]), .ZN(U_dfifo_U_dcore_n92) );
  AOI22_X1 U_dfifo_U_dcore_U33 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[7]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[9]), .ZN(U_dfifo_U_dcore_n54) );
  AOI22_X1 U_dfifo_U_dcore_U32 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[10]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[12]), .ZN(U_dfifo_U_dcore_n94) );
  AOI22_X1 U_dfifo_U_dcore_U31 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[8]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[10]), .ZN(U_dfifo_U_dcore_n90) );
  AOI22_X1 U_dfifo_U_dcore_U30 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[6]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[8]), .ZN(U_dfifo_U_dcore_n49) );
  INV_X2 U_dfifo_U_dcore_U29 ( .A(U_dfifo_U_dcore_n84), .ZN(
        U_dfifo_U_dcore_n85) );
  AOI22_X1 U_dfifo_U_dcore_U28 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[11]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[13]), .ZN(U_dfifo_U_dcore_n96) );
  AOI22_X1 U_dfifo_U_dcore_U27 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[5]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[7]), .ZN(U_dfifo_U_dcore_n46) );
  INV_X2 U_dfifo_U_dcore_U26 ( .A(U_dfifo_U_dcore_n60), .ZN(
        U_dfifo_U_dcore_n61) );
  INV_X2 U_dfifo_U_dcore_U25 ( .A(U_dfifo_U_dcore_n80), .ZN(
        U_dfifo_U_dcore_n81) );
  AOI22_X1 U_dfifo_U_dcore_U24 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[12]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[14]), .ZN(U_dfifo_U_dcore_n98) );
  AOI22_X1 U_dfifo_U_dcore_U23 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[2]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[4]), .ZN(U_dfifo_U_dcore_n37) );
  INV_X2 U_dfifo_U_dcore_U22 ( .A(U_dfifo_U_dcore_n76), .ZN(
        U_dfifo_U_dcore_n77) );
  AOI22_X1 U_dfifo_U_dcore_U21 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[4]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[6]), .ZN(U_dfifo_U_dcore_n43) );
  AOI22_X1 U_dfifo_U_dcore_U20 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[15]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[17]), .ZN(U_dfifo_U_dcore_n105) );
  AOI22_X1 U_dfifo_U_dcore_U19 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[13]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[15]), .ZN(U_dfifo_U_dcore_n100) );
  AOI22_X1 U_dfifo_U_dcore_U18 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[14]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[16]), .ZN(U_dfifo_U_dcore_n102) );
  AOI22_X1 U_dfifo_U_dcore_U17 ( .A1(U_dfifo_U_dcore_n103), .A2(
        U_dfifo_m_btm_data[3]), .B1(U_dfifo_U_dcore_n127), .B2(
        U_dfifo_U_dcore_m_sf_data_out[5]), .ZN(U_dfifo_U_dcore_n40) );
  INV_X2 U_dfifo_U_dcore_U16 ( .A(U_dfifo_U_dcore_n64), .ZN(
        U_dfifo_U_dcore_n65) );
  NAND2_X1 U_dfifo_U_dcore_U15 ( .A1(U_dfifo_U_dcore_n50), .A2(hiu_data[21]), 
        .ZN(U_dfifo_U_dcore_n44) );
  NAND2_X1 U_dfifo_U_dcore_U14 ( .A1(U_dfifo_U_dcore_n50), .A2(hiu_data[17]), 
        .ZN(U_dfifo_U_dcore_n32) );
  NAND2_X1 U_dfifo_U_dcore_U13 ( .A1(U_dfifo_U_dcore_n50), .A2(hiu_data[20]), 
        .ZN(U_dfifo_U_dcore_n41) );
  NAND2_X1 U_dfifo_U_dcore_U12 ( .A1(U_dfifo_U_dcore_n50), .A2(hiu_data[19]), 
        .ZN(U_dfifo_U_dcore_n38) );
  NAND2_X1 U_dfifo_U_dcore_U11 ( .A1(U_dfifo_U_dcore_n50), .A2(hiu_data[23]), 
        .ZN(U_dfifo_U_dcore_n52) );
  NAND2_X1 U_dfifo_U_dcore_U10 ( .A1(hiu_data[16]), .A2(U_dfifo_U_dcore_n50), 
        .ZN(U_dfifo_U_dcore_n29) );
  NAND2_X1 U_dfifo_U_dcore_U9 ( .A1(U_dfifo_U_dcore_n50), .A2(hiu_data[22]), 
        .ZN(U_dfifo_U_dcore_n47) );
  NAND2_X1 U_dfifo_U_dcore_U8 ( .A1(U_dfifo_U_dcore_n50), .A2(hiu_data[18]), 
        .ZN(U_dfifo_U_dcore_n35) );
  INV_X2 U_dfifo_U_dcore_U7 ( .A(U_dfifo_U_dcore_n103), .ZN(
        U_dfifo_U_dcore_n28) );
  INV_X4 U_dfifo_U_dcore_U6 ( .A(U_dfifo_U_dcore_n2), .ZN(U_dfifo_U_dcore_n1)
         );
  NAND2_X1 U_dfifo_U_dcore_U5 ( .A1(U_dfifo_U_dcore_n21), .A2(
        U_dfifo_U_dcore_n22), .ZN(U_dfifo_m_afull) );
  INV_X4 U_dfifo_U_dcore_U4 ( .A(U_dfifo_U_dcore_n23), .ZN(U_dfifo_m_full) );
  NAND2_X2 U_dfifo_U_dcore_U3 ( .A1(U_dfifo_U_dcore_m_sf_full), .A2(
        U_dfifo_U_dcore_f_buf_has_data), .ZN(U_dfifo_U_dcore_n23) );
  DFFR_X2 U_dfifo_U_dcore_f_data_out_reg_18_ ( .D(U_dfifo_U_dcore_n149), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[16]), .QN(U_dfifo_U_dcore_n13) );
  DFFR_X2 U_dfifo_U_dcore_f_data_out_reg_25_ ( .D(U_dfifo_U_dcore_n142), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[23]), .QN(U_dfifo_U_dcore_n14) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_2_ ( .D(U_dfifo_U_dcore_n134), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[0]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_3_ ( .D(U_dfifo_U_dcore_n135), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[1]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_4_ ( .D(U_dfifo_U_dcore_n136), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[2]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_5_ ( .D(U_dfifo_U_dcore_n137), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[3]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_6_ ( .D(U_dfifo_U_dcore_n138), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[4]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_7_ ( .D(U_dfifo_U_dcore_n139), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[5]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_8_ ( .D(U_dfifo_U_dcore_n140), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[6]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_9_ ( .D(U_dfifo_U_dcore_n141), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[7]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_24_ ( .D(U_dfifo_U_dcore_n143), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[22]), .QN(U_dfifo_U_dcore_n15) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_23_ ( .D(U_dfifo_U_dcore_n144), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[21]), .QN(U_dfifo_U_dcore_n16) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_22_ ( .D(U_dfifo_U_dcore_n145), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[20]), .QN(U_dfifo_U_dcore_n17) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_21_ ( .D(U_dfifo_U_dcore_n146), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[19]), .QN(U_dfifo_U_dcore_n18) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_20_ ( .D(U_dfifo_U_dcore_n147), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[18]), .QN(U_dfifo_U_dcore_n19) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_19_ ( .D(U_dfifo_U_dcore_n148), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[17]), .QN(U_dfifo_U_dcore_n20) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_10_ ( .D(U_dfifo_U_dcore_n150), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[8]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_11_ ( .D(U_dfifo_U_dcore_n151), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[9]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_12_ ( .D(U_dfifo_U_dcore_n152), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[10]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_13_ ( .D(U_dfifo_U_dcore_n153), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[11]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_14_ ( .D(U_dfifo_U_dcore_n154), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[12]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_15_ ( .D(U_dfifo_U_dcore_n155), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[13]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_16_ ( .D(U_dfifo_U_dcore_n156), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[14]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_17_ ( .D(U_dfifo_U_dcore_n157), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_btm_data[15]) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_26_ ( .D(U_dfifo_U_dcore_n158), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[24]), .QN(U_dfifo_U_dcore_n5) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_27_ ( .D(U_dfifo_U_dcore_n159), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[25]), .QN(U_dfifo_U_dcore_n6) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_28_ ( .D(U_dfifo_U_dcore_n160), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[26]), .QN(U_dfifo_U_dcore_n12) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_29_ ( .D(U_dfifo_U_dcore_n161), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[27]), .QN(U_dfifo_U_dcore_n7) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_30_ ( .D(U_dfifo_U_dcore_n162), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[28]), .QN(U_dfifo_U_dcore_n8) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_31_ ( .D(U_dfifo_U_dcore_n163), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[29]), .QN(U_dfifo_U_dcore_n9) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_32_ ( .D(U_dfifo_U_dcore_n164), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[30]), .QN(U_dfifo_U_dcore_n10) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_33_ ( .D(U_dfifo_U_dcore_n165), .CK(
        hclk), .RN(hresetn), .Q(hiu_data[31]), .QN(U_dfifo_U_dcore_n11) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_1_ ( .D(U_dfifo_U_dcore_n166), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_data_out_1_) );
  DFFR_X1 U_dfifo_U_dcore_f_data_out_reg_0_ ( .D(U_dfifo_U_dcore_n167), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_m_data_out_0_) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_has_data_reg ( .D(U_dfifo_U_dcore_n203), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_has_data), .QN(
        U_dfifo_U_dcore_n4) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_0_ ( .D(U_dfifo_U_dcore_n168), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_0_), .QN(n60) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_1_ ( .D(U_dfifo_U_dcore_n169), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_1_), .QN(n59) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_2_ ( .D(U_dfifo_U_dcore_n170), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_2_), .QN(n52) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_3_ ( .D(U_dfifo_U_dcore_n171), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_3_), .QN(n58) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_4_ ( .D(U_dfifo_U_dcore_n172), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_4_), .QN(n57) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_5_ ( .D(U_dfifo_U_dcore_n173), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_5_), .QN(n56) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_6_ ( .D(U_dfifo_U_dcore_n174), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_6_), .QN(n55) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_7_ ( .D(U_dfifo_U_dcore_n175), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_7_), .QN(n54) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_8_ ( .D(U_dfifo_U_dcore_n176), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_8_), .QN(n53) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_9_ ( .D(U_dfifo_U_dcore_n177), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_9_), .QN(n67) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_10_ ( .D(U_dfifo_U_dcore_n178), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_10_), .QN(n66) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_11_ ( .D(U_dfifo_U_dcore_n179), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_11_), .QN(n65) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_12_ ( .D(U_dfifo_U_dcore_n180), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_12_), .QN(n64) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_13_ ( .D(U_dfifo_U_dcore_n181), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_13_), .QN(n63) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_14_ ( .D(U_dfifo_U_dcore_n182), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_14_), .QN(n62) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_15_ ( .D(U_dfifo_U_dcore_n183), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_15_), .QN(n61) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_16_ ( .D(U_dfifo_U_dcore_n184), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_16_), .QN(n83) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_17_ ( .D(U_dfifo_U_dcore_n185), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_17_), .QN(n82) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_18_ ( .D(U_dfifo_U_dcore_n186), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_18_), .QN(n81) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_19_ ( .D(U_dfifo_U_dcore_n187), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_19_), .QN(n80) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_20_ ( .D(U_dfifo_U_dcore_n188), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_20_), .QN(n79) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_21_ ( .D(U_dfifo_U_dcore_n189), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_21_), .QN(n78) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_22_ ( .D(U_dfifo_U_dcore_n190), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_22_), .QN(n77) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_23_ ( .D(U_dfifo_U_dcore_n191), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_23_), .QN(n76) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_24_ ( .D(U_dfifo_U_dcore_n192), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_24_), .QN(n75) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_25_ ( .D(U_dfifo_U_dcore_n193), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_25_), .QN(n74) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_26_ ( .D(U_dfifo_U_dcore_n194), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_26_), .QN(n85) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_27_ ( .D(U_dfifo_U_dcore_n195), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_27_), .QN(n84) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_28_ ( .D(U_dfifo_U_dcore_n196), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_28_), .QN(n73) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_29_ ( .D(U_dfifo_U_dcore_n197), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_29_), .QN(n72) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_30_ ( .D(U_dfifo_U_dcore_n198), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_30_), .QN(n71) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_31_ ( .D(U_dfifo_U_dcore_n199), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_31_), .QN(n70) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_32_ ( .D(U_dfifo_U_dcore_n200), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_32_), .QN(n68) );
  DFFR_X1 U_dfifo_U_dcore_f_buf_data_reg_33_ ( .D(U_dfifo_U_dcore_n201), .CK(
        hclk), .RN(hresetn), .Q(U_dfifo_U_dcore_f_buf_data_33_), .QN(n69) );
  DFFS_X2 U_dfifo_U_dcore_f_empty_reg ( .D(U_dfifo_U_dcore_n_empty), .CK(hclk), 
        .SN(hresetn), .Q(U_dfifo_m_empty) );
  AOI22_X1 U_afifo_U_acore_U_sub_fifo_U276 ( .A1(
        U_afifo_U_acore_U_sub_fifo_count_1_), .A2(
        U_afifo_U_acore_U_sub_fifo_n371), .B1(
        U_afifo_U_acore_U_sub_fifo_count_0_), .B2(U_afifo_U_acore_n166), .ZN(
        U_afifo_U_acore_U_sub_fifo_n372) );
  NOR2_X1 U_afifo_U_acore_U_sub_fifo_U275 ( .A1(
        U_afifo_U_acore_U_sub_fifo_count_0_), .A2(U_afifo_U_acore_n166), .ZN(
        U_afifo_U_acore_U_sub_fifo_n371) );
  OAI21_X1 U_afifo_U_acore_U_sub_fifo_U274 ( .B1(
        U_afifo_U_acore_U_sub_fifo_n370), .B2(U_afifo_U_acore_U_sub_fifo_n11), 
        .A(U_afifo_U_acore_U_sub_fifo_n1), .ZN(U_afifo_U_acore_U_sub_fifo_n324) );
  OAI21_X1 U_afifo_U_acore_U_sub_fifo_U273 ( .B1(
        U_afifo_U_acore_U_sub_fifo_n370), .B2(U_afifo_U_acore_U_sub_fifo_n149), 
        .A(U_afifo_U_acore_U_sub_fifo_n369), .ZN(
        U_afifo_U_acore_U_sub_fifo_n323) );
  OAI21_X1 U_afifo_U_acore_U_sub_fifo_U272 ( .B1(U_afifo_U_acore_n166), .B2(
        U_afifo_U_acore_U_sub_fifo_n167), .A(
        U_afifo_U_acore_U_sub_fifo_count_1_), .ZN(
        U_afifo_U_acore_U_sub_fifo_n165) );
  NAND2_X1 U_afifo_U_acore_U_sub_fifo_U271 ( .A1(
        U_afifo_U_acore_U_sub_fifo_count_0_), .A2(U_afifo_U_acore_n166), .ZN(
        U_afifo_U_acore_U_sub_fifo_n166) );
  NAND3_X4 U_afifo_U_acore_U_sub_fifo_U270 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n149), .A2(
        U_afifo_U_acore_U_sub_fifo_in_ptr_1_), .A3(
        U_afifo_U_acore_U_sub_fifo_n370), .ZN(U_afifo_U_acore_U_sub_fifo_n169)
         );
  NAND3_X4 U_afifo_U_acore_U_sub_fifo_U269 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n11), .A2(U_afifo_U_acore_U_sub_fifo_n149), 
        .A3(U_afifo_U_acore_U_sub_fifo_n370), .ZN(
        U_afifo_U_acore_U_sub_fifo_n369) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U267 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n132), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n57), .C1(U_afifo_U_acore_U_sub_fifo_n7), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[18]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U266 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n122), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n77), .C1(U_afifo_U_acore_U_sub_fifo_n28), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[28]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U265 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n123), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n78), .C1(U_afifo_U_acore_U_sub_fifo_n29), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[27]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U264 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n125), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n56), .C1(U_afifo_U_acore_U_sub_fifo_n6), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[25]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U263 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n121), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n76), .C1(U_afifo_U_acore_U_sub_fifo_n27), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[29]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U262 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n124), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n79), .C1(U_afifo_U_acore_U_sub_fifo_n30), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[26]) );
  INV_X4 U_afifo_U_acore_U_sub_fifo_U261 ( .A(U_afifo_U_acore_U_sub_fifo_n162), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n150) );
  INV_X4 U_afifo_U_acore_U_sub_fifo_U260 ( .A(U_afifo_U_acore_U_sub_fifo_n150), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n151) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U259 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n126), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n80), .C1(U_afifo_U_acore_U_sub_fifo_n31), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[24]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U258 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n127), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n81), .C1(U_afifo_U_acore_U_sub_fifo_n32), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[23]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U257 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n128), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n82), .C1(U_afifo_U_acore_U_sub_fifo_n33), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[22]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U256 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n130), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n84), .C1(U_afifo_U_acore_U_sub_fifo_n35), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[20]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U255 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n131), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n85), .C1(U_afifo_U_acore_U_sub_fifo_n36), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[19]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U254 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n129), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n83), .C1(U_afifo_U_acore_U_sub_fifo_n34), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[21]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U253 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n116), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n72), .C1(U_afifo_U_acore_U_sub_fifo_n23), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[34]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U252 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n113), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n54), .C1(U_afifo_U_acore_U_sub_fifo_n4), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[37]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U251 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n114), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n70), .C1(U_afifo_U_acore_U_sub_fifo_n21), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[36]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U250 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n120), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n75), .C1(U_afifo_U_acore_U_sub_fifo_n26), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[30]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U249 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n112), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n69), .C1(U_afifo_U_acore_U_sub_fifo_n20), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[38]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U248 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n117), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n73), .C1(U_afifo_U_acore_U_sub_fifo_n24), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[33]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U247 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n115), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n71), .C1(U_afifo_U_acore_U_sub_fifo_n22), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[35]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U246 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n111), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n68), .C1(U_afifo_U_acore_U_sub_fifo_n19), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[39]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U245 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n119), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n74), .C1(U_afifo_U_acore_U_sub_fifo_n25), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[31]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U244 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n118), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n55), .C1(U_afifo_U_acore_U_sub_fifo_n5), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[32]) );
  INV_X4 U_afifo_U_acore_U_sub_fifo_U243 ( .A(U_afifo_U_acore_n166), .ZN(
        U_afifo_U_acore_U_sub_fifo_n168) );
  INV_X4 U_afifo_U_acore_U_sub_fifo_U242 ( .A(U_afifo_U_acore_n165), .ZN(
        U_afifo_U_acore_U_sub_fifo_n167) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U241 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n68), .B1(
        U_afifo_U_acore_U_sub_fifo_n17), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n231) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U239 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n31), .B1(
        U_afifo_U_acore_U_sub_fifo_n42), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n261) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U238 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n72), .B1(
        U_afifo_U_acore_U_sub_fifo_n19), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n233) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U237 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n90), .B1(
        U_afifo_U_acore_U_sub_fifo_n26), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n242) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U236 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n84), .B1(
        U_afifo_U_acore_U_sub_fifo_n24), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n239) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U235 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n78), .B1(
        U_afifo_U_acore_U_sub_fifo_n21), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n236) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U234 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n167), .B1(
        U_afifo_U_acore_U_sub_fifo_n7), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n254) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U233 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n70), .B1(
        U_afifo_U_acore_U_sub_fifo_n18), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n232) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U232 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n74), .B1(
        U_afifo_U_acore_U_sub_fifo_n20), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n234) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U231 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n82), .B1(
        U_afifo_U_acore_U_sub_fifo_n23), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n238) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U230 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n88), .B1(
        U_afifo_U_acore_U_sub_fifo_n25), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n241) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U229 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n86), .B1(
        U_afifo_U_acore_U_sub_fifo_n5), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n240) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U228 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n80), .B1(
        U_afifo_U_acore_U_sub_fifo_n22), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n237) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U226 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n30), .B1(
        U_afifo_U_acore_U_sub_fifo_n14), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n227) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U224 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n32), .B1(
        U_afifo_U_acore_U_sub_fifo_n43), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n263) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U222 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n29), .B1(
        U_afifo_U_acore_U_sub_fifo_n13), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n226) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U221 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n76), .B1(
        U_afifo_U_acore_U_sub_fifo_n4), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n235) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U219 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n162), .B1(
        U_afifo_U_acore_U_sub_fifo_n36), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n253) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U217 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n199), .B1(
        U_afifo_U_acore_U_sub_fifo_n38), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n256) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U215 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n156), .B1(
        U_afifo_U_acore_U_sub_fifo_n33), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n250) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U213 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n194), .B1(
        U_afifo_U_acore_U_sub_fifo_n16), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n230) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U211 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n203), .B1(
        U_afifo_U_acore_U_sub_fifo_n40), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n258) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U209 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n153), .B1(
        U_afifo_U_acore_U_sub_fifo_n32), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n249) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U207 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n158), .B1(
        U_afifo_U_acore_U_sub_fifo_n34), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n251) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U205 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n94), .B1(
        U_afifo_U_acore_U_sub_fifo_n27), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n243) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U203 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n100), .B1(
        U_afifo_U_acore_U_sub_fifo_n30), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n246) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U201 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n186), .B1(
        U_afifo_U_acore_U_sub_fifo_n61), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n225) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U199 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n160), .B1(
        U_afifo_U_acore_U_sub_fifo_n35), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n252) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U197 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n205), .B1(
        U_afifo_U_acore_U_sub_fifo_n8), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n259) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U195 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n96), .B1(
        U_afifo_U_acore_U_sub_fifo_n28), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n244) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U193 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n102), .B1(
        U_afifo_U_acore_U_sub_fifo_n6), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n247) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U191 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n207), .B1(
        U_afifo_U_acore_U_sub_fifo_n41), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n260) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U189 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n104), .B1(
        U_afifo_U_acore_U_sub_fifo_n31), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n248) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U187 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n201), .B1(
        U_afifo_U_acore_U_sub_fifo_n39), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n257) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U185 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n173), .B1(
        U_afifo_U_acore_U_sub_fifo_n44), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n264) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U183 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n192), .B1(
        U_afifo_U_acore_U_sub_fifo_n15), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n229) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U181 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n197), .B1(
        U_afifo_U_acore_U_sub_fifo_n37), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n255) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U179 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n98), .B1(
        U_afifo_U_acore_U_sub_fifo_n29), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n245) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U177 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n175), .B1(
        U_afifo_U_acore_U_sub_fifo_n45), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n265) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U175 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n190), .B1(
        U_afifo_U_acore_U_sub_fifo_n3), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n228) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U173 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n179), .B1(
        U_afifo_U_acore_U_sub_fifo_n9), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n267) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U171 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n177), .B1(
        U_afifo_U_acore_U_sub_fifo_n46), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n266) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U169 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n33), .B1(
        U_afifo_U_acore_U_sub_fifo_n48), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n269) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U168 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n92), .B1(
        U_afifo_U_acore_U_sub_fifo_n49), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n270) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U166 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n181), .B1(
        U_afifo_U_acore_U_sub_fifo_n47), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n268) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U164 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n210), .B1(
        U_afifo_U_acore_U_sub_fifo_n50), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n272) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U163 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n133), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n86), .C1(U_afifo_U_acore_U_sub_fifo_n37), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[17]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U162 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n134), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n87), .C1(U_afifo_U_acore_U_sub_fifo_n38), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[16]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U161 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n135), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n88), .C1(U_afifo_U_acore_U_sub_fifo_n39), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[15]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U160 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n136), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n89), .C1(U_afifo_U_acore_U_sub_fifo_n40), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[14]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U159 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n148), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n99), .C1(U_afifo_U_acore_U_sub_fifo_n50), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[0]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U158 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n137), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n58), .C1(U_afifo_U_acore_U_sub_fifo_n8), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[13]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U157 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n138), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n90), .C1(U_afifo_U_acore_U_sub_fifo_n41), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[12]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U156 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n107), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n64), .C1(U_afifo_U_acore_U_sub_fifo_n15), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[43]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U155 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n139), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n91), .C1(U_afifo_U_acore_U_sub_fifo_n42), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[11]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U154 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n104), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n62), .C1(U_afifo_U_acore_U_sub_fifo_n13), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[46]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U153 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n103), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n52), .C1(U_afifo_U_acore_U_sub_fifo_n61), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[47]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U152 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n108), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n65), .C1(U_afifo_U_acore_U_sub_fifo_n16), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[42]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U151 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n146), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n97), .C1(U_afifo_U_acore_U_sub_fifo_n48), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[3]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U150 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n144), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n59), .C1(U_afifo_U_acore_U_sub_fifo_n9), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[5]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U149 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n106), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n53), .C1(U_afifo_U_acore_U_sub_fifo_n3), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[44]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U148 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n145), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n96), .C1(U_afifo_U_acore_U_sub_fifo_n47), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[4]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U147 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n140), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n92), .C1(U_afifo_U_acore_U_sub_fifo_n43), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[9]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U146 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n105), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n63), .C1(U_afifo_U_acore_U_sub_fifo_n14), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[45]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U145 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n102), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n51), .C1(U_afifo_U_acore_U_sub_fifo_n60), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[48]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U144 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n142), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n94), .C1(U_afifo_U_acore_U_sub_fifo_n45), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[7]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U143 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n2), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n101), .C1(U_afifo_U_acore_U_sub_fifo_n12), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[49]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U142 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n143), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n95), .C1(U_afifo_U_acore_U_sub_fifo_n46), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[6]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U141 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n141), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n93), .C1(U_afifo_U_acore_U_sub_fifo_n44), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[8]) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U139 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n28), .B1(
        U_afifo_U_acore_U_sub_fifo_n12), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n223) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U137 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n153), .A2(U_afifo_U_acore_n184), .B1(
        U_afifo_U_acore_U_sub_fifo_n60), .B2(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n224) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U136 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n109), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n66), .C1(U_afifo_U_acore_U_sub_fifo_n17), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[41]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U135 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n151), .A2(U_afifo_U_acore_U_sub_fifo_n110), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n67), .C1(U_afifo_U_acore_U_sub_fifo_n18), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[40]) );
  OAI222_X2 U_afifo_U_acore_U_sub_fifo_U134 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n162), .A2(U_afifo_U_acore_U_sub_fifo_n147), 
        .B1(U_afifo_U_acore_U_sub_fifo_n163), .B2(
        U_afifo_U_acore_U_sub_fifo_n98), .C1(U_afifo_U_acore_U_sub_fifo_n49), 
        .C2(U_afifo_U_acore_U_sub_fifo_n161), .ZN(
        U_afifo_U_acore_m_sf_data_out[2]) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U133 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n80), .B1(
        U_afifo_U_acore_U_sub_fifo_n71), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n187) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U132 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n90), .B1(
        U_afifo_U_acore_U_sub_fifo_n75), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n192) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U131 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n72), .B1(
        U_afifo_U_acore_U_sub_fifo_n68), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n183) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U130 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n86), .B1(
        U_afifo_U_acore_U_sub_fifo_n55), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n190) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U129 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n82), .B1(
        U_afifo_U_acore_U_sub_fifo_n72), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n188) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U128 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n68), .B1(
        U_afifo_U_acore_U_sub_fifo_n66), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n181) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U127 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n78), .B1(
        U_afifo_U_acore_U_sub_fifo_n70), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n186) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U126 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n76), .B1(
        U_afifo_U_acore_U_sub_fifo_n54), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n185) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U125 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n74), .B1(
        U_afifo_U_acore_U_sub_fifo_n69), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n184) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U124 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n70), .B1(
        U_afifo_U_acore_U_sub_fifo_n67), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n182) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U123 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n88), .B1(
        U_afifo_U_acore_U_sub_fifo_n74), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n191) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U122 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n28), .B1(
        U_afifo_U_acore_U_sub_fifo_n101), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n173) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U121 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n158), .B1(
        U_afifo_U_acore_U_sub_fifo_n83), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n201) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U120 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n194), .B1(
        U_afifo_U_acore_U_sub_fifo_n65), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n180) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U119 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n205), .B1(
        U_afifo_U_acore_U_sub_fifo_n58), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n209) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U118 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n192), .B1(
        U_afifo_U_acore_U_sub_fifo_n64), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n179) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U117 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n190), .B1(
        U_afifo_U_acore_U_sub_fifo_n53), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n178) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U116 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n156), .B1(
        U_afifo_U_acore_U_sub_fifo_n82), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n200) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U115 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n30), .B1(
        U_afifo_U_acore_U_sub_fifo_n63), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n177) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U114 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n29), .B1(
        U_afifo_U_acore_U_sub_fifo_n62), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n176) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U113 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n186), .B1(
        U_afifo_U_acore_U_sub_fifo_n52), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n175) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U112 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n184), .B1(
        U_afifo_U_acore_U_sub_fifo_n51), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n174) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U111 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n94), .B1(
        U_afifo_U_acore_U_sub_fifo_n76), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n193) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U110 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n96), .B1(
        U_afifo_U_acore_U_sub_fifo_n77), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n194) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U109 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n31), .B1(
        U_afifo_U_acore_U_sub_fifo_n91), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n211) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U108 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n104), .B1(
        U_afifo_U_acore_U_sub_fifo_n80), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n198) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U107 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n98), .B1(
        U_afifo_U_acore_U_sub_fifo_n78), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n195) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U106 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n33), .B1(
        U_afifo_U_acore_U_sub_fifo_n97), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n219) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U105 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n153), .B1(
        U_afifo_U_acore_U_sub_fifo_n81), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n199) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U104 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n100), .B1(
        U_afifo_U_acore_U_sub_fifo_n79), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n196) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U103 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n203), .B1(
        U_afifo_U_acore_U_sub_fifo_n89), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n208) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U102 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n179), .B1(
        U_afifo_U_acore_U_sub_fifo_n59), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n217) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U101 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n207), .B1(
        U_afifo_U_acore_U_sub_fifo_n90), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n210) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U100 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n160), .B1(
        U_afifo_U_acore_U_sub_fifo_n84), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n202) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U99 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n162), .B1(
        U_afifo_U_acore_U_sub_fifo_n85), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n203) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U98 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n177), .B1(
        U_afifo_U_acore_U_sub_fifo_n95), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n216) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U97 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n167), .B1(
        U_afifo_U_acore_U_sub_fifo_n57), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n204) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U96 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n197), .B1(
        U_afifo_U_acore_U_sub_fifo_n86), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n205) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U95 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n175), .B1(
        U_afifo_U_acore_U_sub_fifo_n94), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n215) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U94 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n199), .B1(
        U_afifo_U_acore_U_sub_fifo_n87), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n206) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U93 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n173), .B1(
        U_afifo_U_acore_U_sub_fifo_n93), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n214) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U92 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n201), .B1(
        U_afifo_U_acore_U_sub_fifo_n88), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n207) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U91 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n32), .B1(
        U_afifo_U_acore_U_sub_fifo_n92), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n213) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U90 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n92), .B1(
        U_afifo_U_acore_U_sub_fifo_n98), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n220) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U89 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n84), .B1(
        U_afifo_U_acore_U_sub_fifo_n73), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n189) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U88 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n210), .B1(
        U_afifo_U_acore_U_sub_fifo_n99), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n222) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U87 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n181), .B1(
        U_afifo_U_acore_U_sub_fifo_n96), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n218) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U86 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n212), .A2(U_afifo_U_acore_n102), .B1(
        U_afifo_U_acore_U_sub_fifo_n56), .B2(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n197) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U85 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n33), .B1(
        U_afifo_U_acore_U_sub_fifo_n146), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n319) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U84 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n68), .B1(
        U_afifo_U_acore_U_sub_fifo_n109), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n281) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U83 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n210), .B1(
        U_afifo_U_acore_U_sub_fifo_n148), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n322) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U82 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n192), .B1(
        U_afifo_U_acore_U_sub_fifo_n107), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n279) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U81 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n179), .B1(
        U_afifo_U_acore_U_sub_fifo_n144), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n317) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U80 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n29), .B1(
        U_afifo_U_acore_U_sub_fifo_n104), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n276) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U79 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n186), .B1(
        U_afifo_U_acore_U_sub_fifo_n103), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n275) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U78 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n181), .B1(
        U_afifo_U_acore_U_sub_fifo_n145), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n318) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U77 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n190), .B1(
        U_afifo_U_acore_U_sub_fifo_n106), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n278) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U76 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n76), .B1(
        U_afifo_U_acore_U_sub_fifo_n113), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n285) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U75 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n194), .B1(
        U_afifo_U_acore_U_sub_fifo_n108), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n280) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U74 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n92), .B1(
        U_afifo_U_acore_U_sub_fifo_n147), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n320) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U73 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n78), .B1(
        U_afifo_U_acore_U_sub_fifo_n114), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n286) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U72 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n72), .B1(
        U_afifo_U_acore_U_sub_fifo_n111), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n283) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U71 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n74), .B1(
        U_afifo_U_acore_U_sub_fifo_n112), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n284) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U70 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n177), .B1(
        U_afifo_U_acore_U_sub_fifo_n143), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n316) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U69 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n70), .B1(
        U_afifo_U_acore_U_sub_fifo_n110), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n282) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U68 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n28), .B1(
        U_afifo_U_acore_U_sub_fifo_n2), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n273) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U67 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n84), .B1(
        U_afifo_U_acore_U_sub_fifo_n117), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n289) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U66 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n100), .B1(
        U_afifo_U_acore_U_sub_fifo_n124), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n296) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U65 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n205), .B1(
        U_afifo_U_acore_U_sub_fifo_n137), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n309) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U64 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n86), .B1(
        U_afifo_U_acore_U_sub_fifo_n118), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n290) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U63 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n158), .B1(
        U_afifo_U_acore_U_sub_fifo_n129), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n301) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U62 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n162), .B1(
        U_afifo_U_acore_U_sub_fifo_n131), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n303) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U61 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n94), .B1(
        U_afifo_U_acore_U_sub_fifo_n121), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n293) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U60 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n90), .B1(
        U_afifo_U_acore_U_sub_fifo_n120), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n292) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U59 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n104), .B1(
        U_afifo_U_acore_U_sub_fifo_n126), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n298) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U58 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n201), .B1(
        U_afifo_U_acore_U_sub_fifo_n135), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n307) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U57 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n88), .B1(
        U_afifo_U_acore_U_sub_fifo_n119), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n291) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U56 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n173), .B1(
        U_afifo_U_acore_U_sub_fifo_n141), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n314) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U55 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n203), .B1(
        U_afifo_U_acore_U_sub_fifo_n136), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n308) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U54 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n156), .B1(
        U_afifo_U_acore_U_sub_fifo_n128), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n300) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U53 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n80), .B1(
        U_afifo_U_acore_U_sub_fifo_n115), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n287) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U52 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n197), .B1(
        U_afifo_U_acore_U_sub_fifo_n133), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n305) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U51 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n167), .B1(
        U_afifo_U_acore_U_sub_fifo_n132), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n304) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U50 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n82), .B1(
        U_afifo_U_acore_U_sub_fifo_n116), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n288) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U49 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n102), .B1(
        U_afifo_U_acore_U_sub_fifo_n125), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n297) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U48 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n153), .B1(
        U_afifo_U_acore_U_sub_fifo_n127), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n299) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U47 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n175), .B1(
        U_afifo_U_acore_U_sub_fifo_n142), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n315) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U46 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n184), .B1(
        U_afifo_U_acore_U_sub_fifo_n102), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n274) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U45 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n96), .B1(
        U_afifo_U_acore_U_sub_fifo_n122), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n294) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U44 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n31), .B1(
        U_afifo_U_acore_U_sub_fifo_n139), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n311) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U43 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n32), .B1(
        U_afifo_U_acore_U_sub_fifo_n140), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n313) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U42 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n160), .B1(
        U_afifo_U_acore_U_sub_fifo_n130), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n302) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U41 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n207), .B1(
        U_afifo_U_acore_U_sub_fifo_n138), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n310) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U40 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n98), .B1(
        U_afifo_U_acore_U_sub_fifo_n123), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n295) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U39 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n30), .B1(
        U_afifo_U_acore_U_sub_fifo_n105), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n277) );
  AOI22_X2 U_afifo_U_acore_U_sub_fifo_U38 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n152), .A2(U_afifo_U_acore_n199), .B1(
        U_afifo_U_acore_U_sub_fifo_n134), .B2(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n306) );
  NOR2_X2 U_afifo_U_acore_U_sub_fifo_U37 ( .A1(U_afifo_U_acore_n166), .A2(
        U_afifo_U_acore_n2), .ZN(U_afifo_U_acore_U_sub_fifo_n160) );
  OAI21_X2 U_afifo_U_acore_U_sub_fifo_U36 ( .B1(
        U_afifo_U_acore_U_sub_fifo_n160), .B2(U_afifo_U_acore_U_sub_fifo_n163), 
        .A(U_afifo_U_acore_U_sub_fifo_n159), .ZN(
        U_afifo_U_acore_U_sub_fifo_n171) );
  NAND2_X2 U_afifo_U_acore_U_sub_fifo_U35 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n160), .A2(U_afifo_U_acore_U_sub_fifo_n150), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n158) );
  OAI21_X2 U_afifo_U_acore_U_sub_fifo_U34 ( .B1(
        U_afifo_U_acore_U_sub_fifo_n160), .B2(U_afifo_U_acore_U_sub_fifo_n161), 
        .A(U_afifo_U_acore_U_sub_fifo_n158), .ZN(
        U_afifo_U_acore_U_sub_fifo_n170) );
  OAI211_X1 U_afifo_U_acore_U_sub_fifo_U32 ( .C1(U_afifo_U_acore_n165), .C2(
        U_afifo_U_acore_U_sub_fifo_n166), .A(U_afifo_U_acore_U_sub_fifo_n165), 
        .B(U_afifo_U_acore_m_sf_full), .ZN(U_afifo_U_acore_U_sub_fifo_n172) );
  INV_X8 U_afifo_U_acore_U_sub_fifo_U30 ( .A(U_afifo_U_acore_U_sub_fifo_n1), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n153) );
  INV_X8 U_afifo_U_acore_U_sub_fifo_U28 ( .A(
        U_afifo_U_acore_U_sub_fifo_out_ptr_0_), .ZN(
        U_afifo_U_acore_U_sub_fifo_n161) );
  INV_X8 U_afifo_U_acore_U_sub_fifo_U27 ( .A(
        U_afifo_U_acore_U_sub_fifo_out_ptr_1_), .ZN(
        U_afifo_U_acore_U_sub_fifo_n163) );
  INV_X8 U_afifo_U_acore_U_sub_fifo_U26 ( .A(U_afifo_U_acore_U_sub_fifo_n169), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n212) );
  NAND2_X4 U_afifo_U_acore_U_sub_fifo_U25 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n161), .A2(U_afifo_U_acore_U_sub_fifo_n163), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n162) );
  AND2_X4 U_afifo_U_acore_U_sub_fifo_U24 ( .A1(U_afifo_U_acore_U_sub_fifo_n100), .A2(U_afifo_U_acore_U_sub_fifo_n10), .ZN(U_afifo_U_acore_n2) );
  NAND2_X2 U_afifo_U_acore_U_sub_fifo_U23 ( .A1(
        U_afifo_U_acore_U_sub_fifo_count_1_), .A2(
        U_afifo_U_acore_U_sub_fifo_count_0_), .ZN(U_afifo_U_acore_m_sf_full)
         );
  OAI21_X2 U_afifo_U_acore_U_sub_fifo_U22 ( .B1(U_afifo_U_acore_m_sf_full), 
        .B2(U_afifo_U_acore_U_sub_fifo_n168), .A(
        U_afifo_U_acore_U_sub_fifo_n167), .ZN(U_afifo_U_acore_U_sub_fifo_n373)
         );
  NAND3_X1 U_afifo_U_acore_U_sub_fifo_U21 ( .A1(
        U_afifo_U_acore_U_sub_fifo_n160), .A2(U_afifo_U_acore_U_sub_fifo_n163), 
        .A3(U_afifo_U_acore_U_sub_fifo_out_ptr_0_), .ZN(
        U_afifo_U_acore_U_sub_fifo_n159) );
  INV_X4 U_afifo_U_acore_U_sub_fifo_U20 ( .A(U_afifo_U_acore_U_sub_fifo_n373), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n370) );
  XOR2_X1 U_afifo_U_acore_U_sub_fifo_U19 ( .A(U_afifo_U_acore_U_sub_fifo_n373), 
        .B(U_afifo_U_acore_U_sub_fifo_n372), .Z(
        U_afifo_U_acore_U_sub_fifo_n325) );
  INV_X8 U_afifo_U_acore_U_sub_fifo_U4 ( .A(U_afifo_U_acore_U_sub_fifo_n369), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n152) );
  OR3_X4 U_afifo_U_acore_U_sub_fifo_U3 ( .A1(
        U_afifo_U_acore_U_sub_fifo_in_ptr_1_), .A2(
        U_afifo_U_acore_U_sub_fifo_n373), .A3(U_afifo_U_acore_U_sub_fifo_n149), 
        .ZN(U_afifo_U_acore_U_sub_fifo_n1) );
  DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__0_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n272), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n50) );
  DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__2_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n270), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n49) );
  DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__3_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n269), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n48) );
  DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__4_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n268), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n47) );
  DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__5_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n267), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n9) );
  DFFR_X2 U_afifo_U_acore_U_sub_fifo_mem_reg_1__6_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n266), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n46) );
  DFFR_X2 U_afifo_U_acore_U_sub_fifo_in_ptr_reg_0_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n323), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n149) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_out_ptr_reg_0_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n170), .CK(hclk), .RN(hresetn), .Q(
        U_afifo_U_acore_U_sub_fifo_out_ptr_0_) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_out_ptr_reg_1_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n171), .CK(hclk), .RN(hresetn), .Q(
        U_afifo_U_acore_U_sub_fifo_out_ptr_1_) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_count_reg_1_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n172), .CK(hclk), .RN(hresetn), .Q(
        U_afifo_U_acore_U_sub_fifo_count_1_), .QN(
        U_afifo_U_acore_U_sub_fifo_n100) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__49_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n173), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n101) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__48_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n174), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n51) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__47_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n175), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n52) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__46_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n176), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n62) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__45_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n177), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n63) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__44_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n178), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n53) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__43_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n179), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n64) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__42_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n180), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n65) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__41_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n181), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n66) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__40_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n182), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n67) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__39_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n183), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n68) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__38_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n184), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n69) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__37_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n185), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n54) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__36_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n186), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n70) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__35_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n187), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n71) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__34_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n188), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n72) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__33_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n189), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n73) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__32_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n190), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n55) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__31_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n191), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n74) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__30_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n192), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n75) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__29_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n193), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n76) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__28_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n194), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n77) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__27_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n195), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n78) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__26_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n196), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n79) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__25_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n197), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n56) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__24_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n198), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n80) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__23_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n199), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n81) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__22_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n200), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n82) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__21_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n201), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n83) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__20_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n202), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n84) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__19_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n203), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n85) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__18_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n204), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n57) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__17_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n205), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n86) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__16_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n206), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n87) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__15_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n207), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n88) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__14_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n208), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n89) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__13_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n209), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n58) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__12_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n210), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n90) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__11_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n211), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n91) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__9_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n213), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n92) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__8_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n214), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n93) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__7_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n215), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n94) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__6_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n216), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n95) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__5_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n217), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n59) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__4_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n218), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n96) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__3_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n219), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n97) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__2_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n220), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n98) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_2__0_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n222), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n99) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__49_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n223), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n12) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__48_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n224), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n60) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__47_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n225), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n61) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__46_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n226), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n13) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__45_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n227), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n14) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__44_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n228), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n3) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__43_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n229), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n15) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__42_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n230), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n16) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__41_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n231), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n17) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__40_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n232), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n18) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__39_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n233), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n19) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__38_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n234), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n20) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__37_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n235), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n4) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__36_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n236), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n21) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__35_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n237), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n22) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__34_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n238), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n23) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__33_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n239), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n24) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__32_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n240), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n5) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__31_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n241), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n25) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__30_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n242), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n26) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__29_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n243), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n27) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__28_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n244), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n28) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__27_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n245), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n29) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__26_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n246), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n30) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__25_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n247), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n6) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__24_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n248), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n31) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__23_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n249), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n32) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__22_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n250), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n33) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__21_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n251), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n34) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__20_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n252), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n35) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__19_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n253), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n36) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__18_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n254), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n7) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__17_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n255), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n37) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__16_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n256), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n38) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__15_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n257), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n39) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__14_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n258), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n40) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__13_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n259), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n8) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__12_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n260), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n41) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__11_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n261), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n42) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__9_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n263), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n43) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__8_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n264), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n44) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_1__7_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n265), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n45) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__49_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n273), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n2) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__48_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n274), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n102) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__47_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n275), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n103) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__46_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n276), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n104) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__45_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n277), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n105) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__44_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n278), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n106) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__43_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n279), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n107) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__42_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n280), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n108) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__41_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n281), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n109) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__40_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n282), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n110) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__39_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n283), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n111) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__38_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n284), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n112) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__37_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n285), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n113) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__36_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n286), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n114) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__35_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n287), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n115) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__34_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n288), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n116) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__33_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n289), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n117) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__32_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n290), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n118) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__31_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n291), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n119) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__30_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n292), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n120) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__29_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n293), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n121) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__28_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n294), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n122) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__27_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n295), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n123) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__26_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n296), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n124) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__25_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n297), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n125) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__24_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n298), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n126) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__23_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n299), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n127) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__22_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n300), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n128) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__21_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n301), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n129) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__20_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n302), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n130) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__19_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n303), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n131) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__18_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n304), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n132) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__17_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n305), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n133) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__16_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n306), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n134) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__15_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n307), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n135) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__14_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n308), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n136) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__13_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n309), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n137) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__12_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n310), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n138) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__11_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n311), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n139) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__9_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n313), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n140) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__8_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n314), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n141) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__7_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n315), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n142) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__6_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n316), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n143) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__5_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n317), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n144) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__4_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n318), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n145) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__3_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n319), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n146) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__2_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n320), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n147) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_mem_reg_0__0_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n322), .CK(hclk), .RN(hresetn), .QN(
        U_afifo_U_acore_U_sub_fifo_n148) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_in_ptr_reg_1_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n324), .CK(hclk), .RN(hresetn), .Q(
        U_afifo_U_acore_U_sub_fifo_in_ptr_1_), .QN(
        U_afifo_U_acore_U_sub_fifo_n11) );
  DFFR_X1 U_afifo_U_acore_U_sub_fifo_count_reg_0_ ( .D(
        U_afifo_U_acore_U_sub_fifo_n325), .CK(hclk), .RN(hresetn), .Q(
        U_afifo_U_acore_U_sub_fifo_count_0_), .QN(
        U_afifo_U_acore_U_sub_fifo_n10) );
  OAI21_X1 U_dfifo_U_dcore_U_sub_fifo_U435 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_n603), .B2(U_dfifo_U_dcore_U_sub_fifo_n57), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n12), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n448) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U434 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n60), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n117), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n310) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U433 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n59), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n116), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n309) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U432 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n52), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n115), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n308) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U431 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n58), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n114), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n307) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U430 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n57), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n113), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n306) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U429 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n56), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n112), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n305) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U428 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n55), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n111), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n304) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U427 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n54), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n110), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n303) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U426 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n53), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n109), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n302) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U425 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n67), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n108), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n301) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U424 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n66), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n107), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n300) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U423 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n65), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n106), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n299) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U422 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n64), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n105), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n298) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U421 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n63), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n104), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n297) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U420 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n62), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n103), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n296) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U419 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n61), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n102), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n295) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U418 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n83), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n101), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n294) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U417 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n82), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n100), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n293) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U416 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n81), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n99), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n292) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U415 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n80), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n98), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n291) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U414 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n79), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n97), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n290) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U413 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n78), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n96), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n289) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U412 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n77), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n95), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n288) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U411 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n76), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n94), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n287) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U410 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n75), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n93), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n286) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U409 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n74), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n92), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n285) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U408 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n85), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n91), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n284) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U407 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n84), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n90), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n283) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U406 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n73), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n89), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n282) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U405 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n72), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n88), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n281) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U404 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n71), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n87), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n280) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U403 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n70), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n86), .B2(U_dfifo_U_dcore_U_sub_fifo_n6), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n279) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U402 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n60), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n52), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n276) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U401 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n59), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n51), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n275) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U400 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n52), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n50), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n274) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U399 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n58), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n49), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n273) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U398 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n57), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n48), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n272) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U397 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n56), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n47), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n271) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U396 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n55), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n46), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n270) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U395 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n54), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n45), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n269) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U394 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n53), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n44), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n268) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U393 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n67), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n43), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n267) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U392 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n66), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n42), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n266) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U391 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n65), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n41), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n265) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U390 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n64), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n40), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n264) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U389 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n63), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n39), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n263) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U388 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n62), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n38), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n262) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U387 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n61), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n37), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n261) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U386 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n83), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n36), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n260) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U385 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n82), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n35), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n259) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U384 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n81), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n34), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n258) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U383 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n80), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n33), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n257) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U382 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n79), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n32), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n256) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U381 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n78), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n31), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n255) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U380 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n77), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n30), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n254) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U379 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n76), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n29), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n253) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U378 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n75), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n28), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n252) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U377 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n74), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n27), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n251) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U376 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n85), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n26), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n250) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U375 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n84), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n25), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n249) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U374 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n73), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n24), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n248) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U373 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n72), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n23), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n247) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U372 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n71), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n22), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n246) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U371 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n70), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n21), .B2(U_dfifo_U_dcore_U_sub_fifo_n7), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n245) );
  OR2_X4 U_dfifo_U_dcore_U_sub_fifo_U370 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n602), .A2(U_dfifo_U_dcore_U_sub_fifo_n567), .ZN(U_dfifo_U_dcore_U_sub_fifo_n12) );
  OR2_X4 U_dfifo_U_dcore_U_sub_fifo_U369 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n604), .A2(U_dfifo_U_dcore_U_sub_fifo_n567), .ZN(U_dfifo_U_dcore_U_sub_fifo_n11) );
  OR3_X4 U_dfifo_U_dcore_U_sub_fifo_U368 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_2_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_), .A3(
        U_dfifo_U_dcore_U_sub_fifo_n602), .ZN(U_dfifo_U_dcore_U_sub_fifo_n10)
         );
  OR3_X4 U_dfifo_U_dcore_U_sub_fifo_U367 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_2_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_), .A3(
        U_dfifo_U_dcore_U_sub_fifo_n604), .ZN(U_dfifo_U_dcore_U_sub_fifo_n9)
         );
  AND2_X4 U_dfifo_U_dcore_U_sub_fifo_U366 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n460), .A2(U_dfifo_U_dcore_U_sub_fifo_n18), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n562) );
  AOI21_X1 U_dfifo_U_dcore_U_sub_fifo_U365 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_n13), .B2(U_dfifo_U_dcore_U_sub_fifo_n54), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n17), .ZN(U_dfifo_U_dcore_m_sf_afull) );
  INV_X1 U_dfifo_U_dcore_U_sub_fifo_U364 ( .A(U_dfifo_U_dcore_U_sub_fifo_n602), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n603) );
  NOR3_X1 U_dfifo_U_dcore_U_sub_fifo_U363 ( .A1(U_dfifo_U_dcore_n208), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n609), .A3(U_dfifo_U_dcore_U_sub_fifo_n13), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n456) );
  OAI21_X1 U_dfifo_U_dcore_U_sub_fifo_U362 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_n458), .B2(U_dfifo_U_dcore_U_sub_fifo_n55), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n604), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n449) );
  NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U359 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_1_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n460) );
  NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U358 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n56), .ZN(U_dfifo_U_dcore_U_sub_fifo_n560)
         );
  NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U357 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n18), .A2(U_dfifo_U_dcore_U_sub_fifo_n56), .ZN(U_dfifo_U_dcore_U_sub_fifo_n605) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U356 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__25_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__25_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n605), .ZN(U_dfifo_U_dcore_U_sub_fifo_n514)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U355 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n27), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n92), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n512)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U354 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__25_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n512), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n513) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U353 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__18_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__18_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n490)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U352 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n34), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n99), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n488)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U351 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__18_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n488), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n489) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U350 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__10_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__10_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n466)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U349 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n42), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n107), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n464)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U348 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__10_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n464), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n465) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U347 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n73), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n466), .B(
        U_dfifo_U_dcore_U_sub_fifo_n465), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[10]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U346 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__17_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__17_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n487)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U345 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n35), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n100), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n485)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U344 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__17_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n485), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n486) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U343 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n66), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n487), .B(
        U_dfifo_U_dcore_U_sub_fifo_n486), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[17]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U342 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__9_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__9_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n564)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U341 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n43), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n108), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n561)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U340 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__9_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n561), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n563) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U339 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__2_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__2_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n529)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U338 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n50), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n115), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n527)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U337 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__2_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n527), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n528) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U336 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__24_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__24_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n605), .ZN(U_dfifo_U_dcore_U_sub_fifo_n511)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U335 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n28), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n93), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n509)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U334 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__24_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n509), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n510) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U333 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__14_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__14_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n478)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U332 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n38), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n103), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n476)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U331 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__14_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n476), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n477) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U330 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n69), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n478), .B(
        U_dfifo_U_dcore_U_sub_fifo_n477), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[14]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U329 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__11_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__11_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n469)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U328 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n41), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n106), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n467)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U327 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__11_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n467), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n468) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U326 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n72), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n469), .B(
        U_dfifo_U_dcore_U_sub_fifo_n468), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[11]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U325 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__13_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__13_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n475)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U324 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n39), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n104), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n473)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U323 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__13_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n473), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n474) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U322 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n70), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n475), .B(
        U_dfifo_U_dcore_U_sub_fifo_n474), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[13]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U321 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__12_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__12_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n472)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U320 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n40), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n105), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n470)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U319 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__12_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n470), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n471) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U318 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n71), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n472), .B(
        U_dfifo_U_dcore_U_sub_fifo_n471), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[12]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U317 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__33_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__33_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n541)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U316 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n19), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n84), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n539)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U315 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__33_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n539), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n540) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U314 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n58), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n541), .B(
        U_dfifo_U_dcore_U_sub_fifo_n540), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[33]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U313 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__26_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__26_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n517)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U312 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n26), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n91), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n515)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U311 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__26_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n515), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n516) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U310 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n65), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n517), .B(
        U_dfifo_U_dcore_U_sub_fifo_n516), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[26]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U309 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__23_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__23_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n605), .ZN(U_dfifo_U_dcore_U_sub_fifo_n508)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U308 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n29), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n94), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n506)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U307 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__23_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n506), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n507) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U306 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__16_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__16_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n484)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U305 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n36), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n101), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n482)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U304 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__16_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n482), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n483) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U303 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n67), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n484), .B(
        U_dfifo_U_dcore_U_sub_fifo_n483), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[16]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U302 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__15_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__15_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n481)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U301 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n37), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n102), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n479)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U300 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__15_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n479), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n480) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U299 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n68), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n481), .B(
        U_dfifo_U_dcore_U_sub_fifo_n480), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[15]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U298 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__20_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__20_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n605), .ZN(U_dfifo_U_dcore_U_sub_fifo_n499)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U297 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n32), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n97), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n497)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U296 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__20_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n497), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n498) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U295 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__19_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__19_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n493)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U294 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n33), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n98), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n491)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U293 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__19_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n491), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n492) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U292 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__22_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__22_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n605), .ZN(U_dfifo_U_dcore_U_sub_fifo_n505)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U291 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n30), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n95), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n503)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U290 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__22_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n503), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n504) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U289 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__21_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__21_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n605), .ZN(U_dfifo_U_dcore_U_sub_fifo_n502)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U288 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n31), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n96), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n500)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U287 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__21_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n500), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n501) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U286 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__8_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__8_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n559)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U285 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n44), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n109), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n557)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U284 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__8_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n557), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n558) );
  NAND2_X2 U_dfifo_U_dcore_U_sub_fifo_U282 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n458), .A2(U_dfifo_U_dcore_U_sub_fifo_n55), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n604) );
  NAND2_X2 U_dfifo_U_dcore_U_sub_fifo_U249 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n458), .A2(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_0_), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n602) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U248 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__5_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__5_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n550)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U247 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n47), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n112), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n548)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U246 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__5_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n548), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n549) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U245 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__4_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__4_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n547)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U244 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n48), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n113), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n545)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U243 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__4_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n545), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n546) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U242 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__7_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__7_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n556)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U241 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n45), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n110), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n554)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U240 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__7_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n554), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n555) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U239 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__6_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__6_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n553)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U238 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n46), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n111), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n551)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U237 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__6_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n551), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n552) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U236 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__3_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__3_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n544)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U235 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n49), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n114), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n542)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U234 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__3_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n542), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n543) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U233 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__31_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__31_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n535)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U232 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n21), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n86), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n533)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U231 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__31_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n533), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n534) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U230 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n60), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n535), .B(
        U_dfifo_U_dcore_U_sub_fifo_n534), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[31]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U229 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__32_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n560), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__32_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n538)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U228 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n20), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n85), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n536)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U227 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__32_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n536), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n537) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U226 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n59), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n538), .B(
        U_dfifo_U_dcore_U_sub_fifo_n537), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[32]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U225 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__0_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__0_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n463)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U224 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n52), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n117), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n461)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U223 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__0_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n461), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n462) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U222 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n83), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n463), .B(
        U_dfifo_U_dcore_U_sub_fifo_n462), .ZN(U_dfifo_U_dcore_m_sf_data_out[0]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U221 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n62), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n69), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n364) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U220 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n58), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n80), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n375) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U219 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n82), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n66), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n361) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U218 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n83), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n67), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n362) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U217 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n70), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n60), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n347) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U216 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n76), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n120), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n355) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U215 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n56), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n78), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n373) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U214 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n74), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n118), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n353) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U213 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n80), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n124), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n359) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U212 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n73), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n63), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n350) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U211 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n72), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n62), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n349) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U210 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n61), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n68), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n363) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U209 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n69), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n58), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n345) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U208 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n68), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n59), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n346) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U207 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n66), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n73), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n368) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U206 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n57), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n79), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n374) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U205 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n54), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n76), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n371) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U204 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n85), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n65), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n352) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U203 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n52), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n81), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n376) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U202 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n64), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n71), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n366) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U201 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n84), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n64), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n351) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U200 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n71), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n61), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n348) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U199 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n63), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n70), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n365) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U198 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n65), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n72), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n367) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U197 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n77), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n121), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n356) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U196 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n55), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n77), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n372) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U195 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n67), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n74), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n369) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U194 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n59), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n82), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n377) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U193 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n81), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n125), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n360) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U192 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n75), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n119), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n354) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U191 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n60), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n83), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n378) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U190 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n78), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n122), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n357) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U189 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n53), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n75), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n370) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U188 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n232), .A2(n79), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n123), .B2(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n358) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U187 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n65), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n150), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n333) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U186 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n74), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n136), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n319) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U185 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n81), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n143), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n326) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U184 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n77), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n139), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n322) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U183 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n76), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n138), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n321) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U182 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n66), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n151), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n334) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U181 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n63), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n148), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n331) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U180 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n85), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n135), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n318) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U179 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n64), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n149), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n332) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U178 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n83), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n145), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n328) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U177 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n79), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n141), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n324) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U176 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n84), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n134), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n317) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U175 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n67), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n152), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n335) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U174 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n71), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n131), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n314) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U173 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n62), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n147), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n330) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U172 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n53), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n153), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n336) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U171 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n82), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n144), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n327) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U170 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n75), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n137), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n320) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U169 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n54), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n154), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n337) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U168 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n68), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n129), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n312) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U167 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n55), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n155), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n338) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U166 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n70), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n130), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n313) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U165 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n80), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n142), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n325) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U164 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n56), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n156), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n339) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U163 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n69), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n128), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n311) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U162 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n72), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n132), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n315) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U161 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n78), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n140), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n323) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U160 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n57), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n157), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n340) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U159 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n61), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n146), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n329) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U158 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n73), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n133), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n316) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U157 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n58), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n158), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n341) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U156 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n59), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n160), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n343) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U155 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n60), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n161), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n344) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U154 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n231), .A2(n52), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n159), .B2(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n342) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U153 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__28_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__28_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n523)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U152 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n24), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n89), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n521)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U151 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__28_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n521), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n522) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U150 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n63), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n523), .B(
        U_dfifo_U_dcore_U_sub_fifo_n522), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[28]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U149 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__27_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__27_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n520)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U148 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n25), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n90), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n518)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U147 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__27_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n518), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n519) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U146 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n64), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n520), .B(
        U_dfifo_U_dcore_U_sub_fifo_n519), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[27]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U145 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__29_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__29_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n526)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U144 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n23), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n88), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n524)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U143 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__29_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n524), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n525) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U142 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n62), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n526), .B(
        U_dfifo_U_dcore_U_sub_fifo_n525), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[29]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U141 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__30_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__30_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n532)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U140 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n22), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n87), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n530)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U139 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__30_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n530), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n531) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U138 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n61), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n532), .B(
        U_dfifo_U_dcore_U_sub_fifo_n531), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[30]) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U137 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n56), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n224), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n441) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U136 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n68), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n197), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n414) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U135 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n69), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n196), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n413) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U134 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n71), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n199), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n416) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U133 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n59), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n228), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n445) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U132 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n73), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n201), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n418) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U131 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n72), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n200), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n417) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U130 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n53), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n221), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n438) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U129 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n70), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n198), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n415) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U128 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n60), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n229), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n446) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U127 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n57), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n225), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n442) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U126 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n52), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n227), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n444) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U125 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n55), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n223), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n440) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U124 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n54), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n222), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n439) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U123 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n58), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n226), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n443) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U122 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n63), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n182), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n399) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U121 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n66), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n185), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n402) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U120 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n56), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n190), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n407) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U119 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n61), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n180), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n397) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U118 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n55), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n189), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n406) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U117 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n60), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n195), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n412) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U116 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n54), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n188), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n405) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U115 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n62), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n181), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n398) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U114 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n64), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n183), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n400) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U113 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n57), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n191), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n408) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U112 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n65), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n184), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n401) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U111 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n58), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n192), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n409) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U110 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n53), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n187), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n404) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U109 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n67), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n186), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n403) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U108 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n59), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n194), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n411) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U107 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n52), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n193), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n410) );
  AOI22_X2 U_dfifo_U_dcore_U_sub_fifo_U106 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__1_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n230), .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__1_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n235), .ZN(U_dfifo_U_dcore_U_sub_fifo_n496)
         );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U105 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n51), .A2(U_dfifo_U_dcore_U_sub_fifo_n8), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n116), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n14), .ZN(U_dfifo_U_dcore_U_sub_fifo_n494)
         );
  AOI21_X2 U_dfifo_U_dcore_U_sub_fifo_U104 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__1_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n562), .A(U_dfifo_U_dcore_U_sub_fifo_n494), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n495) );
  OAI211_X2 U_dfifo_U_dcore_U_sub_fifo_U103 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n82), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n496), .B(
        U_dfifo_U_dcore_U_sub_fifo_n495), .ZN(U_dfifo_U_dcore_m_sf_data_out[1]) );
  NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U102 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n608), .A2(U_dfifo_U_dcore_U_sub_fifo_n18), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n607) );
  OAI22_X2 U_dfifo_U_dcore_U_sub_fifo_U101 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n607), .A2(U_dfifo_U_dcore_U_sub_fifo_n56), 
        .B1(U_dfifo_U_dcore_U_sub_fifo_n608), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n53), .ZN(U_dfifo_U_dcore_U_sub_fifo_n451)
         );
  OAI21_X2 U_dfifo_U_dcore_U_sub_fifo_U100 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_n607), .B2(U_dfifo_U_dcore_U_sub_fifo_n126), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n606), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n452) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U98 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n68), .B1(U_dfifo_U_dcore_U_sub_fifo_n85), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n6), .ZN(U_dfifo_U_dcore_U_sub_fifo_n278)
         );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U97 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n16), .A2(n69), .B1(U_dfifo_U_dcore_U_sub_fifo_n84), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n6), .ZN(U_dfifo_U_dcore_U_sub_fifo_n277)
         );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U96 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n69), .B1(U_dfifo_U_dcore_U_sub_fifo_n19), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n7), .ZN(U_dfifo_U_dcore_U_sub_fifo_n243)
         );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U95 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n15), .A2(n68), .B1(U_dfifo_U_dcore_U_sub_fifo_n20), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n7), .ZN(U_dfifo_U_dcore_U_sub_fifo_n244)
         );
  NAND2_X1 U_dfifo_U_dcore_U_sub_fifo_U94 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n57), .ZN(U_dfifo_U_dcore_U_sub_fifo_n567)
         );
  INV_X1 U_dfifo_U_dcore_U_sub_fifo_U93 ( .A(U_dfifo_U_dcore_U_sub_fifo_n609), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n608) );
  NAND3_X1 U_dfifo_U_dcore_U_sub_fifo_U92 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n609), .A2(U_dfifo_U_dcore_U_sub_fifo_n605), 
        .A3(U_dfifo_U_dcore_U_sub_fifo_n126), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n606) );
  NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U88 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n241), .A2(U_dfifo_U_dcore_U_sub_fifo_n17), .ZN(U_dfifo_U_dcore_m_sf_full) );
  NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U87 ( .A1(U_dfifo_U_dcore_n24), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n609), .ZN(U_dfifo_U_dcore_U_sub_fifo_n455)
         );
  NOR3_X2 U_dfifo_U_dcore_U_sub_fifo_U86 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n57), .A3(U_dfifo_U_dcore_U_sub_fifo_n604), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n16) );
  NOR3_X2 U_dfifo_U_dcore_U_sub_fifo_U85 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n57), .A3(U_dfifo_U_dcore_U_sub_fifo_n602), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n15) );
  INV_X4 U_dfifo_U_dcore_U_sub_fifo_U84 ( .A(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n234) );
  INV_X4 U_dfifo_U_dcore_U_sub_fifo_U83 ( .A(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n233) );
  NAND2_X2 U_dfifo_U_dcore_U_sub_fifo_U82 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n13), .A2(U_dfifo_U_dcore_U_sub_fifo_count_1_), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n241) );
  NAND2_X4 U_dfifo_U_dcore_U_sub_fifo_U81 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n460), .ZN(U_dfifo_U_dcore_U_sub_fifo_n53)
         );
  NAND2_X4 U_dfifo_U_dcore_U_sub_fifo_U80 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n18), .ZN(U_dfifo_U_dcore_U_sub_fifo_n14)
         );
  NAND2_X4 U_dfifo_U_dcore_U_sub_fifo_U79 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n8) );
  BUF_X4 U_dfifo_U_dcore_U_sub_fifo_U78 ( .A(U_dfifo_U_dcore_U_sub_fifo_n605), 
        .Z(U_dfifo_U_dcore_U_sub_fifo_n235) );
  BUF_X4 U_dfifo_U_dcore_U_sub_fifo_U77 ( .A(U_dfifo_U_dcore_U_sub_fifo_n560), 
        .Z(U_dfifo_U_dcore_U_sub_fifo_n230) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U76 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n120), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n508), .B(
        U_dfifo_U_dcore_U_sub_fifo_n507), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[23]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U75 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n121), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n505), .B(
        U_dfifo_U_dcore_U_sub_fifo_n504), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[22]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U74 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n122), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n502), .B(
        U_dfifo_U_dcore_U_sub_fifo_n501), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[21]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U73 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n123), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n499), .B(
        U_dfifo_U_dcore_U_sub_fifo_n498), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[20]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U72 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n75), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n559), .B(
        U_dfifo_U_dcore_U_sub_fifo_n558), .ZN(U_dfifo_U_dcore_m_sf_data_out[8]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U71 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n78), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n550), .B(
        U_dfifo_U_dcore_U_sub_fifo_n549), .ZN(U_dfifo_U_dcore_m_sf_data_out[5]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U70 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n77), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n553), .B(
        U_dfifo_U_dcore_U_sub_fifo_n552), .ZN(U_dfifo_U_dcore_m_sf_data_out[6]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U69 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n79), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n547), .B(
        U_dfifo_U_dcore_U_sub_fifo_n546), .ZN(U_dfifo_U_dcore_m_sf_data_out[4]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U68 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n76), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n556), .B(
        U_dfifo_U_dcore_U_sub_fifo_n555), .ZN(U_dfifo_U_dcore_m_sf_data_out[7]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U67 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n80), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n544), .B(
        U_dfifo_U_dcore_U_sub_fifo_n543), .ZN(U_dfifo_U_dcore_m_sf_data_out[3]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U66 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n74), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n564), .B(
        U_dfifo_U_dcore_U_sub_fifo_n563), .ZN(U_dfifo_U_dcore_m_sf_data_out[9]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U65 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n119), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n511), .B(
        U_dfifo_U_dcore_U_sub_fifo_n510), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[24]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U64 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n81), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n529), .B(
        U_dfifo_U_dcore_U_sub_fifo_n528), .ZN(U_dfifo_U_dcore_m_sf_data_out[2]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U63 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n118), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n514), .B(
        U_dfifo_U_dcore_U_sub_fifo_n513), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[25]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U62 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n125), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n490), .B(
        U_dfifo_U_dcore_U_sub_fifo_n489), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[18]) );
  OAI211_X1 U_dfifo_U_dcore_U_sub_fifo_U61 ( .C1(
        U_dfifo_U_dcore_U_sub_fifo_n124), .C2(U_dfifo_U_dcore_U_sub_fifo_n53), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n493), .B(
        U_dfifo_U_dcore_U_sub_fifo_n492), .ZN(
        U_dfifo_U_dcore_m_sf_data_out[19]) );
  NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U60 ( .A1(U_dfifo_U_dcore_n209), .A2(
        U_dfifo_U_dcore_m_sf_empty), .ZN(U_dfifo_U_dcore_U_sub_fifo_n609) );
  NOR2_X1 U_dfifo_U_dcore_U_sub_fifo_U59 ( .A1(U_dfifo_U_dcore_U_sub_fifo_n608), .A2(U_dfifo_U_dcore_U_sub_fifo_count_0_), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n565) );
  NOR2_X2 U_dfifo_U_dcore_U_sub_fifo_U58 ( .A1(U_dfifo_U_dcore_n208), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n455), .ZN(U_dfifo_U_dcore_U_sub_fifo_n458)
         );
  AOI21_X1 U_dfifo_U_dcore_U_sub_fifo_U57 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_n608), .B2(U_dfifo_U_dcore_U_sub_fifo_n18), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n607), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n453) );
  XOR2_X1 U_dfifo_U_dcore_U_sub_fifo_U56 ( .A(U_dfifo_U_dcore_U_sub_fifo_n459), 
        .B(U_dfifo_U_dcore_U_sub_fifo_n458), .Z(
        U_dfifo_U_dcore_U_sub_fifo_n454) );
  XNOR2_X1 U_dfifo_U_dcore_U_sub_fifo_U55 ( .A(
        U_dfifo_U_dcore_U_sub_fifo_count_1_), .B(
        U_dfifo_U_dcore_U_sub_fifo_n566), .ZN(U_dfifo_U_dcore_U_sub_fifo_n242)
         );
  INV_X4 U_dfifo_U_dcore_U_sub_fifo_U54 ( .A(U_dfifo_U_dcore_U_sub_fifo_n9), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n231) );
  INV_X4 U_dfifo_U_dcore_U_sub_fifo_U53 ( .A(U_dfifo_U_dcore_U_sub_fifo_n10), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n232) );
  OAI21_X1 U_dfifo_U_dcore_U_sub_fifo_U52 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_n603), .B2(U_dfifo_U_dcore_U_sub_fifo_n127), 
        .A(U_dfifo_U_dcore_U_sub_fifo_n10), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n447) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U51 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n84), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n202), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n419) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U50 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n75), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n205), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n422) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U49 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n74), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n204), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n421) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U48 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n85), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n203), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n420) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U47 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n77), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n207), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n424) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U46 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n78), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n208), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n425) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U45 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n79), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n209), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n426) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U44 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n80), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n210), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n427) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U43 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n76), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n206), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n423) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U42 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n81), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n211), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n428) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U41 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n82), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n212), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n429) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U40 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n83), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n213), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n430) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U39 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n61), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n214), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n431) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U38 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n62), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n215), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n432) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U37 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n63), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n216), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n433) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U36 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n64), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n217), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n434) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U35 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n65), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n218), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n435) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U34 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n66), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n219), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n436) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U33 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n234), .A2(n67), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n220), .B2(U_dfifo_U_dcore_U_sub_fifo_n12), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n437) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U32 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n69), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n162), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n379) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U31 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n68), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n163), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n380) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U30 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n70), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n164), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n381) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U29 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n71), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n165), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n382) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U28 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n72), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n166), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n383) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U27 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n73), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n167), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n384) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U26 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n84), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n168), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n385) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U25 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n85), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n169), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n386) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U24 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n74), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n170), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n387) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U23 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n75), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n171), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n388) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U22 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n76), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n172), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n389) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U21 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n77), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n173), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n390) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U20 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n78), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n174), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n391) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U19 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n79), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n175), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n392) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U18 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n80), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n176), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n393) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U17 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n81), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n177), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n394) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U16 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n82), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n178), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n395) );
  AOI22_X1 U_dfifo_U_dcore_U_sub_fifo_U15 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_n233), .A2(n83), .B1(
        U_dfifo_U_dcore_U_sub_fifo_n179), .B2(U_dfifo_U_dcore_U_sub_fifo_n11), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n396) );
  NOR3_X2 U_dfifo_U_dcore_U_sub_fifo_U14 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_count_2_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_count_0_), .A3(
        U_dfifo_U_dcore_U_sub_fifo_count_1_), .ZN(U_dfifo_U_dcore_m_sf_empty)
         );
  MUX2_X1 U_dfifo_U_dcore_U_sub_fifo_U13 ( .A(U_dfifo_U_dcore_U_sub_fifo_n609), 
        .B(U_dfifo_U_dcore_n209), .S(U_dfifo_U_dcore_U_sub_fifo_count_0_), .Z(
        U_dfifo_U_dcore_U_sub_fifo_n459) );
  AOI21_X1 U_dfifo_U_dcore_U_sub_fifo_U12 ( .B1(U_dfifo_U_dcore_n208), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n565), .A(U_dfifo_U_dcore_U_sub_fifo_n456), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n566) );
  INV_X4 U_dfifo_U_dcore_U_sub_fifo_U11 ( .A(U_dfifo_U_dcore_U_sub_fifo_n15), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n7) );
  INV_X4 U_dfifo_U_dcore_U_sub_fifo_U10 ( .A(U_dfifo_U_dcore_U_sub_fifo_n16), 
        .ZN(U_dfifo_U_dcore_U_sub_fifo_n6) );
  OAI221_X1 U_dfifo_U_dcore_U_sub_fifo_U8 ( .B1(
        U_dfifo_U_dcore_U_sub_fifo_count_2_), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n1), .C1(U_dfifo_U_dcore_U_sub_fifo_n17), 
        .C2(U_dfifo_U_dcore_U_sub_fifo_n5), .A(U_dfifo_U_dcore_n24), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n450) );
  AOI21_X1 U_dfifo_U_dcore_U_sub_fifo_U7 ( .B1(U_dfifo_U_dcore_n208), .B2(
        U_dfifo_U_dcore_U_sub_fifo_count_0_), .A(U_dfifo_U_dcore_U_sub_fifo_n4), .ZN(U_dfifo_U_dcore_U_sub_fifo_n5) );
  OAI22_X1 U_dfifo_U_dcore_U_sub_fifo_U6 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_count_1_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n3), .B1(U_dfifo_U_dcore_n208), .B2(
        U_dfifo_U_dcore_U_sub_fifo_n608), .ZN(U_dfifo_U_dcore_U_sub_fifo_n4)
         );
  INV_X1 U_dfifo_U_dcore_U_sub_fifo_U5 ( .A(U_dfifo_U_dcore_n209), .ZN(
        U_dfifo_U_dcore_U_sub_fifo_n3) );
  NAND2_X1 U_dfifo_U_dcore_U_sub_fifo_U3 ( .A1(
        U_dfifo_U_dcore_U_sub_fifo_count_1_), .A2(
        U_dfifo_U_dcore_U_sub_fifo_n456), .ZN(U_dfifo_U_dcore_U_sub_fifo_n1)
         );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_out_ptr_reg_0_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n453), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_0_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n18) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_out_ptr_reg_1_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n451), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_1_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n56) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_out_ptr_reg_2_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n452), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_out_ptr_2_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n126) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__5_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n373), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n78) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__6_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n372), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n77) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__7_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n371), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n76) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__8_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n370), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n75) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__9_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n369), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n74) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__10_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n368), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n73) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__11_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n367), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n72) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__12_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n366), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n71) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__13_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n365), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n70) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__14_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n364), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n69) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__15_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n363), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n68) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__16_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n362), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n67) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__17_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n361), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n66) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__18_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n360), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n125) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__19_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n359), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n124) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__20_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n358), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n123) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__21_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n357), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n122) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__22_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n356), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n121) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__23_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n355), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n120) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__24_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n354), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n119) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__25_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n353), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n118) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__26_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n352), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n65) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__27_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n351), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n64) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__28_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n350), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n63) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__29_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n349), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n62) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__30_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n348), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n61) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__31_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n347), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n60) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__32_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n346), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n59) );
  DFFR_X2 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__33_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n345), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n58) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_count_reg_1_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n242), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_count_1_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n54) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__33_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n243), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n19) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__32_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n244), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n20) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__31_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n245), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n21) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__30_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n246), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n22) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__29_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n247), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n23) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__28_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n248), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n24) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__27_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n249), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n25) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__26_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n250), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n26) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__25_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n251), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n27) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__24_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n252), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n28) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__23_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n253), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n29) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__22_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n254), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n30) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__21_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n255), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n31) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__20_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n256), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n32) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__19_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n257), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n33) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__18_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n258), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n34) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__17_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n259), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n35) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__16_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n260), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n36) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__15_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n261), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n37) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__14_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n262), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n38) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__13_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n263), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n39) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__12_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n264), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n40) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__11_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n265), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n41) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__10_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n266), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n42) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__9_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n267), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n43) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__8_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n268), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n44) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__7_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n269), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n45) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__6_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n270), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n46) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__5_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n271), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n47) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__4_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n272), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n48) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__3_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n273), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n49) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__2_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n274), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n50) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__1_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n275), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n51) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_5__0_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n276), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n52) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__33_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n277), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n84) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__32_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n278), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n85) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__31_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n279), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n86) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__30_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n280), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n87) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__29_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n281), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n88) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__28_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n282), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n89) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__27_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n283), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n90) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__26_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n284), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n91) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__25_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n285), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n92) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__24_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n286), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n93) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__23_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n287), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n94) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__22_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n288), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n95) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__21_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n289), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n96) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__20_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n290), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n97) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__19_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n291), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n98) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__18_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n292), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n99) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__17_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n293), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n100) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__16_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n294), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n101) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__15_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n295), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n102) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__14_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n296), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n103) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__13_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n297), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n104) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__12_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n298), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n105) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__11_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n299), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n106) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__10_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n300), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n107) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__9_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n301), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n108) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__8_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n302), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n109) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__7_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n303), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n110) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__6_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n304), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n111) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__5_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n305), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n112) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__4_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n306), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n113) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__3_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n307), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n114) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__2_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n308), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n115) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__1_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n309), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n116) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_4__0_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n310), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n117) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__33_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n311), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__33_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n128) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__32_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n312), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__32_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n129) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__31_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n313), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__31_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n130) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__30_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n314), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__30_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n131) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__29_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n315), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__29_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n132) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__28_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n316), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__28_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n133) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__27_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n317), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__27_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n134) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__26_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n318), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__26_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n135) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__25_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n319), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__25_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n136) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__24_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n320), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__24_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n137) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__23_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n321), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__23_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n138) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__22_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n322), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__22_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n139) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__21_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n323), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__21_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n140) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__20_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n324), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__20_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n141) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__19_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n325), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__19_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n142) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__18_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n326), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__18_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n143) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__17_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n327), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__17_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n144) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__16_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n328), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__16_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n145) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__15_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n329), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__15_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n146) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__14_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n330), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__14_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n147) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__13_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n331), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__13_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n148) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__12_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n332), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__12_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n149) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__11_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n333), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__11_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n150) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__10_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n334), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__10_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n151) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__9_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n335), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__9_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n152) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__8_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n336), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__8_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n153) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__7_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n337), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__7_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n154) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__6_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n338), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__6_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n155) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__5_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n339), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__5_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n156) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__4_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n340), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__4_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n157) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__3_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n341), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__3_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n158) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__2_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n342), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__2_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n159) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__1_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n343), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__1_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n160) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_0__0_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n344), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_0__0_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n161) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__4_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n374), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n79) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__3_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n375), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n80) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__2_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n376), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n81) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__1_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n377), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n82) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_1__0_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n378), .CK(hclk), .RN(hresetn), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n83) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__33_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n379), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__33_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n162) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__32_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n380), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__32_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n163) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__31_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n381), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__31_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n164) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__30_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n382), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__30_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n165) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__29_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n383), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__29_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n166) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__28_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n384), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__28_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n167) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__27_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n385), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__27_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n168) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__26_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n386), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__26_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n169) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__25_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n387), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__25_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n170) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__24_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n388), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__24_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n171) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__23_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n389), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__23_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n172) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__22_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n390), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__22_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n173) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__21_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n391), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__21_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n174) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__20_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n392), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__20_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n175) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__19_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n393), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__19_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n176) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__18_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n394), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__18_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n177) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__17_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n395), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__17_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n178) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__16_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n396), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__16_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n179) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__15_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n397), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__15_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n180) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__14_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n398), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__14_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n181) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__13_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n399), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__13_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n182) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__12_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n400), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__12_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n183) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__11_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n401), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__11_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n184) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__10_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n402), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__10_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n185) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__9_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n403), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__9_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n186) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__8_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n404), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__8_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n187) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__7_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n405), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__7_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n188) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__6_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n406), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__6_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n189) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__5_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n407), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__5_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n190) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__4_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n408), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__4_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n191) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__3_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n409), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__3_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n192) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__2_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n410), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__2_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n193) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__1_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n411), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__1_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n194) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_2__0_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n412), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_2__0_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n195) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__33_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n413), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__33_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n196) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__32_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n414), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__32_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n197) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__31_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n415), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__31_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n198) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__30_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n416), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__30_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n199) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__29_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n417), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__29_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n200) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__28_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n418), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__28_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n201) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__27_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n419), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__27_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n202) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__26_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n420), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__26_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n203) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__25_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n421), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__25_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n204) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__24_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n422), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__24_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n205) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__23_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n423), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__23_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n206) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__22_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n424), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__22_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n207) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__21_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n425), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__21_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n208) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__20_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n426), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__20_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n209) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__19_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n427), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__19_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n210) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__18_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n428), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__18_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n211) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__17_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n429), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__17_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n212) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__16_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n430), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__16_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n213) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__15_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n431), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__15_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n214) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__14_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n432), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__14_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n215) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__13_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n433), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__13_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n216) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__12_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n434), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__12_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n217) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__11_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n435), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__11_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n218) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__10_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n436), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__10_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n219) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__9_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n437), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__9_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n220) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__8_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n438), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__8_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n221) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__7_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n439), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__7_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n222) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__6_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n440), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__6_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n223) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__5_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n441), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__5_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n224) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__4_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n442), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__4_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n225) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__3_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n443), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__3_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n226) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__2_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n444), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__2_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n227) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__1_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n445), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__1_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n228) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_mem_reg_3__0_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n446), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_mem_3__0_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n229) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_in_ptr_reg_1_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n447), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_1_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n127) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_in_ptr_reg_2_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n448), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_2_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n57) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_in_ptr_reg_0_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n449), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_in_ptr_0_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n55) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_count_reg_2_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n450), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_count_2_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n17) );
  DFFR_X1 U_dfifo_U_dcore_U_sub_fifo_count_reg_0_ ( .D(
        U_dfifo_U_dcore_U_sub_fifo_n454), .CK(hclk), .RN(hresetn), .Q(
        U_dfifo_U_dcore_U_sub_fifo_count_0_), .QN(
        U_dfifo_U_dcore_U_sub_fifo_n13) );
  NOR2_X1 U3 ( .A1(U_ctl_n400), .A2(U_ctl_n288), .ZN(n10) );
  AOI22_X1 U4 ( .A1(U_afifo_n54), .A2(U_afifo_f_data2_12_), .B1(U_afifo_n140), 
        .B2(n10), .ZN(n11) );
  INV_X1 U5 ( .A(n11), .ZN(U_afifo_m_data_in[12]) );
  AOI22_X1 U6 ( .A1(haddr[6]), .A2(U_afifo_n93), .B1(U_afifo_f_data2_16_), 
        .B2(U_afifo_n54), .ZN(n12) );
  INV_X1 U7 ( .A(n12), .ZN(U_afifo_m_data_in[16]) );
  AOI22_X1 U8 ( .A1(haddr[31]), .A2(U_afifo_n99), .B1(U_afifo_f_data2_41_), 
        .B2(U_afifo_n54), .ZN(n13) );
  INV_X1 U9 ( .A(n13), .ZN(U_afifo_m_data_in[41]) );
  AOI22_X1 U10 ( .A1(haddr[26]), .A2(U_afifo_n98), .B1(U_afifo_f_data2_36_), 
        .B2(U_afifo_n54), .ZN(n14) );
  INV_X1 U11 ( .A(n14), .ZN(U_afifo_m_data_in[36]) );
  AOI22_X1 U12 ( .A1(haddr[18]), .A2(U_afifo_n147), .B1(U_afifo_f_data2_28_), 
        .B2(U_afifo_n54), .ZN(n15) );
  INV_X1 U13 ( .A(n15), .ZN(U_afifo_m_data_in[28]) );
  AOI22_X1 U14 ( .A1(haddr[7]), .A2(U_afifo_n93), .B1(U_afifo_f_data2_17_), 
        .B2(U_afifo_n54), .ZN(n16) );
  INV_X1 U15 ( .A(n16), .ZN(U_afifo_m_data_in[17]) );
  AOI22_X1 U16 ( .A1(haddr[30]), .A2(U_afifo_n140), .B1(U_afifo_f_data2_40_), 
        .B2(U_afifo_n54), .ZN(n17) );
  INV_X1 U17 ( .A(n17), .ZN(U_afifo_m_data_in[40]) );
  AOI22_X1 U18 ( .A1(haddr[25]), .A2(U_afifo_n98), .B1(U_afifo_f_data2_35_), 
        .B2(U_afifo_n54), .ZN(n18) );
  INV_X1 U19 ( .A(n18), .ZN(U_afifo_m_data_in[35]) );
  AOI22_X1 U20 ( .A1(haddr[21]), .A2(U_afifo_n99), .B1(U_afifo_f_data2_31_), 
        .B2(U_afifo_n54), .ZN(n19) );
  INV_X1 U21 ( .A(n19), .ZN(U_afifo_m_data_in[31]) );
  AOI22_X1 U22 ( .A1(haddr[17]), .A2(U_afifo_n147), .B1(U_afifo_f_data2_27_), 
        .B2(U_afifo_n54), .ZN(n20) );
  INV_X1 U23 ( .A(n20), .ZN(U_afifo_m_data_in[27]) );
  INV_X1 U24 ( .A(U_ctl_n308), .ZN(n21) );
  NOR3_X1 U25 ( .A1(U_ctl_fr_prv_1wrap), .A2(U_ctl_n97), .A3(n21), .ZN(n22) );
  NOR4_X1 U26 ( .A1(miu_pop_n), .A2(hiu_rw), .A3(n22), .A4(m_df_push_n), .ZN(
        n23) );
  OAI221_X1 U27 ( .B1(U_dfifo_m_empty), .B2(U_dfifo_n5), .C1(U_dfifo_m_empty), 
        .C2(U_dfifo_m_aempty), .A(n23), .ZN(U_ctl_n304) );
  AOI22_X1 U28 ( .A1(haddr[29]), .A2(U_afifo_n93), .B1(U_afifo_f_data2_39_), 
        .B2(U_afifo_n54), .ZN(n24) );
  INV_X1 U29 ( .A(n24), .ZN(U_afifo_m_data_in[39]) );
  AOI22_X1 U30 ( .A1(haddr[24]), .A2(U_afifo_n98), .B1(U_afifo_f_data2_34_), 
        .B2(U_afifo_n54), .ZN(n25) );
  INV_X1 U31 ( .A(n25), .ZN(U_afifo_m_data_in[34]) );
  AOI22_X1 U32 ( .A1(haddr[23]), .A2(U_afifo_n140), .B1(U_afifo_f_data2_33_), 
        .B2(U_afifo_n54), .ZN(n26) );
  INV_X1 U33 ( .A(n26), .ZN(U_afifo_m_data_in[33]) );
  AOI22_X1 U34 ( .A1(haddr[16]), .A2(U_afifo_n147), .B1(U_afifo_f_data2_26_), 
        .B2(U_afifo_n54), .ZN(n27) );
  INV_X1 U35 ( .A(n27), .ZN(U_afifo_m_data_in[26]) );
  AOI22_X1 U36 ( .A1(haddr[14]), .A2(U_afifo_n99), .B1(U_afifo_f_data2_24_), 
        .B2(U_afifo_n54), .ZN(n28) );
  INV_X1 U37 ( .A(n28), .ZN(U_afifo_m_data_in[24]) );
  OAI22_X1 U38 ( .A1(U_afifo_U_acore_n1), .A2(U_afifo_U_acore_n8), .B1(
        U_afifo_U_acore_n35), .B2(U_afifo_U_acore_n32), .ZN(hiu_burst_size[5])
         );
  AOI22_X1 U39 ( .A1(haddr[27]), .A2(U_afifo_n93), .B1(U_afifo_f_data2_37_), 
        .B2(U_afifo_n54), .ZN(n29) );
  INV_X1 U40 ( .A(n29), .ZN(U_afifo_m_data_in[37]) );
  AOI22_X1 U41 ( .A1(haddr[20]), .A2(U_afifo_n140), .B1(U_afifo_f_data2_30_), 
        .B2(U_afifo_n54), .ZN(n30) );
  INV_X1 U42 ( .A(n30), .ZN(U_afifo_m_data_in[30]) );
  AOI22_X1 U43 ( .A1(haddr[19]), .A2(U_afifo_n98), .B1(U_afifo_f_data2_29_), 
        .B2(U_afifo_n54), .ZN(n31) );
  INV_X1 U44 ( .A(n31), .ZN(U_afifo_m_data_in[29]) );
  AOI22_X1 U45 ( .A1(haddr[10]), .A2(U_afifo_n147), .B1(U_afifo_f_data2_20_), 
        .B2(U_afifo_n54), .ZN(n32) );
  INV_X1 U46 ( .A(n32), .ZN(U_afifo_m_data_in[20]) );
  AOI22_X1 U47 ( .A1(m_af_data1_in_2_), .A2(U_afifo_n99), .B1(
        U_afifo_f_data2_2_), .B2(U_afifo_n54), .ZN(n33) );
  INV_X1 U48 ( .A(n33), .ZN(U_afifo_m_data_in[2]) );
  INV_X1 U49 ( .A(U_rbuf_n123), .ZN(n34) );
  AOI21_X1 U50 ( .B1(U_rbuf_n34), .B2(n34), .A(miu_push_n), .ZN(U_rbuf_n161)
         );
  OAI22_X1 U51 ( .A1(U_afifo_U_acore_n1), .A2(U_afifo_U_acore_n4), .B1(
        U_afifo_U_acore_n35), .B2(U_afifo_U_acore_n181), .ZN(hiu_burst_size[0]) );
  INV_X1 U52 ( .A(U_ctl_n288), .ZN(n35) );
  INV_X1 U53 ( .A(U_ctl_n189), .ZN(n36) );
  AOI22_X1 U54 ( .A1(U_ctl_n189), .A2(U_ctl_f_amba_bsz2[0]), .B1(n35), .B2(n36), .ZN(U_ctl_n163) );
  AOI22_X1 U55 ( .A1(haddr[15]), .A2(U_afifo_n93), .B1(U_afifo_f_data2_25_), 
        .B2(U_afifo_n54), .ZN(n37) );
  INV_X1 U56 ( .A(n37), .ZN(U_afifo_m_data_in[25]) );
  AOI22_X1 U57 ( .A1(haddr[13]), .A2(U_afifo_n99), .B1(U_afifo_f_data2_23_), 
        .B2(U_afifo_n54), .ZN(n38) );
  INV_X1 U58 ( .A(n38), .ZN(U_afifo_m_data_in[23]) );
  AOI22_X1 U59 ( .A1(haddr[12]), .A2(U_afifo_n98), .B1(U_afifo_f_data2_22_), 
        .B2(U_afifo_n54), .ZN(n39) );
  INV_X1 U60 ( .A(n39), .ZN(U_afifo_m_data_in[22]) );
  AOI22_X1 U61 ( .A1(haddr[11]), .A2(U_afifo_n140), .B1(U_afifo_f_data2_21_), 
        .B2(U_afifo_n54), .ZN(n40) );
  INV_X1 U62 ( .A(n40), .ZN(U_afifo_m_data_in[21]) );
  AOI22_X1 U63 ( .A1(haddr[9]), .A2(U_afifo_n147), .B1(U_afifo_f_data2_19_), 
        .B2(U_afifo_n54), .ZN(n41) );
  INV_X1 U64 ( .A(n41), .ZN(U_afifo_m_data_in[19]) );
  INV_X1 U65 ( .A(U_ctl_fd_amba_bcnt_1_), .ZN(n42) );
  NOR4_X1 U66 ( .A1(U_ctl_n338), .A2(U_ctl_n382), .A3(U_ctl_fd_amba_bcnt_0_), 
        .A4(n42), .ZN(n43) );
  AOI211_X1 U67 ( .C1(U_ctl_n395), .C2(U_ctl_n145), .A(n43), .B(U_ctl_n323), 
        .ZN(U_ctl_n118) );
  NOR3_X1 U68 ( .A1(U_ctl_n381), .A2(U_ctl_n238), .A3(U_ctl_n237), .ZN(n44) );
  NAND2_X1 U69 ( .A1(n47), .A2(haddr[7]), .ZN(n45) );
  OAI22_X1 U70 ( .A1(n44), .A2(n45), .B1(U_afifo_n164), .B2(n47), .ZN(
        U_afifo_n21) );
  NAND3_X1 U71 ( .A1(n47), .A2(U_ctl_n92), .A3(U_ctl_n150), .ZN(n46) );
  OAI21_X1 U72 ( .B1(U_afifo_n158), .B2(n47), .A(n46), .ZN(U_afifo_n12) );
  INV_X2 U73 ( .A(U_afifo_n15), .ZN(U_afifo_m_data_in[48]) );
  INV_X2 U74 ( .A(U_ctl_n68), .ZN(U_ctl_n67) );
  NOR2_X2 U75 ( .A1(n8), .A2(U_ctl_n190), .ZN(U_ctl_n68) );
  INV_X2 U76 ( .A(miu_data[0]), .ZN(U_rbuf_n181) );
  INV_X2 U77 ( .A(miu_data[1]), .ZN(U_rbuf_n182) );
  INV_X2 U78 ( .A(miu_data[3]), .ZN(U_rbuf_n184) );
  INV_X2 U79 ( .A(miu_data[5]), .ZN(U_rbuf_n186) );
  INV_X2 U80 ( .A(miu_data[6]), .ZN(U_rbuf_n187) );
  INV_X2 U81 ( .A(miu_data[7]), .ZN(U_rbuf_n188) );
  INV_X2 U82 ( .A(miu_data[9]), .ZN(U_rbuf_n190) );
  INV_X2 U83 ( .A(miu_data[10]), .ZN(U_rbuf_n191) );
  INV_X2 U84 ( .A(miu_data[12]), .ZN(U_rbuf_n193) );
  INV_X8 U85 ( .A(n47), .ZN(U_afifo_n176) );
  INV_X8 U86 ( .A(n47), .ZN(U_afifo_n174) );
  AND2_X4 U87 ( .A1(m_af_data1_in_3_), .A2(hready), .ZN(n47) );
  OR2_X2 U88 ( .A1(U_ctl_n90), .A2(U_ctl_n298), .ZN(n49) );
  AND2_X2 U89 ( .A1(U_rbuf_n145), .A2(U_rbuf_f_top_data_13_), .ZN(n50) );
  OR2_X4 U90 ( .A1(U_ctl_n332), .A2(U_ctl_n278), .ZN(n51) );
endmodule


module DW_memctl_miu ( hclk, hclk_2x, hresetn, scan_mode, hiu_mem_req, 
        hiu_reg_req, hiu_rw, hiu_burst_size, hiu_wrapped_burst, hiu_terminate, 
        hiu_addr, hiu_haddr, hiu_hsize, hiu_wr_data, s_rd_data, miu_burst_done, 
        miu_pop_n, miu_push_n, miu_col_addr_width, miu_data_width, m_addr, 
        s_addr, s_bank_addr, s_ras_n, s_cas_n, s_sel_n, s_cke, sf_cke, s_we_n, 
        s_wr_data, s_dqm, s_dout_valid, s_rd_ready, s_rd_start, s_rd_pop, 
        s_rd_end, s_rd_dqs_mask, s_cas_latency, s_read_pipe, sf_cas_latency, 
        s_sa, s_scl, s_dqs, s_rp_n, s_sda_out, s_sda_in, s_sda_oe_n, sm_addr, 
        sm_oe_n, sm_we_n, sm_bs_n, sm_dout_valid, sm_rp_n, sm_wp_n, sm_adv_n, 
        sm_rd_data, sm_wr_data, remap, sm_clken, sm_ready, sm_data_width_set0, 
        sm_access, m_wr_data, m_dout_valid, m_precharge_bit, s_ebi_req, 
        s_ebi_gnt, sm_ebi_req, sm_ebi_gnt, power_down, sf_power_down, 
        sm_power_down, clear_sr_dp, sf_clear_dp, big_endian, miu_rd_data_out, 
        gpi, gpo, debug_ad_bank_addr, debug_ad_row_addr, debug_ad_sf_bank_addr, 
        debug_ad_sf_row_addr, debug_ad_sf_col_addr, debug_sm_burst_done, 
        debug_sm_pop_n, debug_sm_push_n, debug_smc_cs, debug_ref_req, 
        debug_ad_col_addr_15_, debug_ad_col_addr_14_, debug_ad_col_addr_11_, 
        debug_ad_col_addr_10_, debug_ad_col_addr_9_, debug_ad_col_addr_8_, 
        debug_ad_col_addr_7_, debug_ad_col_addr_6_, debug_ad_col_addr_5_, 
        debug_ad_col_addr_4_, debug_ad_col_addr_3_, debug_ad_col_addr_2_, 
        debug_ad_col_addr_1_, debug_ad_col_addr_0_, 
        debug_ad_col_addr_13__BAR_BAR, debug_ad_col_addr_12__BAR_BAR );
  input [5:0] hiu_burst_size;
  input [31:0] hiu_addr;
  input [3:0] hiu_haddr;
  input [2:0] hiu_hsize;
  input [31:0] hiu_wr_data;
  input [31:0] s_rd_data;
  output [3:0] miu_col_addr_width;
  output [1:0] miu_data_width;
  output [15:0] m_addr;
  output [15:0] s_addr;
  output [1:0] s_bank_addr;
  output [0:0] s_sel_n;
  output [15:0] s_wr_data;
  output [1:0] s_dqm;
  output [1:0] s_dout_valid;
  output [2:0] s_cas_latency;
  output [2:0] s_read_pipe;
  output [2:0] sf_cas_latency;
  output [2:0] s_sa;
  output [1:0] s_dqs;
  output [22:0] sm_addr;
  output [3:0] sm_bs_n;
  output [3:0] sm_dout_valid;
  output [2:0] sm_wp_n;
  input [31:0] sm_rd_data;
  output [31:0] sm_wr_data;
  input [2:0] sm_data_width_set0;
  output [15:0] m_wr_data;
  output [1:0] m_dout_valid;
  output [31:0] miu_rd_data_out;
  input [7:0] gpi;
  output [7:0] gpo;
  output [1:0] debug_ad_bank_addr;
  output [15:0] debug_ad_row_addr;
  output [1:0] debug_ad_sf_bank_addr;
  output [15:0] debug_ad_sf_row_addr;
  output [15:0] debug_ad_sf_col_addr;
  output [3:0] debug_smc_cs;
  input hclk, hclk_2x, hresetn, scan_mode, hiu_mem_req, hiu_reg_req, hiu_rw,
         hiu_wrapped_burst, hiu_terminate, s_rd_ready, s_sda_in, remap,
         sm_clken, sm_ready, s_ebi_gnt, sm_ebi_gnt, power_down, sf_power_down,
         sm_power_down, clear_sr_dp, sf_clear_dp, big_endian;
  output miu_burst_done, miu_pop_n, miu_push_n, s_ras_n, s_cas_n, s_cke,
         sf_cke, s_we_n, s_rd_start, s_rd_pop, s_rd_end, s_rd_dqs_mask, s_scl,
         s_rp_n, s_sda_out, s_sda_oe_n, sm_oe_n, sm_we_n, sm_rp_n, sm_adv_n,
         sm_access, m_precharge_bit, s_ebi_req, sm_ebi_req,
         debug_sm_burst_done, debug_sm_pop_n, debug_sm_push_n, debug_ref_req,
         debug_ad_col_addr_15_, debug_ad_col_addr_14_, debug_ad_col_addr_11_,
         debug_ad_col_addr_10_, debug_ad_col_addr_9_, debug_ad_col_addr_8_,
         debug_ad_col_addr_7_, debug_ad_col_addr_6_, debug_ad_col_addr_5_,
         debug_ad_col_addr_4_, debug_ad_col_addr_3_, debug_ad_col_addr_2_,
         debug_ad_col_addr_1_, debug_ad_col_addr_0_,
         debug_ad_col_addr_13__BAR_BAR, debug_ad_col_addr_12__BAR_BAR;
  wire   n27, n44, debug_ad_col_addr_13_, debug_ad_col_addr_12_,
         ad_static_mem_req, cr_do_self_ref_rp, ctl_burst_done, ctl_pop_n,
         cr_pop_n, dmc_pop_n, ctl_push_n, cr_push_reg_n, dmc_push_n,
         sdram_req_i, ctl_auto_ref_en, ctl_ext_mode_reg_done, ctl_ref_ack,
         cr_push_n, ad_sdram_type_0_, ctl_chip_select_0_, pre_amble,
         pre_rd_dqs_mask, ad_sdram_chip_select_0_, cr_s_ready_valid,
         cr_do_initialize, cr_do_power_down, cr_mode_reg_update,
         cr_exn_mode_reg_update, cr_delayed_precharge, cr_ref_all_before_sr,
         cr_ref_all_after_sr, ctl_init_done, ctl_mode_reg_done,
         ctl_sd_in_sf_mode, cr_s_data_width_early_0_, N28, n1, n2, n3, n4, n5,
         n6, n7, n14, n16, n17, n18, n19, n21, U_dsdc_n2085, U_dsdc_n2084,
         U_dsdc_n2083, U_dsdc_n2082, U_dsdc_n2081, U_dsdc_n2080, U_dsdc_n2079,
         U_dsdc_n2078, U_dsdc_n2077, U_dsdc_n2076, U_dsdc_n2075, U_dsdc_n2074,
         U_dsdc_n2073, U_dsdc_n2072, U_dsdc_n2071, U_dsdc_n2070, U_dsdc_n2069,
         U_dsdc_n2068, U_dsdc_n2067, U_dsdc_n2066, U_dsdc_n2065, U_dsdc_n2064,
         U_dsdc_n2063, U_dsdc_n2062, U_dsdc_n2061, U_dsdc_n2060, U_dsdc_n2059,
         U_dsdc_n2058, U_dsdc_n2057, U_dsdc_n2056, U_dsdc_n2055, U_dsdc_n2054,
         U_dsdc_n2053, U_dsdc_n2052, U_dsdc_n2051, U_dsdc_n2050, U_dsdc_n2049,
         U_dsdc_n2048, U_dsdc_n2047, U_dsdc_n2046, U_dsdc_n2045, U_dsdc_n2044,
         U_dsdc_n2043, U_dsdc_n2042, U_dsdc_n2041, U_dsdc_n2040, U_dsdc_n2039,
         U_dsdc_n2038, U_dsdc_n2037, U_dsdc_n2036, U_dsdc_n2035, U_dsdc_n2034,
         U_dsdc_n2033, U_dsdc_n2032, U_dsdc_n2031, U_dsdc_n2030, U_dsdc_n2029,
         U_dsdc_n2028, U_dsdc_n2027, U_dsdc_n2026, U_dsdc_n2025, U_dsdc_n2024,
         U_dsdc_n2023, U_dsdc_n2022, U_dsdc_n2021, U_dsdc_n2020, U_dsdc_n2019,
         U_dsdc_n2018, U_dsdc_n2017, U_dsdc_n2016, U_dsdc_n2015, U_dsdc_n2014,
         U_dsdc_n2013, U_dsdc_n2012, U_dsdc_n2010, U_dsdc_n2009, U_dsdc_n2008,
         U_dsdc_n2007, U_dsdc_n2006, U_dsdc_n2005, U_dsdc_n2003, U_dsdc_n2001,
         U_dsdc_n1999, U_dsdc_n1997, U_dsdc_n1995, U_dsdc_n1994, U_dsdc_n1993,
         U_dsdc_n1992, U_dsdc_n1991, U_dsdc_n1990, U_dsdc_n1989, U_dsdc_n1988,
         U_dsdc_n1987, U_dsdc_n1986, U_dsdc_n1985, U_dsdc_n1984, U_dsdc_n1983,
         U_dsdc_n1982, U_dsdc_n1981, U_dsdc_n1980, U_dsdc_n1979, U_dsdc_n1978,
         U_dsdc_n1977, U_dsdc_n1976, U_dsdc_n1975, U_dsdc_n1974, U_dsdc_n1973,
         U_dsdc_n1972, U_dsdc_n1971, U_dsdc_n1970, U_dsdc_n1969, U_dsdc_n1968,
         U_dsdc_n1967, U_dsdc_n1966, U_dsdc_n1965, U_dsdc_n1964, U_dsdc_n1963,
         U_dsdc_n1962, U_dsdc_n1961, U_dsdc_n1960, U_dsdc_n1959, U_dsdc_n1958,
         U_dsdc_n1957, U_dsdc_n1956, U_dsdc_n1954, U_dsdc_n1953, U_dsdc_n1951,
         U_dsdc_n1948, U_dsdc_n1947, U_dsdc_n1946, U_dsdc_n1945, U_dsdc_n1944,
         U_dsdc_n1943, U_dsdc_n1942, U_dsdc_n1941, U_dsdc_n1940, U_dsdc_n1939,
         U_dsdc_n1938, U_dsdc_n1937, U_dsdc_n1936, U_dsdc_n1935, U_dsdc_n1934,
         U_dsdc_n1933, U_dsdc_n1932, U_dsdc_n1931, U_dsdc_n1930, U_dsdc_n1929,
         U_dsdc_n1928, U_dsdc_n1927, U_dsdc_n1926, U_dsdc_n1925, U_dsdc_n1924,
         U_dsdc_n1923, U_dsdc_n1922, U_dsdc_n1921, U_dsdc_n1920, U_dsdc_n1919,
         U_dsdc_n1918, U_dsdc_n1917, U_dsdc_n1916, U_dsdc_n1915, U_dsdc_n1914,
         U_dsdc_n1913, U_dsdc_n1912, U_dsdc_n1911, U_dsdc_n1910, U_dsdc_n1909,
         U_dsdc_n1908, U_dsdc_n1907, U_dsdc_n1906, U_dsdc_n1905, U_dsdc_n1904,
         U_dsdc_n1903, U_dsdc_n1902, U_dsdc_n1901, U_dsdc_n1900, U_dsdc_n1899,
         U_dsdc_n1898, U_dsdc_n1897, U_dsdc_n1896, U_dsdc_n1895, U_dsdc_n1894,
         U_dsdc_n1893, U_dsdc_n1892, U_dsdc_n1891, U_dsdc_n1890, U_dsdc_n1889,
         U_dsdc_n1888, U_dsdc_n1887, U_dsdc_n1886, U_dsdc_n1885, U_dsdc_n1884,
         U_dsdc_n1883, U_dsdc_n1882, U_dsdc_n1881, U_dsdc_n1880, U_dsdc_n1879,
         U_dsdc_n1878, U_dsdc_n1877, U_dsdc_n1876, U_dsdc_n1875, U_dsdc_n1874,
         U_dsdc_n1872, U_dsdc_n1871, U_dsdc_n1870, U_dsdc_n1869, U_dsdc_n1868,
         U_dsdc_n1867, U_dsdc_n1866, U_dsdc_n1865, U_dsdc_n1864, U_dsdc_n1863,
         U_dsdc_n1862, U_dsdc_n1861, U_dsdc_n1860, U_dsdc_n1859, U_dsdc_n1858,
         U_dsdc_n1857, U_dsdc_n1856, U_dsdc_n1855, U_dsdc_n1854, U_dsdc_n1853,
         U_dsdc_n1852, U_dsdc_n1851, U_dsdc_n1850, U_dsdc_n1849, U_dsdc_n1848,
         U_dsdc_n1847, U_dsdc_n1846, U_dsdc_n1844, U_dsdc_n1843, U_dsdc_n1842,
         U_dsdc_n1841, U_dsdc_n1840, U_dsdc_n1839, U_dsdc_n1837, U_dsdc_n1836,
         U_dsdc_n1834, U_dsdc_n1833, U_dsdc_n1832, U_dsdc_n1831, U_dsdc_n1830,
         U_dsdc_n1829, U_dsdc_n1828, U_dsdc_n1827, U_dsdc_n1826, U_dsdc_n1825,
         U_dsdc_n1824, U_dsdc_n1823, U_dsdc_n1822, U_dsdc_n1821, U_dsdc_n1820,
         U_dsdc_n1819, U_dsdc_n1818, U_dsdc_n1817, U_dsdc_n1816, U_dsdc_n1815,
         U_dsdc_n1814, U_dsdc_n1813, U_dsdc_n1812, U_dsdc_n1811, U_dsdc_n1810,
         U_dsdc_n1809, U_dsdc_n1808, U_dsdc_n1807, U_dsdc_n1806, U_dsdc_n1805,
         U_dsdc_n1804, U_dsdc_n1803, U_dsdc_n1802, U_dsdc_n1801, U_dsdc_n1800,
         U_dsdc_n1799, U_dsdc_n1798, U_dsdc_n1797, U_dsdc_n1796, U_dsdc_n1795,
         U_dsdc_n1794, U_dsdc_n1793, U_dsdc_n1792, U_dsdc_n1791, U_dsdc_n1790,
         U_dsdc_n1789, U_dsdc_n1788, U_dsdc_n1787, U_dsdc_n1786, U_dsdc_n1785,
         U_dsdc_n1784, U_dsdc_n1783, U_dsdc_n1782, U_dsdc_n1781, U_dsdc_n1780,
         U_dsdc_n1779, U_dsdc_n1778, U_dsdc_n1777, U_dsdc_n1776, U_dsdc_n1775,
         U_dsdc_n1774, U_dsdc_n1773, U_dsdc_n1772, U_dsdc_n1771, U_dsdc_n1770,
         U_dsdc_n1769, U_dsdc_n1768, U_dsdc_n1767, U_dsdc_n1766, U_dsdc_n1765,
         U_dsdc_n1764, U_dsdc_n1763, U_dsdc_n1762, U_dsdc_n1761, U_dsdc_n1760,
         U_dsdc_n1759, U_dsdc_n1758, U_dsdc_n1757, U_dsdc_n1756, U_dsdc_n1755,
         U_dsdc_n1754, U_dsdc_n1753, U_dsdc_n1752, U_dsdc_n1751, U_dsdc_n1750,
         U_dsdc_n1749, U_dsdc_n1748, U_dsdc_n1747, U_dsdc_n1746, U_dsdc_n1745,
         U_dsdc_n1744, U_dsdc_n1743, U_dsdc_n1742, U_dsdc_n1741, U_dsdc_n1740,
         U_dsdc_n1739, U_dsdc_n1738, U_dsdc_n1737, U_dsdc_n1736, U_dsdc_n1735,
         U_dsdc_n1734, U_dsdc_n1733, U_dsdc_n1732, U_dsdc_n1731, U_dsdc_n1730,
         U_dsdc_n1729, U_dsdc_n1728, U_dsdc_n1727, U_dsdc_n1726, U_dsdc_n1725,
         U_dsdc_n1724, U_dsdc_n1723, U_dsdc_n1722, U_dsdc_n1721, U_dsdc_n1720,
         U_dsdc_n1719, U_dsdc_n1718, U_dsdc_n1717, U_dsdc_n1716, U_dsdc_n1715,
         U_dsdc_n1714, U_dsdc_n1713, U_dsdc_n1712, U_dsdc_n1711, U_dsdc_n1710,
         U_dsdc_n1709, U_dsdc_n1708, U_dsdc_n1707, U_dsdc_n1706, U_dsdc_n1705,
         U_dsdc_n1704, U_dsdc_n1703, U_dsdc_n1702, U_dsdc_n1701, U_dsdc_n1700,
         U_dsdc_n1699, U_dsdc_n1698, U_dsdc_n1697, U_dsdc_n1696, U_dsdc_n1695,
         U_dsdc_n1694, U_dsdc_n1693, U_dsdc_n1692, U_dsdc_n1691, U_dsdc_n1690,
         U_dsdc_n1689, U_dsdc_n1688, U_dsdc_n1687, U_dsdc_n1686, U_dsdc_n1685,
         U_dsdc_n1684, U_dsdc_n1683, U_dsdc_n1682, U_dsdc_n1681, U_dsdc_n1680,
         U_dsdc_n1679, U_dsdc_n1678, U_dsdc_n1677, U_dsdc_n1676, U_dsdc_n1675,
         U_dsdc_n1674, U_dsdc_n1673, U_dsdc_n1672, U_dsdc_n1671, U_dsdc_n1670,
         U_dsdc_n1669, U_dsdc_n1668, U_dsdc_n1667, U_dsdc_n1666, U_dsdc_n1662,
         U_dsdc_n1661, U_dsdc_n1660, U_dsdc_n1659, U_dsdc_n1658, U_dsdc_n1657,
         U_dsdc_n1656, U_dsdc_n1655, U_dsdc_n1654, U_dsdc_n1653, U_dsdc_n1652,
         U_dsdc_n1651, U_dsdc_n1650, U_dsdc_n1649, U_dsdc_n1648, U_dsdc_n1647,
         U_dsdc_n1646, U_dsdc_n1645, U_dsdc_n1644, U_dsdc_n1643, U_dsdc_n1642,
         U_dsdc_n1641, U_dsdc_n1640, U_dsdc_n1639, U_dsdc_n1638, U_dsdc_n1637,
         U_dsdc_n1636, U_dsdc_n1635, U_dsdc_n1634, U_dsdc_n1633, U_dsdc_n1632,
         U_dsdc_n1631, U_dsdc_n1630, U_dsdc_n1629, U_dsdc_n1628, U_dsdc_n1627,
         U_dsdc_n1626, U_dsdc_n1625, U_dsdc_n1624, U_dsdc_n1623, U_dsdc_n1622,
         U_dsdc_n1621, U_dsdc_n1620, U_dsdc_n1619, U_dsdc_n1618, U_dsdc_n1617,
         U_dsdc_n1616, U_dsdc_n1615, U_dsdc_n1614, U_dsdc_n1612, U_dsdc_n1611,
         U_dsdc_n1610, U_dsdc_n1609, U_dsdc_n1608, U_dsdc_n1606, U_dsdc_n1605,
         U_dsdc_n1604, U_dsdc_n1603, U_dsdc_n1602, U_dsdc_n1601, U_dsdc_n1600,
         U_dsdc_n1598, U_dsdc_n1597, U_dsdc_n1596, U_dsdc_n1594, U_dsdc_n1593,
         U_dsdc_n1592, U_dsdc_n1591, U_dsdc_n1590, U_dsdc_n1589, U_dsdc_n1588,
         U_dsdc_n1587, U_dsdc_n1586, U_dsdc_n1585, U_dsdc_n1584, U_dsdc_n1583,
         U_dsdc_n1582, U_dsdc_n1581, U_dsdc_n1580, U_dsdc_n1579, U_dsdc_n1578,
         U_dsdc_n1577, U_dsdc_n1576, U_dsdc_n1575, U_dsdc_n1574, U_dsdc_n1573,
         U_dsdc_n1572, U_dsdc_n1571, U_dsdc_n1570, U_dsdc_n1569, U_dsdc_n1568,
         U_dsdc_n1567, U_dsdc_n1566, U_dsdc_n1565, U_dsdc_n1564, U_dsdc_n1563,
         U_dsdc_n1562, U_dsdc_n1561, U_dsdc_n1560, U_dsdc_n1559, U_dsdc_n1558,
         U_dsdc_n1557, U_dsdc_n1556, U_dsdc_n1555, U_dsdc_n1554, U_dsdc_n1553,
         U_dsdc_n1552, U_dsdc_n1551, U_dsdc_n1550, U_dsdc_n1549, U_dsdc_n1548,
         U_dsdc_n1547, U_dsdc_n1546, U_dsdc_n1545, U_dsdc_n1544, U_dsdc_n1543,
         U_dsdc_n1542, U_dsdc_n1541, U_dsdc_n1540, U_dsdc_n1539, U_dsdc_n1538,
         U_dsdc_n1537, U_dsdc_n1536, U_dsdc_n1535, U_dsdc_n1534, U_dsdc_n1533,
         U_dsdc_n1532, U_dsdc_n1531, U_dsdc_n1530, U_dsdc_n1529, U_dsdc_n1528,
         U_dsdc_n1527, U_dsdc_n1526, U_dsdc_n1525, U_dsdc_n1524, U_dsdc_n1523,
         U_dsdc_n1522, U_dsdc_n1521, U_dsdc_n1520, U_dsdc_n1519, U_dsdc_n1518,
         U_dsdc_n1517, U_dsdc_n1516, U_dsdc_n1515, U_dsdc_n1514, U_dsdc_n1513,
         U_dsdc_n1512, U_dsdc_n1511, U_dsdc_n1510, U_dsdc_n1509, U_dsdc_n1508,
         U_dsdc_n1507, U_dsdc_n1506, U_dsdc_n1505, U_dsdc_n1504, U_dsdc_n1503,
         U_dsdc_n1502, U_dsdc_n1501, U_dsdc_n1500, U_dsdc_n1499, U_dsdc_n1498,
         U_dsdc_n1497, U_dsdc_n1496, U_dsdc_n1495, U_dsdc_n1493, U_dsdc_n1492,
         U_dsdc_n1491, U_dsdc_n1490, U_dsdc_n1489, U_dsdc_n1488, U_dsdc_n1487,
         U_dsdc_n1486, U_dsdc_n1485, U_dsdc_n1484, U_dsdc_n1483, U_dsdc_n1482,
         U_dsdc_n1481, U_dsdc_n1480, U_dsdc_n1479, U_dsdc_n1478, U_dsdc_n1477,
         U_dsdc_n1476, U_dsdc_n1475, U_dsdc_n1474, U_dsdc_n1473, U_dsdc_n1472,
         U_dsdc_n1471, U_dsdc_n1470, U_dsdc_n1469, U_dsdc_n1468, U_dsdc_n1467,
         U_dsdc_n1466, U_dsdc_n1465, U_dsdc_n1464, U_dsdc_n1462, U_dsdc_n1461,
         U_dsdc_n1460, U_dsdc_n1458, U_dsdc_n1457, U_dsdc_n1456, U_dsdc_n1455,
         U_dsdc_n1454, U_dsdc_n1453, U_dsdc_n1452, U_dsdc_n1451, U_dsdc_n1450,
         U_dsdc_n1449, U_dsdc_n1448, U_dsdc_n1447, U_dsdc_n1446, U_dsdc_n1445,
         U_dsdc_n1444, U_dsdc_n1438, U_dsdc_n1437, U_dsdc_n1436, U_dsdc_n1435,
         U_dsdc_n1434, U_dsdc_n1433, U_dsdc_n1432, U_dsdc_n1431, U_dsdc_n1430,
         U_dsdc_n1429, U_dsdc_n1428, U_dsdc_n1427, U_dsdc_n1426, U_dsdc_n1425,
         U_dsdc_n1424, U_dsdc_n1423, U_dsdc_n1422, U_dsdc_n1421, U_dsdc_n1420,
         U_dsdc_n1419, U_dsdc_n1418, U_dsdc_n1417, U_dsdc_n1416, U_dsdc_n1415,
         U_dsdc_n1414, U_dsdc_n1413, U_dsdc_n1412, U_dsdc_n1411, U_dsdc_n1410,
         U_dsdc_n1409, U_dsdc_n1408, U_dsdc_n1407, U_dsdc_n1406, U_dsdc_n1405,
         U_dsdc_n1404, U_dsdc_n1403, U_dsdc_n1402, U_dsdc_n1401, U_dsdc_n1400,
         U_dsdc_n1399, U_dsdc_n1398, U_dsdc_n1397, U_dsdc_n1396, U_dsdc_n1395,
         U_dsdc_n1394, U_dsdc_n1393, U_dsdc_n1392, U_dsdc_n1391, U_dsdc_n1390,
         U_dsdc_n1389, U_dsdc_n1388, U_dsdc_n1387, U_dsdc_n1386, U_dsdc_n1385,
         U_dsdc_n1384, U_dsdc_n1383, U_dsdc_n1382, U_dsdc_n1381, U_dsdc_n1380,
         U_dsdc_n1379, U_dsdc_n1377, U_dsdc_n1376, U_dsdc_n1375, U_dsdc_n1374,
         U_dsdc_n1373, U_dsdc_n1372, U_dsdc_n1371, U_dsdc_n1370, U_dsdc_n1369,
         U_dsdc_n1368, U_dsdc_n1367, U_dsdc_n1366, U_dsdc_n1365, U_dsdc_n1364,
         U_dsdc_n1363, U_dsdc_n1362, U_dsdc_n1361, U_dsdc_n1360, U_dsdc_n1359,
         U_dsdc_n1358, U_dsdc_n1357, U_dsdc_n1356, U_dsdc_n1355, U_dsdc_n1354,
         U_dsdc_n1353, U_dsdc_n1352, U_dsdc_n1351, U_dsdc_n1350, U_dsdc_n1349,
         U_dsdc_n1348, U_dsdc_n1347, U_dsdc_n1346, U_dsdc_n1345, U_dsdc_n1344,
         U_dsdc_n1343, U_dsdc_n1342, U_dsdc_n1341, U_dsdc_n1340, U_dsdc_n1339,
         U_dsdc_n1338, U_dsdc_n1337, U_dsdc_n1336, U_dsdc_n1335, U_dsdc_n1334,
         U_dsdc_n1333, U_dsdc_n1332, U_dsdc_n1331, U_dsdc_n1330, U_dsdc_n1329,
         U_dsdc_n1328, U_dsdc_n1327, U_dsdc_n1326, U_dsdc_n1325, U_dsdc_n1324,
         U_dsdc_n1323, U_dsdc_n1322, U_dsdc_n1321, U_dsdc_n1320, U_dsdc_n1319,
         U_dsdc_n1318, U_dsdc_n1317, U_dsdc_n1316, U_dsdc_n1315, U_dsdc_n1314,
         U_dsdc_n1313, U_dsdc_n1312, U_dsdc_n1311, U_dsdc_n1310, U_dsdc_n1309,
         U_dsdc_n1308, U_dsdc_n1307, U_dsdc_n1306, U_dsdc_n1305, U_dsdc_n1304,
         U_dsdc_n1303, U_dsdc_n1302, U_dsdc_n1301, U_dsdc_n1300, U_dsdc_n1299,
         U_dsdc_n1298, U_dsdc_n1297, U_dsdc_n1296, U_dsdc_n1295, U_dsdc_n1294,
         U_dsdc_n1293, U_dsdc_n1292, U_dsdc_n1291, U_dsdc_n1290, U_dsdc_n1289,
         U_dsdc_n1288, U_dsdc_n1287, U_dsdc_n1286, U_dsdc_n1285, U_dsdc_n1284,
         U_dsdc_n1283, U_dsdc_n1282, U_dsdc_n1281, U_dsdc_n1280, U_dsdc_n1279,
         U_dsdc_n1278, U_dsdc_n1277, U_dsdc_n1276, U_dsdc_n1275, U_dsdc_n1274,
         U_dsdc_n1273, U_dsdc_n1272, U_dsdc_n1271, U_dsdc_n1270, U_dsdc_n1269,
         U_dsdc_n1268, U_dsdc_n1267, U_dsdc_n1266, U_dsdc_n1264, U_dsdc_n1263,
         U_dsdc_n1262, U_dsdc_n1261, U_dsdc_n1260, U_dsdc_n1259, U_dsdc_n1258,
         U_dsdc_n1254, U_dsdc_n1253, U_dsdc_n1252, U_dsdc_n1251, U_dsdc_n1250,
         U_dsdc_n1249, U_dsdc_n1248, U_dsdc_n1247, U_dsdc_n1246, U_dsdc_n1245,
         U_dsdc_n1244, U_dsdc_n1243, U_dsdc_n1241, U_dsdc_n1239, U_dsdc_n1238,
         U_dsdc_n1237, U_dsdc_n1235, U_dsdc_n1234, U_dsdc_n1233, U_dsdc_n1231,
         U_dsdc_n1229, U_dsdc_n1228, U_dsdc_n1227, U_dsdc_n1225, U_dsdc_n1224,
         U_dsdc_n1223, U_dsdc_n1222, U_dsdc_n1221, U_dsdc_n1220, U_dsdc_n1219,
         U_dsdc_n1218, U_dsdc_n1217, U_dsdc_n1216, U_dsdc_n1215, U_dsdc_n1214,
         U_dsdc_n1213, U_dsdc_n1212, U_dsdc_n1211, U_dsdc_n1210, U_dsdc_n1209,
         U_dsdc_n1208, U_dsdc_n1207, U_dsdc_n1206, U_dsdc_n1205, U_dsdc_n1204,
         U_dsdc_n1203, U_dsdc_n1202, U_dsdc_n1201, U_dsdc_n1200, U_dsdc_n1199,
         U_dsdc_n1198, U_dsdc_n1197, U_dsdc_n1196, U_dsdc_n1195, U_dsdc_n1194,
         U_dsdc_n1193, U_dsdc_n1192, U_dsdc_n1191, U_dsdc_n1190, U_dsdc_n1189,
         U_dsdc_n1188, U_dsdc_n1187, U_dsdc_n1186, U_dsdc_n1185, U_dsdc_n1184,
         U_dsdc_n1183, U_dsdc_n1182, U_dsdc_n1181, U_dsdc_n1180, U_dsdc_n1179,
         U_dsdc_n1178, U_dsdc_n1177, U_dsdc_n1176, U_dsdc_n1175, U_dsdc_n1174,
         U_dsdc_n1173, U_dsdc_n1172, U_dsdc_n1171, U_dsdc_n1170, U_dsdc_n1169,
         U_dsdc_n1168, U_dsdc_n1167, U_dsdc_n1166, U_dsdc_n1165, U_dsdc_n1164,
         U_dsdc_n1163, U_dsdc_n1162, U_dsdc_n1161, U_dsdc_n1160, U_dsdc_n1159,
         U_dsdc_n1158, U_dsdc_n1157, U_dsdc_n1156, U_dsdc_n1155, U_dsdc_n1154,
         U_dsdc_n1153, U_dsdc_n1152, U_dsdc_n1151, U_dsdc_n1150, U_dsdc_n1149,
         U_dsdc_n1148, U_dsdc_n1147, U_dsdc_n1146, U_dsdc_n1145, U_dsdc_n1144,
         U_dsdc_n1143, U_dsdc_n1142, U_dsdc_n1141, U_dsdc_n1140, U_dsdc_n1139,
         U_dsdc_n1138, U_dsdc_n1137, U_dsdc_n1136, U_dsdc_n1135, U_dsdc_n1134,
         U_dsdc_n1133, U_dsdc_n1132, U_dsdc_n1131, U_dsdc_n1130, U_dsdc_n1129,
         U_dsdc_n1128, U_dsdc_n1127, U_dsdc_n1126, U_dsdc_n1125, U_dsdc_n1124,
         U_dsdc_n1123, U_dsdc_n1122, U_dsdc_n1121, U_dsdc_n1119, U_dsdc_n1118,
         U_dsdc_n1117, U_dsdc_n1116, U_dsdc_n1115, U_dsdc_n1114, U_dsdc_n1113,
         U_dsdc_n1112, U_dsdc_n1111, U_dsdc_n1110, U_dsdc_n1109, U_dsdc_n1108,
         U_dsdc_n1107, U_dsdc_n1106, U_dsdc_n1105, U_dsdc_n1104, U_dsdc_n1103,
         U_dsdc_n1101, U_dsdc_n1100, U_dsdc_n1099, U_dsdc_n1098, U_dsdc_n1097,
         U_dsdc_n1096, U_dsdc_n1095, U_dsdc_n1094, U_dsdc_n1093, U_dsdc_n1092,
         U_dsdc_n1091, U_dsdc_n1090, U_dsdc_n1089, U_dsdc_n1088, U_dsdc_n1087,
         U_dsdc_n1085, U_dsdc_n1084, U_dsdc_n1082, U_dsdc_n1081, U_dsdc_n1079,
         U_dsdc_n1078, U_dsdc_n1077, U_dsdc_n1076, U_dsdc_n1075, U_dsdc_n1074,
         U_dsdc_n1073, U_dsdc_n1072, U_dsdc_n1071, U_dsdc_n1070, U_dsdc_n1069,
         U_dsdc_n1068, U_dsdc_n1067, U_dsdc_n1066, U_dsdc_n1065, U_dsdc_n1064,
         U_dsdc_n1063, U_dsdc_n1062, U_dsdc_n1061, U_dsdc_n1060, U_dsdc_n1059,
         U_dsdc_n1058, U_dsdc_n1057, U_dsdc_n1056, U_dsdc_n1053, U_dsdc_n1052,
         U_dsdc_n1051, U_dsdc_n1050, U_dsdc_n1049, U_dsdc_n1048, U_dsdc_n1047,
         U_dsdc_n1046, U_dsdc_n1045, U_dsdc_n1044, U_dsdc_n1043, U_dsdc_n1042,
         U_dsdc_n1041, U_dsdc_n1040, U_dsdc_n1039, U_dsdc_n1038, U_dsdc_n1037,
         U_dsdc_n1036, U_dsdc_n1035, U_dsdc_n1033, U_dsdc_n1032, U_dsdc_n1031,
         U_dsdc_n1030, U_dsdc_n1029, U_dsdc_n1028, U_dsdc_n1027, U_dsdc_n1026,
         U_dsdc_n1025, U_dsdc_n1024, U_dsdc_n1023, U_dsdc_n1022, U_dsdc_n1021,
         U_dsdc_n1020, U_dsdc_n1019, U_dsdc_n1018, U_dsdc_n1017, U_dsdc_n1016,
         U_dsdc_n1015, U_dsdc_n1014, U_dsdc_n1013, U_dsdc_n1012, U_dsdc_n1011,
         U_dsdc_n1010, U_dsdc_n1009, U_dsdc_n1008, U_dsdc_n1007, U_dsdc_n1006,
         U_dsdc_n1005, U_dsdc_n1004, U_dsdc_n1003, U_dsdc_n1002, U_dsdc_n1001,
         U_dsdc_n1000, U_dsdc_n999, U_dsdc_n998, U_dsdc_n997, U_dsdc_n996,
         U_dsdc_n995, U_dsdc_n994, U_dsdc_n993, U_dsdc_n992, U_dsdc_n991,
         U_dsdc_n990, U_dsdc_n989, U_dsdc_n988, U_dsdc_n987, U_dsdc_n986,
         U_dsdc_n985, U_dsdc_n984, U_dsdc_n983, U_dsdc_n982, U_dsdc_n981,
         U_dsdc_n980, U_dsdc_n979, U_dsdc_n978, U_dsdc_n977, U_dsdc_n976,
         U_dsdc_n975, U_dsdc_n974, U_dsdc_n973, U_dsdc_n972, U_dsdc_n971,
         U_dsdc_n970, U_dsdc_n969, U_dsdc_n968, U_dsdc_n967, U_dsdc_n966,
         U_dsdc_n965, U_dsdc_n964, U_dsdc_n963, U_dsdc_n962, U_dsdc_n961,
         U_dsdc_n960, U_dsdc_n959, U_dsdc_n958, U_dsdc_n957, U_dsdc_n956,
         U_dsdc_n955, U_dsdc_n954, U_dsdc_n953, U_dsdc_n952, U_dsdc_n951,
         U_dsdc_n950, U_dsdc_n949, U_dsdc_n948, U_dsdc_n947, U_dsdc_n946,
         U_dsdc_n945, U_dsdc_n944, U_dsdc_n943, U_dsdc_n942, U_dsdc_n941,
         U_dsdc_n940, U_dsdc_n939, U_dsdc_n938, U_dsdc_n937, U_dsdc_n936,
         U_dsdc_n935, U_dsdc_n934, U_dsdc_n933, U_dsdc_n932, U_dsdc_n931,
         U_dsdc_n930, U_dsdc_n929, U_dsdc_n928, U_dsdc_n927, U_dsdc_n926,
         U_dsdc_n925, U_dsdc_n924, U_dsdc_n923, U_dsdc_n922, U_dsdc_n921,
         U_dsdc_n920, U_dsdc_n919, U_dsdc_n918, U_dsdc_n917, U_dsdc_n916,
         U_dsdc_n915, U_dsdc_n914, U_dsdc_n913, U_dsdc_n912, U_dsdc_n911,
         U_dsdc_n910, U_dsdc_n909, U_dsdc_n908, U_dsdc_n907, U_dsdc_n906,
         U_dsdc_n905, U_dsdc_n904, U_dsdc_n903, U_dsdc_n902, U_dsdc_n901,
         U_dsdc_n900, U_dsdc_n899, U_dsdc_n898, U_dsdc_n897, U_dsdc_n896,
         U_dsdc_n895, U_dsdc_n894, U_dsdc_n893, U_dsdc_n892, U_dsdc_n891,
         U_dsdc_n890, U_dsdc_n889, U_dsdc_n887, U_dsdc_n886, U_dsdc_n885,
         U_dsdc_n884, U_dsdc_n883, U_dsdc_n881, U_dsdc_n880, U_dsdc_n879,
         U_dsdc_n878, U_dsdc_n877, U_dsdc_n876, U_dsdc_n875, U_dsdc_n874,
         U_dsdc_n873, U_dsdc_n872, U_dsdc_n871, U_dsdc_n870, U_dsdc_n869,
         U_dsdc_n868, U_dsdc_n867, U_dsdc_n866, U_dsdc_n865, U_dsdc_n864,
         U_dsdc_n863, U_dsdc_n862, U_dsdc_n861, U_dsdc_n860, U_dsdc_n859,
         U_dsdc_n858, U_dsdc_n857, U_dsdc_n856, U_dsdc_n855, U_dsdc_n854,
         U_dsdc_n853, U_dsdc_n852, U_dsdc_n851, U_dsdc_n850, U_dsdc_n849,
         U_dsdc_n848, U_dsdc_n847, U_dsdc_n846, U_dsdc_n845, U_dsdc_n844,
         U_dsdc_n843, U_dsdc_n842, U_dsdc_n841, U_dsdc_n840, U_dsdc_n839,
         U_dsdc_n838, U_dsdc_n837, U_dsdc_n836, U_dsdc_n835, U_dsdc_n834,
         U_dsdc_n833, U_dsdc_n832, U_dsdc_n831, U_dsdc_n830, U_dsdc_n829,
         U_dsdc_n828, U_dsdc_n827, U_dsdc_n826, U_dsdc_n825, U_dsdc_n824,
         U_dsdc_n822, U_dsdc_n821, U_dsdc_n820, U_dsdc_n819, U_dsdc_n818,
         U_dsdc_n817, U_dsdc_n816, U_dsdc_n815, U_dsdc_n814, U_dsdc_n813,
         U_dsdc_n812, U_dsdc_n810, U_dsdc_n809, U_dsdc_n808, U_dsdc_n807,
         U_dsdc_n806, U_dsdc_n805, U_dsdc_n804, U_dsdc_n803, U_dsdc_n802,
         U_dsdc_n801, U_dsdc_n800, U_dsdc_n799, U_dsdc_n798, U_dsdc_n797,
         U_dsdc_n796, U_dsdc_n795, U_dsdc_n794, U_dsdc_n793, U_dsdc_n792,
         U_dsdc_n791, U_dsdc_n790, U_dsdc_n789, U_dsdc_n788, U_dsdc_n787,
         U_dsdc_n786, U_dsdc_n785, U_dsdc_n784, U_dsdc_n783, U_dsdc_n782,
         U_dsdc_n778, U_dsdc_n777, U_dsdc_n776, U_dsdc_n775, U_dsdc_n774,
         U_dsdc_n773, U_dsdc_n772, U_dsdc_n770, U_dsdc_n767, U_dsdc_n766,
         U_dsdc_n765, U_dsdc_n764, U_dsdc_n763, U_dsdc_n762, U_dsdc_n761,
         U_dsdc_n760, U_dsdc_n759, U_dsdc_n758, U_dsdc_n757, U_dsdc_n756,
         U_dsdc_n755, U_dsdc_n754, U_dsdc_n753, U_dsdc_n752, U_dsdc_n751,
         U_dsdc_n750, U_dsdc_n749, U_dsdc_n748, U_dsdc_n747, U_dsdc_n746,
         U_dsdc_n745, U_dsdc_n744, U_dsdc_n741, U_dsdc_n740, U_dsdc_n739,
         U_dsdc_n738, U_dsdc_n737, U_dsdc_n736, U_dsdc_n735, U_dsdc_n734,
         U_dsdc_n733, U_dsdc_n732, U_dsdc_n731, U_dsdc_n730, U_dsdc_n729,
         U_dsdc_n728, U_dsdc_n727, U_dsdc_n726, U_dsdc_n725, U_dsdc_n724,
         U_dsdc_n723, U_dsdc_n722, U_dsdc_n721, U_dsdc_n720, U_dsdc_n719,
         U_dsdc_n718, U_dsdc_n717, U_dsdc_n716, U_dsdc_n715, U_dsdc_n714,
         U_dsdc_n713, U_dsdc_n712, U_dsdc_n711, U_dsdc_n710, U_dsdc_n708,
         U_dsdc_n705, U_dsdc_n704, U_dsdc_n703, U_dsdc_n702, U_dsdc_n701,
         U_dsdc_n700, U_dsdc_n699, U_dsdc_n698, U_dsdc_n697, U_dsdc_n696,
         U_dsdc_n695, U_dsdc_n694, U_dsdc_n693, U_dsdc_n692, U_dsdc_n691,
         U_dsdc_n690, U_dsdc_n689, U_dsdc_n688, U_dsdc_n687, U_dsdc_n686,
         U_dsdc_n685, U_dsdc_n684, U_dsdc_n683, U_dsdc_n682, U_dsdc_n681,
         U_dsdc_n680, U_dsdc_n679, U_dsdc_n678, U_dsdc_n677, U_dsdc_n676,
         U_dsdc_n675, U_dsdc_n674, U_dsdc_n673, U_dsdc_n672, U_dsdc_n671,
         U_dsdc_n670, U_dsdc_n669, U_dsdc_n668, U_dsdc_n667, U_dsdc_n666,
         U_dsdc_n663, U_dsdc_n662, U_dsdc_n661, U_dsdc_n660, U_dsdc_n659,
         U_dsdc_n658, U_dsdc_n657, U_dsdc_n654, U_dsdc_n653, U_dsdc_n652,
         U_dsdc_n651, U_dsdc_n650, U_dsdc_n649, U_dsdc_n648, U_dsdc_n646,
         U_dsdc_n645, U_dsdc_n644, U_dsdc_n643, U_dsdc_n642, U_dsdc_n641,
         U_dsdc_n621, U_dsdc_n620, U_dsdc_n619, U_dsdc_n618, U_dsdc_n617,
         U_dsdc_n616, U_dsdc_n615, U_dsdc_n614, U_dsdc_n613, U_dsdc_n612,
         U_dsdc_n611, U_dsdc_n610, U_dsdc_n609, U_dsdc_n608, U_dsdc_n607,
         U_dsdc_n606, U_dsdc_n605, U_dsdc_n604, U_dsdc_n603, U_dsdc_n602,
         U_dsdc_n601, U_dsdc_n600, U_dsdc_n599, U_dsdc_n598, U_dsdc_n597,
         U_dsdc_n596, U_dsdc_n595, U_dsdc_n594, U_dsdc_n593, U_dsdc_n592,
         U_dsdc_n591, U_dsdc_n590, U_dsdc_n589, U_dsdc_n588, U_dsdc_n587,
         U_dsdc_n586, U_dsdc_n585, U_dsdc_n584, U_dsdc_n583, U_dsdc_n582,
         U_dsdc_n581, U_dsdc_n580, U_dsdc_n579, U_dsdc_n578, U_dsdc_n577,
         U_dsdc_n576, U_dsdc_n575, U_dsdc_n574, U_dsdc_n573, U_dsdc_n572,
         U_dsdc_n571, U_dsdc_n570, U_dsdc_n569, U_dsdc_n568, U_dsdc_n567,
         U_dsdc_n566, U_dsdc_n565, U_dsdc_n564, U_dsdc_n563, U_dsdc_n562,
         U_dsdc_n561, U_dsdc_n560, U_dsdc_n559, U_dsdc_n558, U_dsdc_n557,
         U_dsdc_n556, U_dsdc_n555, U_dsdc_n553, U_dsdc_n552, U_dsdc_n551,
         U_dsdc_n550, U_dsdc_n549, U_dsdc_n548, U_dsdc_n547, U_dsdc_n546,
         U_dsdc_n545, U_dsdc_n544, U_dsdc_n543, U_dsdc_n542, U_dsdc_n541,
         U_dsdc_n540, U_dsdc_n539, U_dsdc_n538, U_dsdc_n537, U_dsdc_n536,
         U_dsdc_n535, U_dsdc_n534, U_dsdc_n533, U_dsdc_n532, U_dsdc_n531,
         U_dsdc_n530, U_dsdc_n529, U_dsdc_n528, U_dsdc_n527, U_dsdc_n526,
         U_dsdc_n525, U_dsdc_n524, U_dsdc_n523, U_dsdc_n522, U_dsdc_n519,
         U_dsdc_n517, U_dsdc_n516, U_dsdc_n515, U_dsdc_n514, U_dsdc_n513,
         U_dsdc_n512, U_dsdc_n511, U_dsdc_n510, U_dsdc_n509, U_dsdc_n508,
         U_dsdc_n507, U_dsdc_n504, U_dsdc_n503, U_dsdc_n502, U_dsdc_n501,
         U_dsdc_n500, U_dsdc_n499, U_dsdc_n498, U_dsdc_n497, U_dsdc_n496,
         U_dsdc_n495, U_dsdc_n494, U_dsdc_n493, U_dsdc_n492, U_dsdc_n491,
         U_dsdc_n488, U_dsdc_n487, U_dsdc_n486, U_dsdc_n485, U_dsdc_n484,
         U_dsdc_n483, U_dsdc_n482, U_dsdc_n481, U_dsdc_n480, U_dsdc_n479,
         U_dsdc_n478, U_dsdc_n477, U_dsdc_n476, U_dsdc_n475, U_dsdc_n474,
         U_dsdc_n473, U_dsdc_n472, U_dsdc_n471, U_dsdc_n470, U_dsdc_n469,
         U_dsdc_n468, U_dsdc_n467, U_dsdc_n466, U_dsdc_n465, U_dsdc_n464,
         U_dsdc_n463, U_dsdc_n462, U_dsdc_n461, U_dsdc_n460, U_dsdc_n459,
         U_dsdc_n458, U_dsdc_n457, U_dsdc_n456, U_dsdc_n455, U_dsdc_n454,
         U_dsdc_n453, U_dsdc_n452, U_dsdc_n451, U_dsdc_n450, U_dsdc_n449,
         U_dsdc_n448, U_dsdc_n447, U_dsdc_n446, U_dsdc_n445, U_dsdc_n444,
         U_dsdc_n443, U_dsdc_n442, U_dsdc_n441, U_dsdc_n440, U_dsdc_n439,
         U_dsdc_n438, U_dsdc_n437, U_dsdc_n436, U_dsdc_n435, U_dsdc_n434,
         U_dsdc_n433, U_dsdc_n432, U_dsdc_n430, U_dsdc_n429, U_dsdc_n428,
         U_dsdc_n427, U_dsdc_n426, U_dsdc_n425, U_dsdc_n424, U_dsdc_n422,
         U_dsdc_n421, U_dsdc_n420, U_dsdc_n419, U_dsdc_n402, U_dsdc_n401,
         U_dsdc_n400, U_dsdc_n399, U_dsdc_n398, U_dsdc_n397, U_dsdc_n396,
         U_dsdc_n395, U_dsdc_n385, U_dsdc_n384, U_dsdc_n383, U_dsdc_n382,
         U_dsdc_n365, U_dsdc_n364, U_dsdc_n363, U_dsdc_n362, U_dsdc_n361,
         U_dsdc_n360, U_dsdc_n359, U_dsdc_n358, U_dsdc_n357, U_dsdc_n356,
         U_dsdc_n355, U_dsdc_n354, U_dsdc_n353, U_dsdc_n352, U_dsdc_n351,
         U_dsdc_n350, U_dsdc_n349, U_dsdc_n347, U_dsdc_n346, U_dsdc_n345,
         U_dsdc_n344, U_dsdc_n343, U_dsdc_n342, U_dsdc_n341, U_dsdc_n340,
         U_dsdc_n339, U_dsdc_n338, U_dsdc_n337, U_dsdc_n336, U_dsdc_n335,
         U_dsdc_n334, U_dsdc_n333, U_dsdc_n332, U_dsdc_n331, U_dsdc_n330,
         U_dsdc_n328, U_dsdc_n327, U_dsdc_n326, U_dsdc_n325, U_dsdc_n318,
         U_dsdc_n314, U_dsdc_n312, U_dsdc_n309, U_dsdc_n308, U_dsdc_n306,
         U_dsdc_n305, U_dsdc_n304, U_dsdc_n303, U_dsdc_n302, U_dsdc_n301,
         U_dsdc_n299, U_dsdc_n298, U_dsdc_n292, U_dsdc_n284, U_dsdc_n239,
         U_dsdc_n208, U_dsdc_n207, U_dsdc_n206, U_dsdc_n205, U_dsdc_n204,
         U_dsdc_n203, U_dsdc_n202, U_dsdc_n201, U_dsdc_n200, U_dsdc_n199,
         U_dsdc_n198, U_dsdc_n197, U_dsdc_n196, U_dsdc_n195, U_dsdc_n194,
         U_dsdc_n193, U_dsdc_n192, U_dsdc_n191, U_dsdc_n190, U_dsdc_n189,
         U_dsdc_n188, U_dsdc_n187, U_dsdc_n186, U_dsdc_n185, U_dsdc_n184,
         U_dsdc_n183, U_dsdc_n182, U_dsdc_n181, U_dsdc_n180, U_dsdc_n179,
         U_dsdc_n178, U_dsdc_n177, U_dsdc_n176, U_dsdc_n174, U_dsdc_n173,
         U_dsdc_n172, U_dsdc_n171, U_dsdc_n170, U_dsdc_n169, U_dsdc_n168,
         U_dsdc_n167, U_dsdc_n166, U_dsdc_n165, U_dsdc_n164, U_dsdc_n163,
         U_dsdc_n162, U_dsdc_n159, U_dsdc_n158, U_dsdc_n157, U_dsdc_n156,
         U_dsdc_n155, U_dsdc_n154, U_dsdc_n153, U_dsdc_n152, U_dsdc_n151,
         U_dsdc_n150, U_dsdc_n149, U_dsdc_n148, U_dsdc_n147, U_dsdc_n145,
         U_dsdc_n144, U_dsdc_n143, U_dsdc_n142, U_dsdc_n141, U_dsdc_n140,
         U_dsdc_n139, U_dsdc_n137, U_dsdc_n134, U_dsdc_n133, U_dsdc_n131,
         U_dsdc_n130, U_dsdc_n129, U_dsdc_n128, U_dsdc_n126, U_dsdc_n125,
         U_dsdc_n124, U_dsdc_n123, U_dsdc_n121, U_dsdc_n120, U_dsdc_n119,
         U_dsdc_n118, U_dsdc_n117, U_dsdc_n116, U_dsdc_n115, U_dsdc_n114,
         U_dsdc_n113, U_dsdc_n112, U_dsdc_n111, U_dsdc_n109, U_dsdc_n108,
         U_dsdc_n107, U_dsdc_n106, U_dsdc_n105, U_dsdc_n104, U_dsdc_n103,
         U_dsdc_n102, U_dsdc_n101, U_dsdc_n100, U_dsdc_n99, U_dsdc_n98,
         U_dsdc_n97, U_dsdc_n96, U_dsdc_n95, U_dsdc_n94, U_dsdc_n93,
         U_dsdc_n92, U_dsdc_n91, U_dsdc_n90, U_dsdc_n89, U_dsdc_n88,
         U_dsdc_n87, U_dsdc_n86, U_dsdc_n84, U_dsdc_n82, U_dsdc_n81,
         U_dsdc_n80, U_dsdc_n79, U_dsdc_n78, U_dsdc_n75, U_dsdc_n74,
         U_dsdc_n73, U_dsdc_n72, U_dsdc_n71, U_dsdc_n70, U_dsdc_n69,
         U_dsdc_n68, U_dsdc_n67, U_dsdc_n66, U_dsdc_n65, U_dsdc_n63,
         U_dsdc_n62, U_dsdc_n60, U_dsdc_n59, U_dsdc_n58, U_dsdc_n57,
         U_dsdc_n56, U_dsdc_n53, U_dsdc_n52, U_dsdc_n51, U_dsdc_n50,
         U_dsdc_n49, U_dsdc_n48, U_dsdc_n47, U_dsdc_n46, U_dsdc_n45,
         U_dsdc_n44, U_dsdc_n43, U_dsdc_n42, U_dsdc_n41, U_dsdc_n40,
         U_dsdc_n39, U_dsdc_n38, U_dsdc_n37, U_dsdc_n36, U_dsdc_n35,
         U_dsdc_n34, U_dsdc_n33, U_dsdc_n32, U_dsdc_n31, U_dsdc_n30,
         U_dsdc_n29, U_dsdc_n28, U_dsdc_n27, U_dsdc_n26, U_dsdc_n25,
         U_dsdc_n24, U_dsdc_n23, U_dsdc_n22, U_dsdc_n20, U_dsdc_n19,
         U_dsdc_n18, U_dsdc_n17, U_dsdc_n16, U_dsdc_n15, U_dsdc_n14,
         U_dsdc_n12, U_dsdc_n11, U_dsdc_n10, U_dsdc_n9, U_dsdc_n8, U_dsdc_n7,
         U_dsdc_n6, U_dsdc_n5, U_dsdc_n4, U_dsdc_n3, U_dsdc_n2, U_dsdc_n1,
         U_dsdc_DP_OP_1642_126_2028_n1, U_dsdc_DP_OP_1642_126_2028_n2,
         U_dsdc_DP_OP_1642_126_2028_n3, U_dsdc_DP_OP_1642_126_2028_n4,
         U_dsdc_DP_OP_1642_126_2028_n5, U_dsdc_DP_OP_1642_126_2028_n6,
         U_dsdc_DP_OP_1642_126_2028_n7, U_dsdc_DP_OP_1642_126_2028_n8,
         U_dsdc_DP_OP_1642_126_2028_n9, U_dsdc_DP_OP_1642_126_2028_n11,
         U_dsdc_DP_OP_1642_126_2028_n12, U_dsdc_DP_OP_1642_126_2028_n13,
         U_dsdc_DP_OP_1642_126_2028_n14, U_dsdc_DP_OP_1642_126_2028_n15,
         U_dsdc_DP_OP_1642_126_2028_n19, U_dsdc_DP_OP_1642_126_2028_n20,
         U_dsdc_DP_OP_1642_126_2028_n21, U_dsdc_DP_OP_1642_126_2028_n23,
         U_dsdc_DP_OP_1642_126_2028_n24, U_dsdc_DP_OP_1642_126_2028_n25,
         U_dsdc_DP_OP_1642_126_2028_n26, U_dsdc_DP_OP_1642_126_2028_n27,
         U_dsdc_DP_OP_1642_126_2028_n28, U_dsdc_DP_OP_1642_126_2028_n30,
         U_dsdc_DP_OP_1642_126_2028_n31, U_dsdc_DP_OP_1642_126_2028_n34,
         U_dsdc_DP_OP_1642_126_2028_n35, U_dsdc_DP_OP_1642_126_2028_n36,
         U_dsdc_DP_OP_1642_126_2028_n37, U_dsdc_DP_OP_1642_126_2028_n38,
         U_dsdc_DP_OP_1642_126_2028_n39, U_dsdc_DP_OP_1642_126_2028_n40,
         U_dsdc_DP_OP_1642_126_2028_n42, U_dsdc_DP_OP_1642_126_2028_n43,
         U_dsdc_DP_OP_1642_126_2028_n44, U_dsdc_DP_OP_1642_126_2028_n45,
         U_dsdc_DP_OP_1642_126_2028_n46, U_dsdc_DP_OP_1642_126_2028_n47,
         U_dsdc_DP_OP_1642_126_2028_n48, U_dsdc_DP_OP_1642_126_2028_n49,
         U_dsdc_DP_OP_1642_126_2028_n50, U_dsdc_DP_OP_1642_126_2028_n51,
         U_dsdc_DP_OP_1642_126_2028_n52, U_dsdc_DP_OP_1642_126_2028_n58,
         U_dsdc_DP_OP_1642_126_2028_n59, U_dsdc_DP_OP_1642_126_2028_n60,
         U_dsdc_DP_OP_1642_126_2028_n61, U_dsdc_DP_OP_1642_126_2028_n62,
         U_dsdc_DP_OP_1642_126_2028_n85, U_dsdc_DP_OP_1642_126_2028_n86,
         U_dsdc_DP_OP_1642_126_2028_I6, U_dsdc_DP_OP_1642_126_2028_I5_0_,
         U_dsdc_DP_OP_1642_126_2028_I5_1_, U_dsdc_DP_OP_1642_126_2028_I5_2_,
         U_dsdc_DP_OP_1642_126_2028_I5_3_, U_dsdc_DP_OP_1642_126_2028_I5_4_,
         U_dsdc_DP_OP_1642_126_2028_I5_5_, U_dsdc_DP_OP_1642_126_2028_I4,
         U_dsdc_RSOP_1683_C2_CONTROL1, U_dsdc_n554, U_dsdc_n431, U_dsdc_n423,
         U_dsdc_n418, U_dsdc_n417, U_dsdc_n416, U_dsdc_n415, U_dsdc_n414,
         U_dsdc_n413, U_dsdc_n412, U_dsdc_n411, U_dsdc_n410, U_dsdc_n409,
         U_dsdc_n408, U_dsdc_n407, U_dsdc_n406, U_dsdc_n405, U_dsdc_n404,
         U_dsdc_n403, U_dsdc_n394, U_dsdc_n393, U_dsdc_n392, U_dsdc_n391,
         U_dsdc_n390, U_dsdc_n389, U_dsdc_n388, U_dsdc_n387, U_dsdc_n386,
         U_dsdc_n381, U_dsdc_n380, U_dsdc_n379, U_dsdc_n378, U_dsdc_n377,
         U_dsdc_n376, U_dsdc_n375, U_dsdc_n374, U_dsdc_n373, U_dsdc_n372,
         U_dsdc_n371, U_dsdc_n370, U_dsdc_n369, U_dsdc_n368, U_dsdc_n367,
         U_dsdc_n366, U_dsdc_n348, U_dsdc_n329, U_dsdc_n324, U_dsdc_n323,
         U_dsdc_n322, U_dsdc_n321, U_dsdc_n320, U_dsdc_n319, U_dsdc_n317,
         U_dsdc_n316, U_dsdc_n315, U_dsdc_n313, U_dsdc_n310, U_dsdc_n307,
         U_dsdc_n300, U_dsdc_n297, U_dsdc_n296, U_dsdc_n295, U_dsdc_n294,
         U_dsdc_n293, U_dsdc_n291, U_dsdc_n290, U_dsdc_n289, U_dsdc_n288,
         U_dsdc_n287, U_dsdc_n286, U_dsdc_n283, U_dsdc_n282, U_dsdc_n281,
         U_dsdc_n280, U_dsdc_n279, U_dsdc_n278, U_dsdc_n277, U_dsdc_n276,
         U_dsdc_n275, U_dsdc_n274, U_dsdc_n273, U_dsdc_n272, U_dsdc_n271,
         U_dsdc_n270, U_dsdc_n269, U_dsdc_n268, U_dsdc_n267, U_dsdc_n266,
         U_dsdc_n265, U_dsdc_n264, U_dsdc_n263, U_dsdc_n262, U_dsdc_n261,
         U_dsdc_n260, U_dsdc_n259, U_dsdc_n258, U_dsdc_n257, U_dsdc_n256,
         U_dsdc_n255, U_dsdc_n254, U_dsdc_n253, U_dsdc_n252, U_dsdc_n251,
         U_dsdc_n250, U_dsdc_n249, U_dsdc_n248, U_dsdc_n247, U_dsdc_n246,
         U_dsdc_n245, U_dsdc_n244, U_dsdc_n243, U_dsdc_n242, U_dsdc_n241,
         U_dsdc_n240, U_dsdc_n238, U_dsdc_n237, U_dsdc_n236, U_dsdc_n235,
         U_dsdc_n234, U_dsdc_n233, U_dsdc_n232, U_dsdc_n231, U_dsdc_n230,
         U_dsdc_n229, U_dsdc_n228, U_dsdc_n227, U_dsdc_n226, U_dsdc_n225,
         U_dsdc_n224, U_dsdc_n223, U_dsdc_n222, U_dsdc_n221, U_dsdc_n220,
         U_dsdc_n219, U_dsdc_n218, U_dsdc_n217, U_dsdc_n216, U_dsdc_n215,
         U_dsdc_n214, U_dsdc_n213, U_dsdc_n212, U_dsdc_n211, U_dsdc_n210,
         U_dsdc_n209, U_dsdc_add_x_2600_1_n8, U_dsdc_C880_DATA5_5,
         U_dsdc_C880_DATA5_3, U_dsdc_C880_DATA5_1, U_dsdc_bm_bank_age_0__0_,
         U_dsdc_bm_bank_age_0__1_, U_dsdc_bm_bank_age_0__2_,
         U_dsdc_bm_bank_age_0__3_, U_dsdc_bm_bank_age_0__4_,
         U_dsdc_bm_bank_age_1__0_, U_dsdc_bm_bank_age_1__1_,
         U_dsdc_bm_bank_age_1__2_, U_dsdc_bm_bank_age_1__3_,
         U_dsdc_bm_bank_age_1__4_, U_dsdc_bm_bank_age_2__0_,
         U_dsdc_bm_bank_age_2__1_, U_dsdc_bm_bank_age_2__2_,
         U_dsdc_bm_bank_age_2__3_, U_dsdc_bm_bank_age_2__4_,
         U_dsdc_bm_bank_age_3__0_, U_dsdc_bm_bank_age_3__1_,
         U_dsdc_bm_bank_age_3__2_, U_dsdc_bm_bank_age_3__3_,
         U_dsdc_bm_bank_age_3__4_, U_dsdc_N4496, U_dsdc_N4492, U_dsdc_N4491,
         U_dsdc_N4490, U_dsdc_N4489, U_dsdc_N4488, U_dsdc_N4487, U_dsdc_N4486,
         U_dsdc_N4485, U_dsdc_N4484, U_dsdc_N4483, U_dsdc_N4482, U_dsdc_N4481,
         U_dsdc_N4480, U_dsdc_N4479, U_dsdc_N4478, U_dsdc_N4477, U_dsdc_N4476,
         U_dsdc_N4475, U_dsdc_N4474, U_dsdc_N4473, U_dsdc_N4463, U_dsdc_N4462,
         U_dsdc_N4461, U_dsdc_N4460, U_dsdc_N4449, U_dsdc_N4445, U_dsdc_N4444,
         U_dsdc_N4443, U_dsdc_N4442, U_dsdc_N4441, U_dsdc_N4440, U_dsdc_N4439,
         U_dsdc_N4438, U_dsdc_N4437, U_dsdc_N4436, U_dsdc_N4435, U_dsdc_N4434,
         U_dsdc_N4433, U_dsdc_N4432, U_dsdc_N4431, U_dsdc_N4430, U_dsdc_N4429,
         U_dsdc_N4428, U_dsdc_N4427, U_dsdc_N4426, U_dsdc_N4416, U_dsdc_N4415,
         U_dsdc_N4414, U_dsdc_N4413, U_dsdc_N4402, U_dsdc_N4398, U_dsdc_N4397,
         U_dsdc_N4396, U_dsdc_N4395, U_dsdc_N4394, U_dsdc_N4393, U_dsdc_N4392,
         U_dsdc_N4391, U_dsdc_N4390, U_dsdc_N4389, U_dsdc_N4388, U_dsdc_N4387,
         U_dsdc_N4386, U_dsdc_N4385, U_dsdc_N4384, U_dsdc_N4383, U_dsdc_N4382,
         U_dsdc_N4381, U_dsdc_N4380, U_dsdc_N4379, U_dsdc_N4369, U_dsdc_N4368,
         U_dsdc_N4367, U_dsdc_N4366, U_dsdc_N4355, U_dsdc_N4351, U_dsdc_N4350,
         U_dsdc_N4349, U_dsdc_N4348, U_dsdc_N4347, U_dsdc_N4346, U_dsdc_N4345,
         U_dsdc_N4344, U_dsdc_N4343, U_dsdc_N4342, U_dsdc_N4341, U_dsdc_N4340,
         U_dsdc_N4339, U_dsdc_N4338, U_dsdc_N4337, U_dsdc_N4336, U_dsdc_N4335,
         U_dsdc_N4334, U_dsdc_N4333, U_dsdc_N4332, U_dsdc_N4322, U_dsdc_N4321,
         U_dsdc_N4320, U_dsdc_N4319, U_dsdc_N4284, U_dsdc_N4283, U_dsdc_N4282,
         U_dsdc_N4281, U_dsdc_bm_ras_cnt_0__0_, U_dsdc_bm_ras_cnt_0__1_,
         U_dsdc_bm_ras_cnt_0__2_, U_dsdc_bm_ras_cnt_0__3_,
         U_dsdc_bm_ras_cnt_1__0_, U_dsdc_bm_ras_cnt_1__1_,
         U_dsdc_bm_ras_cnt_1__2_, U_dsdc_bm_ras_cnt_1__3_,
         U_dsdc_bm_ras_cnt_2__0_, U_dsdc_bm_ras_cnt_2__1_,
         U_dsdc_bm_ras_cnt_2__2_, U_dsdc_bm_ras_cnt_2__3_,
         U_dsdc_bm_ras_cnt_3__0_, U_dsdc_bm_ras_cnt_3__1_,
         U_dsdc_bm_ras_cnt_3__2_, U_dsdc_bm_ras_cnt_3__3_,
         U_dsdc_bm_rc_cnt_0__0_, U_dsdc_bm_rc_cnt_0__1_,
         U_dsdc_bm_rc_cnt_0__2_, U_dsdc_bm_rc_cnt_0__3_,
         U_dsdc_bm_rc_cnt_1__0_, U_dsdc_bm_rc_cnt_1__1_,
         U_dsdc_bm_rc_cnt_1__2_, U_dsdc_bm_rc_cnt_1__3_,
         U_dsdc_bm_rc_cnt_2__0_, U_dsdc_bm_rc_cnt_2__1_,
         U_dsdc_bm_rc_cnt_2__2_, U_dsdc_bm_rc_cnt_2__3_,
         U_dsdc_bm_rc_cnt_3__0_, U_dsdc_bm_rc_cnt_3__1_,
         U_dsdc_bm_rc_cnt_3__2_, U_dsdc_bm_rc_cnt_3__3_,
         U_dsdc_bm_row_addr_0__0_, U_dsdc_bm_row_addr_0__1_,
         U_dsdc_bm_row_addr_0__2_, U_dsdc_bm_row_addr_0__3_,
         U_dsdc_bm_row_addr_0__4_, U_dsdc_bm_row_addr_0__5_,
         U_dsdc_bm_row_addr_0__6_, U_dsdc_bm_row_addr_0__7_,
         U_dsdc_bm_row_addr_0__8_, U_dsdc_bm_row_addr_0__9_,
         U_dsdc_bm_row_addr_0__10_, U_dsdc_bm_row_addr_0__11_,
         U_dsdc_bm_row_addr_0__12_, U_dsdc_bm_row_addr_0__13_,
         U_dsdc_bm_row_addr_0__14_, U_dsdc_bm_row_addr_0__15_,
         U_dsdc_bm_row_addr_1__0_, U_dsdc_bm_row_addr_1__1_,
         U_dsdc_bm_row_addr_1__2_, U_dsdc_bm_row_addr_1__3_,
         U_dsdc_bm_row_addr_1__4_, U_dsdc_bm_row_addr_1__5_,
         U_dsdc_bm_row_addr_1__6_, U_dsdc_bm_row_addr_1__7_,
         U_dsdc_bm_row_addr_1__8_, U_dsdc_bm_row_addr_1__9_,
         U_dsdc_bm_row_addr_1__10_, U_dsdc_bm_row_addr_1__11_,
         U_dsdc_bm_row_addr_1__12_, U_dsdc_bm_row_addr_1__13_,
         U_dsdc_bm_row_addr_1__14_, U_dsdc_bm_row_addr_1__15_,
         U_dsdc_bm_row_addr_2__0_, U_dsdc_bm_row_addr_2__1_,
         U_dsdc_bm_row_addr_2__2_, U_dsdc_bm_row_addr_2__3_,
         U_dsdc_bm_row_addr_2__4_, U_dsdc_bm_row_addr_2__5_,
         U_dsdc_bm_row_addr_2__6_, U_dsdc_bm_row_addr_2__7_,
         U_dsdc_bm_row_addr_2__8_, U_dsdc_bm_row_addr_2__9_,
         U_dsdc_bm_row_addr_2__10_, U_dsdc_bm_row_addr_2__11_,
         U_dsdc_bm_row_addr_2__12_, U_dsdc_bm_row_addr_2__13_,
         U_dsdc_bm_row_addr_2__14_, U_dsdc_bm_row_addr_2__15_,
         U_dsdc_bm_row_addr_3__0_, U_dsdc_bm_row_addr_3__1_,
         U_dsdc_bm_row_addr_3__2_, U_dsdc_bm_row_addr_3__3_,
         U_dsdc_bm_row_addr_3__4_, U_dsdc_bm_row_addr_3__5_,
         U_dsdc_bm_row_addr_3__6_, U_dsdc_bm_row_addr_3__7_,
         U_dsdc_bm_row_addr_3__8_, U_dsdc_bm_row_addr_3__9_,
         U_dsdc_bm_row_addr_3__10_, U_dsdc_bm_row_addr_3__11_,
         U_dsdc_bm_row_addr_3__12_, U_dsdc_bm_row_addr_3__13_,
         U_dsdc_bm_row_addr_3__14_, U_dsdc_bm_row_addr_3__15_, U_dsdc_N4253,
         U_dsdc_N4252, U_dsdc_N4250, U_dsdc_N4248, U_dsdc_N4246, U_dsdc_N4244,
         U_dsdc_N4242, U_dsdc_N4241, U_dsdc_N4240, U_dsdc_N4239, U_dsdc_N4229,
         U_dsdc_N4228, U_dsdc_t_xp_cnt_0_, U_dsdc_t_xp_cnt_1_, U_dsdc_N4174,
         U_dsdc_N4141, U_dsdc_N4140, U_dsdc_N4139, U_dsdc_N4129, U_dsdc_N4128,
         U_dsdc_N4127, U_dsdc_N2002, U_dsdc_N1991, U_dsdc_N1990, U_dsdc_N1989,
         U_dsdc_N1988, U_dsdc_N1987, U_dsdc_N1767, U_dsdc_N1766, U_dsdc_N1765,
         U_dsdc_N1764, U_dsdc_N1763, U_dsdc_N1762, U_dsdc_N1685,
         U_dsdc_rcd_cnt_0_, U_dsdc_rcd_cnt_2_, U_dsdc_bm_num_open_bank_0_,
         U_dsdc_bm_num_open_bank_1_, U_dsdc_bm_num_open_bank_2_,
         U_dsdc_bm_num_open_bank_3_, U_dsdc_bm_num_open_bank_4_,
         U_dsdc_cas_latency_cnt_0_, U_dsdc_cas_latency_cnt_1_,
         U_dsdc_cas_latency_cnt_2_, U_dsdc_cas_latency_cnt_3_,
         U_dsdc_oldest_bank_0_, U_dsdc_oldest_bank_1_,
         U_dsdc_bm_ras_cnt_max_0_, U_dsdc_bm_ras_cnt_max_1_,
         U_dsdc_bm_ras_cnt_max_2_, U_dsdc_bm_ras_cnt_max_3_,
         U_dsdc_bm_bank_status_0_, U_dsdc_bm_bank_status_1_,
         U_dsdc_bm_bank_status_2_, U_dsdc_bm_bank_status_3_,
         U_dsdc_init_cnt_0_, U_dsdc_init_cnt_1_, U_dsdc_init_cnt_2_,
         U_dsdc_init_cnt_3_, U_dsdc_init_cnt_4_, U_dsdc_init_cnt_5_,
         U_dsdc_init_cnt_6_, U_dsdc_init_cnt_7_, U_dsdc_init_cnt_8_,
         U_dsdc_init_cnt_9_, U_dsdc_init_cnt_10_, U_dsdc_init_cnt_11_,
         U_dsdc_init_cnt_12_, U_dsdc_init_cnt_13_, U_dsdc_init_cnt_14_,
         U_dsdc_init_cnt_15_, U_dsdc_xsr_cnt_0_, U_dsdc_xsr_cnt_1_,
         U_dsdc_xsr_cnt_2_, U_dsdc_xsr_cnt_3_, U_dsdc_xsr_cnt_4_,
         U_dsdc_xsr_cnt_5_, U_dsdc_xsr_cnt_7_, U_dsdc_xsr_cnt_8_,
         U_dsdc_mrd_cnt_0_, U_dsdc_mrd_cnt_1_, U_dsdc_dqs_mask_end_nxt,
         U_dsdc_s_rd_end_nxt, U_dsdc_close_bank_addr_0_,
         U_dsdc_close_bank_addr_1_, U_dsdc_bm_close_bank_0_,
         U_dsdc_bm_close_bank_1_, U_dsdc_bm_close_bank_2_,
         U_dsdc_bm_close_bank_3_, U_dsdc_write_start_nxt,
         U_dsdc_wrapped_pop_flag_nxt, U_dsdc_cas_latency_1_,
         U_dsdc_cas_latency_2_, U_dsdc_N430, U_dsdc_auto_ref_en_nxt,
         U_dsdc_N429, U_dsdc_pre_amble_nxt, U_dsdc_N428, U_dsdc_N427,
         U_dsdc_N426, U_dsdc_N425, U_dsdc_N422, U_dsdc_s_bank_addr_nxt_a_1_,
         U_dsdc_N420, U_dsdc_N419, U_dsdc_N418, U_dsdc_N417, U_dsdc_N416,
         U_dsdc_N415, U_dsdc_N414, U_dsdc_N413, U_dsdc_N412, U_dsdc_N411,
         U_dsdc_N410, U_dsdc_N409, U_dsdc_N408, U_dsdc_N404, U_dsdc_N403,
         U_dsdc_N402, U_dsdc_N401, U_dsdc_i_dqs, U_dsdc_dqs_mask_end,
         U_dsdc_r_bm_close_all, U_dsdc_r_close_bank_addr_0_,
         U_dsdc_r_close_bank_addr_1_, U_dsdc_r_bm_close_bank_0_,
         U_dsdc_r_bm_close_bank_1_, U_dsdc_r_bm_close_bank_2_,
         U_dsdc_r_bm_close_bank_3_, U_dsdc_pre_amble_mute, U_dsdc_data_flag,
         U_dsdc_delta_delay_0_, U_dsdc_delta_delay_1_, U_dsdc_delta_delay_2_,
         U_dsdc_wrapped_pop_flag, U_dsdc_early_term_flag, U_dsdc_i_col_addr_1_,
         U_dsdc_i_col_addr_2_, U_dsdc_i_col_addr_4_, U_dsdc_i_col_addr_5_,
         U_dsdc_i_col_addr_6_, U_dsdc_i_col_addr_7_, U_dsdc_i_col_addr_8_,
         U_dsdc_i_col_addr_9_, U_dsdc_i_col_addr_11_, U_dsdc_i_col_addr_12_,
         U_dsdc_i_col_addr_13_, U_dsdc_i_col_addr_14_, U_dsdc_r_cas_latency_0_,
         U_dsdc_r_cas_latency_1_, U_dsdc_r_cas_latency_2_,
         U_dsdc_r_cas_latency_3_, U_dsdc_r_wrapped_burst,
         U_dsdc_r_burst_size_0_, U_dsdc_r_burst_size_1_,
         U_dsdc_r_burst_size_2_, U_dsdc_r_burst_size_3_,
         U_dsdc_r_burst_size_4_, U_dsdc_r_burst_size_5_, U_dsdc_r_rw,
         U_dsdc_r_col_addr_0_, U_dsdc_r_col_addr_1_, U_dsdc_r_col_addr_2_,
         U_dsdc_r_col_addr_3_, U_dsdc_r_col_addr_4_, U_dsdc_r_col_addr_5_,
         U_dsdc_r_col_addr_6_, U_dsdc_r_col_addr_7_, U_dsdc_r_col_addr_8_,
         U_dsdc_r_col_addr_9_, U_dsdc_r_col_addr_10_, U_dsdc_r_col_addr_11_,
         U_dsdc_r_col_addr_12_, U_dsdc_r_col_addr_13_, U_dsdc_r_col_addr_14_,
         U_dsdc_r_row_addr_0_, U_dsdc_r_row_addr_1_, U_dsdc_r_row_addr_2_,
         U_dsdc_r_row_addr_3_, U_dsdc_r_row_addr_4_, U_dsdc_r_row_addr_5_,
         U_dsdc_r_row_addr_6_, U_dsdc_r_row_addr_7_, U_dsdc_r_row_addr_8_,
         U_dsdc_r_row_addr_9_, U_dsdc_r_row_addr_10_, U_dsdc_r_row_addr_11_,
         U_dsdc_r_row_addr_12_, U_dsdc_r_row_addr_13_, U_dsdc_r_row_addr_14_,
         U_dsdc_r_row_addr_15_, U_dsdc_r_bank_addr_0_, U_dsdc_r_bank_addr_1_,
         U_dsdc_r_chip_slct_0_, U_dsdc_data_cnt_0_, U_dsdc_data_cnt_1_,
         U_dsdc_data_cnt_2_, U_dsdc_data_cnt_3_, U_dsdc_data_cnt_4_,
         U_dsdc_data_cnt_5_, U_dsdc_cas_cnt_1_, U_dsdc_cas_cnt_2_,
         U_dsdc_cas_cnt_3_, U_dsdc_cas_cnt_4_, U_dsdc_cas_cnt_5_,
         U_dsdc_row_cnt_0_, U_dsdc_row_cnt_1_, U_dsdc_row_cnt_2_,
         U_dsdc_row_cnt_3_, U_dsdc_row_cnt_4_, U_dsdc_row_cnt_5_,
         U_dsdc_row_cnt_6_, U_dsdc_row_cnt_7_, U_dsdc_row_cnt_8_,
         U_dsdc_row_cnt_9_, U_dsdc_row_cnt_10_, U_dsdc_row_cnt_11_,
         U_dsdc_row_cnt_12_, U_dsdc_row_cnt_13_, U_dsdc_row_cnt_14_,
         U_dsdc_row_cnt_15_, U_dsdc_num_init_ref_cnt_0_,
         U_dsdc_num_init_ref_cnt_1_, U_dsdc_num_init_ref_cnt_2_,
         U_dsdc_num_init_ref_cnt_3_, U_dsdc_wtr_cnt_0_, U_dsdc_wtr_cnt_2_,
         U_dsdc_wr_cnt_0_, U_dsdc_wr_cnt_2_, U_dsdc_term_cnt_0_,
         U_dsdc_term_cnt_1_, U_dsdc_term_cnt_2_, U_dsdc_term_cnt_3_,
         U_dsdc_term_cnt_4_, U_dsdc_rp_cnt2_2_, U_dsdc_rp_cnt1_0_,
         U_dsdc_rp_cnt1_1_, U_dsdc_rp_cnt1_2_, U_dsdc_rcar_cnt2_0_,
         U_dsdc_rcar_cnt2_1_, U_dsdc_rcar_cnt2_2_, U_dsdc_rcar_cnt2_3_,
         U_dsdc_rcar_cnt1_0_, U_dsdc_rcar_cnt1_1_, U_dsdc_rcar_cnt1_2_,
         U_dsdc_rcar_cnt1_3_, U_dsdc_i_dqs_d, U_dsdc_operation_cs_0_,
         U_dsdc_operation_cs_1_, U_dsdc_operation_cs_2_,
         U_dsdc_operation_cs_3_, U_dsdc_access_cs_0_, U_dsdc_access_cs_1_,
         U_dsdc_access_cs_2_, U_dsdc_access_cs_3_, U_dsdc_access_cs_4_,
         U_dsdc_s_dout_valid_nxt, U_dsdc_i_dqs_nxt, U_dsdc_n2097, U_dsdc_n2096,
         U_dsdc_n2095, U_dsdc_n2094, U_dsdc_n2093, U_ddrwr_n54, U_ddrwr_n53,
         U_ddrwr_n52, U_ddrwr_n51, U_ddrwr_n50, U_ddrwr_n49, U_ddrwr_n48,
         U_ddrwr_n47, U_ddrwr_n46, U_ddrwr_n45, U_ddrwr_n44, U_ddrwr_n43,
         U_ddrwr_n42, U_ddrwr_n41, U_ddrwr_n40, U_ddrwr_n39, U_ddrwr_n38,
         U_ddrwr_n37, U_ddrwr_n36, U_ddrwr_n35, U_ddrwr_n33, U_ddrwr_n32,
         U_ddrwr_n31, U_ddrwr_n30, U_ddrwr_n29, U_ddrwr_n28, U_ddrwr_n26,
         U_ddrwr_n27, U_ddrwr_n18, U_ddrwr_n17, U_ddrwr_n16, U_ddrwr_n15,
         U_ddrwr_n14, U_ddrwr_n13, U_ddrwr_n12, U_ddrwr_n11, U_ddrwr_n10,
         U_ddrwr_n9, U_ddrwr_n8, U_ddrwr_n7, U_ddrwr_n6, U_ddrwr_n5,
         U_ddrwr_n4, U_ddrwr_n3, U_ddrwr_n2, U_ddrwr_n1,
         U_ddrwr_hclk_2x_scan_clk, U_ddrwr_r_pre_dqm_0_, U_ddrwr_r_pre_dqm_1_,
         U_ddrwr_r_pre_dqm_2_, U_ddrwr_r_pre_dqm_3_, U_ddrwr_r_wr_data_0_,
         U_ddrwr_r_wr_data_1_, U_ddrwr_r_wr_data_2_, U_ddrwr_r_wr_data_3_,
         U_ddrwr_r_wr_data_4_, U_ddrwr_r_wr_data_5_, U_ddrwr_r_wr_data_6_,
         U_ddrwr_r_wr_data_7_, U_ddrwr_r_wr_data_8_, U_ddrwr_r_wr_data_9_,
         U_ddrwr_r_wr_data_10_, U_ddrwr_r_wr_data_11_, U_ddrwr_r_wr_data_12_,
         U_ddrwr_r_wr_data_13_, U_ddrwr_r_wr_data_14_, U_ddrwr_r_wr_data_15_,
         U_ddrwr_r_wr_data_16_, U_ddrwr_r_wr_data_17_, U_ddrwr_r_wr_data_18_,
         U_ddrwr_r_wr_data_19_, U_ddrwr_r_wr_data_20_, U_ddrwr_r_wr_data_21_,
         U_ddrwr_r_wr_data_22_, U_ddrwr_r_wr_data_23_, U_ddrwr_r_wr_data_24_,
         U_ddrwr_r_wr_data_25_, U_ddrwr_r_wr_data_26_, U_ddrwr_r_wr_data_27_,
         U_ddrwr_r_wr_data_28_, U_ddrwr_r_wr_data_29_, U_ddrwr_r_wr_data_30_,
         U_ddrwr_r_wr_data_31_, U_ddrwr_i_dqs_1_, U_ddrwr_N44,
         U_ddrwr_r_pre_dqs_hclk_2x, U_ddrwr_r_dqs, U_ddrwr_N41,
         U_ddrwr_rd_dqs_mask_d_0_, U_ddrwr_rd_dqs_mask_d_1_,
         U_ddrwr_rd_dqs_mask_d_2_, U_ddrwr_rd_dqs_mask_d_3_,
         U_ddrwr_rd_dqs_mask_d_4_, U_ddrwr_rd_dqs_mask_d_5_, U_cr_n550,
         U_cr_n549, U_cr_n548, U_cr_n547, U_cr_n546, U_cr_n545, U_cr_n544,
         U_cr_n543, U_cr_n542, U_cr_n541, U_cr_n540, U_cr_n539, U_cr_n538,
         U_cr_n537, U_cr_n536, U_cr_n535, U_cr_n534, U_cr_n533, U_cr_n532,
         U_cr_n531, U_cr_n530, U_cr_n529, U_cr_n528, U_cr_n527, U_cr_n526,
         U_cr_n525, U_cr_n524, U_cr_n523, U_cr_n522, U_cr_n521, U_cr_n520,
         U_cr_n519, U_cr_n518, U_cr_n517, U_cr_n516, U_cr_n515, U_cr_n514,
         U_cr_n513, U_cr_n512, U_cr_n511, U_cr_n510, U_cr_n509, U_cr_n508,
         U_cr_n507, U_cr_n506, U_cr_n505, U_cr_n504, U_cr_n503, U_cr_n502,
         U_cr_n501, U_cr_n500, U_cr_n499, U_cr_n498, U_cr_n497, U_cr_n496,
         U_cr_n495, U_cr_n494, U_cr_n493, U_cr_n492, U_cr_n491, U_cr_n490,
         U_cr_n489, U_cr_n488, U_cr_n487, U_cr_n486, U_cr_n485, U_cr_n484,
         U_cr_n483, U_cr_n482, U_cr_n481, U_cr_n480, U_cr_n479, U_cr_n478,
         U_cr_n477, U_cr_n476, U_cr_n475, U_cr_n474, U_cr_n473, U_cr_n472,
         U_cr_n471, U_cr_n470, U_cr_n469, U_cr_n468, U_cr_n467, U_cr_n466,
         U_cr_n465, U_cr_n464, U_cr_n463, U_cr_n462, U_cr_n461, U_cr_n460,
         U_cr_n459, U_cr_n458, U_cr_n457, U_cr_n456, U_cr_n455, U_cr_n454,
         U_cr_n453, U_cr_n452, U_cr_n451, U_cr_n450, U_cr_n449, U_cr_n448,
         U_cr_n447, U_cr_n446, U_cr_n445, U_cr_n444, U_cr_n443, U_cr_n442,
         U_cr_n441, U_cr_n440, U_cr_n439, U_cr_n438, U_cr_n437, U_cr_n436,
         U_cr_n435, U_cr_n434, U_cr_n433, U_cr_n432, U_cr_n431, U_cr_n430,
         U_cr_n429, U_cr_n428, U_cr_n427, U_cr_n426, U_cr_n425, U_cr_n424,
         U_cr_n423, U_cr_n422, U_cr_n421, U_cr_n420, U_cr_n419, U_cr_n418,
         U_cr_n417, U_cr_n416, U_cr_n415, U_cr_n414, U_cr_n413, U_cr_n412,
         U_cr_n411, U_cr_n410, U_cr_n409, U_cr_n408, U_cr_n407, U_cr_n406,
         U_cr_n405, U_cr_n404, U_cr_n403, U_cr_n402, U_cr_n401, U_cr_n400,
         U_cr_n399, U_cr_n398, U_cr_n397, U_cr_n396, U_cr_n395, U_cr_n394,
         U_cr_n393, U_cr_n392, U_cr_n391, U_cr_n390, U_cr_n389, U_cr_n388,
         U_cr_n387, U_cr_n386, U_cr_n385, U_cr_n384, U_cr_n383, U_cr_n382,
         U_cr_n381, U_cr_n380, U_cr_n379, U_cr_n378, U_cr_n377, U_cr_n376,
         U_cr_n375, U_cr_n374, U_cr_n373, U_cr_n372, U_cr_n371, U_cr_n370,
         U_cr_n369, U_cr_n368, U_cr_n367, U_cr_n366, U_cr_n365, U_cr_n364,
         U_cr_n363, U_cr_n362, U_cr_n361, U_cr_n360, U_cr_n359, U_cr_n358,
         U_cr_n357, U_cr_n356, U_cr_n355, U_cr_n354, U_cr_n353, U_cr_n352,
         U_cr_n351, U_cr_n350, U_cr_n349, U_cr_n348, U_cr_n347, U_cr_n346,
         U_cr_n345, U_cr_n344, U_cr_n343, U_cr_n342, U_cr_n341, U_cr_n340,
         U_cr_n339, U_cr_n338, U_cr_n337, U_cr_n336, U_cr_n335, U_cr_n334,
         U_cr_n333, U_cr_n332, U_cr_n331, U_cr_n330, U_cr_n329, U_cr_n328,
         U_cr_n327, U_cr_n326, U_cr_n325, U_cr_n324, U_cr_n323, U_cr_n322,
         U_cr_n321, U_cr_n320, U_cr_n319, U_cr_n318, U_cr_n317, U_cr_n316,
         U_cr_n315, U_cr_n314, U_cr_n313, U_cr_n312, U_cr_n311, U_cr_n310,
         U_cr_n309, U_cr_n308, U_cr_n307, U_cr_n306, U_cr_n305, U_cr_n304,
         U_cr_n303, U_cr_n302, U_cr_n301, U_cr_n300, U_cr_n299, U_cr_n298,
         U_cr_n297, U_cr_n296, U_cr_n295, U_cr_n294, U_cr_n293, U_cr_n292,
         U_cr_n291, U_cr_n290, U_cr_n289, U_cr_n288, U_cr_n287, U_cr_n286,
         U_cr_n285, U_cr_n284, U_cr_n283, U_cr_n282, U_cr_n281, U_cr_n280,
         U_cr_n279, U_cr_n278, U_cr_n277, U_cr_n276, U_cr_n275, U_cr_n274,
         U_cr_n273, U_cr_n272, U_cr_n271, U_cr_n270, U_cr_n269, U_cr_n268,
         U_cr_n267, U_cr_n266, U_cr_n265, U_cr_n264, U_cr_n263, U_cr_n262,
         U_cr_n261, U_cr_n260, U_cr_n259, U_cr_n258, U_cr_n257, U_cr_n256,
         U_cr_n255, U_cr_n254, U_cr_n253, U_cr_n252, U_cr_n251, U_cr_n250,
         U_cr_n249, U_cr_n248, U_cr_n247, U_cr_n246, U_cr_n245, U_cr_n244,
         U_cr_n243, U_cr_n242, U_cr_n241, U_cr_n240, U_cr_n239, U_cr_n238,
         U_cr_n237, U_cr_n236, U_cr_n235, U_cr_n234, U_cr_n233, U_cr_n232,
         U_cr_n231, U_cr_n230, U_cr_n229, U_cr_n228, U_cr_n227, U_cr_n226,
         U_cr_n225, U_cr_n224, U_cr_n223, U_cr_n222, U_cr_n221, U_cr_n220,
         U_cr_n219, U_cr_n218, U_cr_n217, U_cr_n216, U_cr_n215, U_cr_n214,
         U_cr_n213, U_cr_n212, U_cr_n211, U_cr_n210, U_cr_n209, U_cr_n208,
         U_cr_n207, U_cr_n206, U_cr_n205, U_cr_n204, U_cr_n203, U_cr_n202,
         U_cr_n201, U_cr_n200, U_cr_n199, U_cr_n198, U_cr_n197, U_cr_n196,
         U_cr_n195, U_cr_n194, U_cr_n193, U_cr_n192, U_cr_n191, U_cr_n190,
         U_cr_n189, U_cr_n188, U_cr_n187, U_cr_n186, U_cr_n185, U_cr_n184,
         U_cr_n182, U_cr_n181, U_cr_n180, U_cr_n179, U_cr_n178, U_cr_n177,
         U_cr_n176, U_cr_n175, U_cr_n174, U_cr_n171, U_cr_n170, U_cr_n169,
         U_cr_n168, U_cr_n167, U_cr_n166, U_cr_n165, U_cr_n164, U_cr_n163,
         U_cr_n162, U_cr_n161, U_cr_n160, U_cr_n159, U_cr_n158, U_cr_n157,
         U_cr_n156, U_cr_n155, U_cr_n154, U_cr_n153, U_cr_n152, U_cr_n151,
         U_cr_n150, U_cr_n149, U_cr_n148, U_cr_n147, U_cr_n146, U_cr_n145,
         U_cr_n144, U_cr_n143, U_cr_n142, U_cr_n141, U_cr_n140, U_cr_n139,
         U_cr_n138, U_cr_n137, U_cr_n136, U_cr_n135, U_cr_n134, U_cr_n133,
         U_cr_n132, U_cr_n131, U_cr_n130, U_cr_n129, U_cr_n128, U_cr_n127,
         U_cr_n126, U_cr_n125, U_cr_n124, U_cr_n123, U_cr_n122, U_cr_n121,
         U_cr_n120, U_cr_n119, U_cr_n118, U_cr_n117, U_cr_n116, U_cr_n115,
         U_cr_n114, U_cr_n113, U_cr_n112, U_cr_n111, U_cr_n110, U_cr_n109,
         U_cr_n108, U_cr_n107, U_cr_n106, U_cr_n105, U_cr_n104, U_cr_n103,
         U_cr_n102, U_cr_n101, U_cr_n100, U_cr_n97, U_cr_n72, U_cr_n71,
         U_cr_n70, U_cr_n69, U_cr_n68, U_cr_n67, U_cr_n66, U_cr_n65, U_cr_n64,
         U_cr_n63, U_cr_n62, U_cr_n61, U_cr_n60, U_cr_n59, U_cr_n58, U_cr_n57,
         U_cr_n56, U_cr_n55, U_cr_n54, U_cr_n53, U_cr_n52, U_cr_n51, U_cr_n50,
         U_cr_n49, U_cr_n48, U_cr_n47, U_cr_n46, U_cr_n45, U_cr_n44, U_cr_n43,
         U_cr_n42, U_cr_n41, U_cr_n40, U_cr_n39, U_cr_n38, U_cr_n37, U_cr_n36,
         U_cr_n35, U_cr_n34, U_cr_n33, U_cr_n32, U_cr_n31, U_cr_n30, U_cr_n29,
         U_cr_n28, U_cr_n27, U_cr_n26, U_cr_n25, U_cr_n24, U_cr_n23, U_cr_n22,
         U_cr_n21, U_cr_n20, U_cr_n19, U_cr_n18, U_cr_n17, U_cr_n16, U_cr_n13,
         U_cr_n12, U_cr_n11, U_cr_n10, U_cr_n9, U_cr_n8, U_cr_n7, U_cr_n6,
         U_cr_n5, U_cr_n4, U_cr_n3, U_cr_n2, U_cr_n1, U_cr_n99, U_cr_n98,
         U_cr_n96, U_cr_n95, U_cr_n94, U_cr_n93, U_cr_n92, U_cr_n91, U_cr_n90,
         U_cr_n89, U_cr_n88, U_cr_n87, U_cr_n86, U_cr_n85, U_cr_n84, U_cr_n83,
         U_cr_n82, U_cr_n81, U_cr_n80, U_cr_n79, U_cr_n78, U_cr_n77, U_cr_n76,
         U_cr_n75, U_cr_n74, U_cr_n73, U_cr_cr_cs_0_, U_cr_cr_cs_1_,
         U_cr_cr_cs_2_, U_cr_s_sda_d, U_cr_s_sda_d1, U_cr_N745, U_cr_N740,
         U_cr_N739, U_cr_N738, U_cr_N737, U_cr_N736, U_cr_N735, U_cr_N734,
         U_cr_N733, U_cr_N700, U_cr_N699, U_cr_N698, U_cr_N697, U_cr_N696,
         U_cr_N695, U_cr_N694, U_cr_N693, U_cr_N692, U_cr_N691, U_cr_N690,
         U_cr_N689, U_cr_N688, U_cr_N655, U_cr_N654, U_cr_N653, U_cr_N652,
         U_cr_N651, U_cr_N650, U_cr_N649, U_cr_N648, U_cr_N647, U_cr_N646,
         U_cr_N645, U_cr_N644, U_cr_N643, U_cr_N642, U_cr_N641, U_cr_N640,
         U_cr_N639, U_cr_N638, U_cr_N637, U_cr_N636, U_cr_N635, U_cr_N634,
         U_cr_N577, U_cr_N576, U_cr_N574, U_cr_N573, U_cr_N572, U_cr_N571,
         U_cr_N567, U_cr_N566, U_cr_N565, U_cr_N564, U_cr_N563, U_cr_N562,
         U_cr_N561, U_cr_N560, U_cr_N559, U_cr_N558, U_cr_N557, U_cr_N556,
         U_cr_N555, U_cr_N554, U_cr_N553, U_cr_N552, U_cr_N551, U_cr_N550,
         U_cr_N479, U_cr_N478, U_cr_N477, U_cr_N476, U_cr_N475, U_cr_N474,
         U_cr_N473, U_cr_N472, U_cr_N471, U_cr_N470, U_cr_N469, U_cr_N468,
         U_cr_N467, U_cr_N466, U_cr_N465, U_cr_N464, U_cr_N420, U_cr_N419,
         U_cr_N418, U_cr_N417, U_cr_N416, U_cr_N415, U_cr_N414, U_cr_N413,
         U_cr_N412, U_cr_N411, U_cr_N410, U_cr_N409, U_cr_N408, U_cr_N407,
         U_cr_N406, U_cr_N405, U_cr_N404, U_cr_N403, U_cr_N402, U_cr_N401,
         U_cr_N400, U_cr_N399, U_cr_N398, U_cr_N397, U_cr_N396, U_cr_N395,
         U_cr_N394, U_cr_N393, U_cr_N392, U_cr_N391, U_cr_N390, U_cr_N389,
         U_cr_N315, U_cr_N314, U_cr_N313, U_cr_N312, U_cr_N311, U_cr_N310,
         U_cr_N308, U_cr_N307, U_cr_N306, U_cr_N305, U_cr_N304, U_cr_N303,
         U_cr_N302, U_cr_N301, U_cr_N300, U_cr_N299, U_cr_N298,
         U_cr_sctlr_default_11, U_cr_stmg0r_0_, U_cr_stmg0r_1_, U_cr_stmg0r_26,
         U_cr_sctlr_12_, U_cr_sctlr_13_, U_cr_sctlr_14_, U_cr_sctlr_15_,
         U_cr_sctlr_16_, U_cr_n572, U_cr_n571, U_cr_n570, U_cr_n569, U_cr_n568,
         U_cr_n567, U_cr_n566, U_cr_n565, U_cr_n564, U_cr_n563, U_cr_n562,
         U_cr_n561, U_cr_n560, U_cr_n559, U_cr_n558, U_cr_n557, U_cr_n556,
         U_cr_n555, U_cr_n554, U_cr_n553, U_cr_n552, U_cr_n551, U_addrdec_n311,
         U_addrdec_n310, U_addrdec_n309, U_addrdec_n306, U_addrdec_n305,
         U_addrdec_n304, U_addrdec_n303, U_addrdec_n302, U_addrdec_n301,
         U_addrdec_n300, U_addrdec_n299, U_addrdec_n298, U_addrdec_n297,
         U_addrdec_n296, U_addrdec_n295, U_addrdec_n294, U_addrdec_n293,
         U_addrdec_n292, U_addrdec_n291, U_addrdec_n290, U_addrdec_n287,
         U_addrdec_n286, U_addrdec_n285, U_addrdec_n284, U_addrdec_n283,
         U_addrdec_n282, U_addrdec_n281, U_addrdec_n280, U_addrdec_n278,
         U_addrdec_n277, U_addrdec_n276, U_addrdec_n275, U_addrdec_n274,
         U_addrdec_n273, U_addrdec_n272, U_addrdec_n271, U_addrdec_n270,
         U_addrdec_n269, U_addrdec_n268, U_addrdec_n267, U_addrdec_n266,
         U_addrdec_n265, U_addrdec_n264, U_addrdec_n263, U_addrdec_n262,
         U_addrdec_n261, U_addrdec_n260, U_addrdec_n259, U_addrdec_n258,
         U_addrdec_n257, U_addrdec_n256, U_addrdec_n255, U_addrdec_n254,
         U_addrdec_n253, U_addrdec_n252, U_addrdec_n251, U_addrdec_n250,
         U_addrdec_n249, U_addrdec_n248, U_addrdec_n247, U_addrdec_n246,
         U_addrdec_n245, U_addrdec_n244, U_addrdec_n243, U_addrdec_n242,
         U_addrdec_n241, U_addrdec_n240, U_addrdec_n239, U_addrdec_n238,
         U_addrdec_n237, U_addrdec_n236, U_addrdec_n235, U_addrdec_n234,
         U_addrdec_n233, U_addrdec_n232, U_addrdec_n231, U_addrdec_n230,
         U_addrdec_n229, U_addrdec_n228, U_addrdec_n227, U_addrdec_n226,
         U_addrdec_n225, U_addrdec_n224, U_addrdec_n223, U_addrdec_n222,
         U_addrdec_n221, U_addrdec_n220, U_addrdec_n219, U_addrdec_n218,
         U_addrdec_n217, U_addrdec_n216, U_addrdec_n215, U_addrdec_n214,
         U_addrdec_n213, U_addrdec_n212, U_addrdec_n211, U_addrdec_n210,
         U_addrdec_n209, U_addrdec_n208, U_addrdec_n207, U_addrdec_n206,
         U_addrdec_n205, U_addrdec_n204, U_addrdec_n203, U_addrdec_n202,
         U_addrdec_n201, U_addrdec_n200, U_addrdec_n199, U_addrdec_n198,
         U_addrdec_n197, U_addrdec_n196, U_addrdec_n195, U_addrdec_n194,
         U_addrdec_n193, U_addrdec_n192, U_addrdec_n191, U_addrdec_n190,
         U_addrdec_n189, U_addrdec_n188, U_addrdec_n187, U_addrdec_n186,
         U_addrdec_n185, U_addrdec_n184, U_addrdec_n183, U_addrdec_n182,
         U_addrdec_n181, U_addrdec_n180, U_addrdec_n179, U_addrdec_n178,
         U_addrdec_n177, U_addrdec_n176, U_addrdec_n175, U_addrdec_n174,
         U_addrdec_n173, U_addrdec_n172, U_addrdec_n171, U_addrdec_n170,
         U_addrdec_n169, U_addrdec_n168, U_addrdec_n167, U_addrdec_n166,
         U_addrdec_n165, U_addrdec_n164, U_addrdec_n163, U_addrdec_n162,
         U_addrdec_n161, U_addrdec_n160, U_addrdec_n159, U_addrdec_n158,
         U_addrdec_n156, U_addrdec_n155, U_addrdec_n154, U_addrdec_n153,
         U_addrdec_n152, U_addrdec_n151, U_addrdec_n150, U_addrdec_n149,
         U_addrdec_n148, U_addrdec_n147, U_addrdec_n145, U_addrdec_n144,
         U_addrdec_n143, U_addrdec_n142, U_addrdec_n141, U_addrdec_n140,
         U_addrdec_n139, U_addrdec_n138, U_addrdec_n137, U_addrdec_n136,
         U_addrdec_n135, U_addrdec_n134, U_addrdec_n133, U_addrdec_n132,
         U_addrdec_n131, U_addrdec_n130, U_addrdec_n129, U_addrdec_n128,
         U_addrdec_n127, U_addrdec_n126, U_addrdec_n125, U_addrdec_n124,
         U_addrdec_n123, U_addrdec_n122, U_addrdec_n121, U_addrdec_n120,
         U_addrdec_n119, U_addrdec_n118, U_addrdec_n117, U_addrdec_n116,
         U_addrdec_n115, U_addrdec_n114, U_addrdec_n113, U_addrdec_n112,
         U_addrdec_n111, U_addrdec_n110, U_addrdec_n109, U_addrdec_n108,
         U_addrdec_n107, U_addrdec_n106, U_addrdec_n105, U_addrdec_n104,
         U_addrdec_n103, U_addrdec_n102, U_addrdec_n101, U_addrdec_n100,
         U_addrdec_n99, U_addrdec_n98, U_addrdec_n97, U_addrdec_n96,
         U_addrdec_n95, U_addrdec_n94, U_addrdec_n93, U_addrdec_n92,
         U_addrdec_n91, U_addrdec_n90, U_addrdec_n88, U_addrdec_n87,
         U_addrdec_n86, U_addrdec_n85, U_addrdec_n84, U_addrdec_n83,
         U_addrdec_n82, U_addrdec_n81, U_addrdec_n80, U_addrdec_n79,
         U_addrdec_n78, U_addrdec_n77, U_addrdec_n76, U_addrdec_n75,
         U_addrdec_n74, U_addrdec_n73, U_addrdec_n71, U_addrdec_n70,
         U_addrdec_n67, U_addrdec_n66, U_addrdec_n65, U_addrdec_n64,
         U_addrdec_n63, U_addrdec_n62, U_addrdec_n61, U_addrdec_n60,
         U_addrdec_n59, U_addrdec_n57, U_addrdec_n56, U_addrdec_n54,
         U_addrdec_n53, U_addrdec_n44, U_addrdec_n43, U_addrdec_n42,
         U_addrdec_n41, U_addrdec_n40, U_addrdec_n39, U_addrdec_n38,
         U_addrdec_n37, U_addrdec_n36, U_addrdec_n35, U_addrdec_n34,
         U_addrdec_n32, U_addrdec_n30, U_addrdec_n28, U_addrdec_n27,
         U_addrdec_n26, U_addrdec_n25, U_addrdec_n24, U_addrdec_n23,
         U_addrdec_n22, U_addrdec_n21, U_addrdec_n20, U_addrdec_n18,
         U_addrdec_n17, U_addrdec_n16, U_addrdec_n15, U_addrdec_n14,
         U_addrdec_n13, U_addrdec_n11, U_addrdec_n10, U_addrdec_n9,
         U_addrdec_n7, U_addrdec_n5, U_addrdec_n4, U_addrdec_n3, U_addrdec_n2,
         U_addrdec_n1, U_addrdec_n348, U_addrdec_n347, U_addrdec_n346,
         U_addrdec_n345, U_addrdec_n58, U_addrdec_N133, U_addrdec_N131,
         U_addrdec_N130, U_addrdec_N129, U_addrdec_N119, U_addrdec_N111,
         U_addrdec_N110, U_addrdec_N109, U_addrdec_N108, U_addrdec_N107,
         U_addrdec_bank_addr_mask_1_, U_addrdec_bcawp_0_, U_addrdec_bcawp_1_,
         U_addrdec_bcawp_2_, U_addrdec_bcawp_3_, U_addrdec_bcawp_4_,
         U_addrdec_flash_select_0_, U_addrdec_sram_select_0_,
         U_addrdec_rom_select_0_, U_refctl_n127, U_refctl_n126, U_refctl_n124,
         U_refctl_n123, U_refctl_n122, U_refctl_n121, U_refctl_n120,
         U_refctl_n119, U_refctl_n118, U_refctl_n117, U_refctl_n116,
         U_refctl_n115, U_refctl_n114, U_refctl_n113, U_refctl_n112,
         U_refctl_n111, U_refctl_n110, U_refctl_n109, U_refctl_n108,
         U_refctl_n107, U_refctl_n106, U_refctl_n105, U_refctl_n104,
         U_refctl_n103, U_refctl_n102, U_refctl_n101, U_refctl_n100,
         U_refctl_n99, U_refctl_n98, U_refctl_n97, U_refctl_n96, U_refctl_n95,
         U_refctl_n94, U_refctl_n93, U_refctl_n92, U_refctl_n91, U_refctl_n90,
         U_refctl_n89, U_refctl_n88, U_refctl_n87, U_refctl_n86, U_refctl_n85,
         U_refctl_n84, U_refctl_n83, U_refctl_n82, U_refctl_n81, U_refctl_n80,
         U_refctl_n79, U_refctl_n78, U_refctl_n77, U_refctl_n76, U_refctl_n75,
         U_refctl_n74, U_refctl_n73, U_refctl_n66, U_refctl_n65, U_refctl_n64,
         U_refctl_n63, U_refctl_n62, U_refctl_n61, U_refctl_n60, U_refctl_n59,
         U_refctl_n58, U_refctl_n57, U_refctl_n56, U_refctl_n55, U_refctl_n54,
         U_refctl_n53, U_refctl_n52, U_refctl_n51, U_refctl_n50, U_refctl_n49,
         U_refctl_n48, U_refctl_n47, U_refctl_n46, U_refctl_n45, U_refctl_n44,
         U_refctl_n43, U_refctl_n42, U_refctl_n41, U_refctl_n40, U_refctl_n39,
         U_refctl_n38, U_refctl_n37, U_refctl_n36, U_refctl_n35, U_refctl_n34,
         U_refctl_n33, U_refctl_n32, U_refctl_n30, U_refctl_n29, U_refctl_n28,
         U_refctl_n27, U_refctl_n25, U_refctl_n23, U_refctl_n22, U_refctl_n21,
         U_refctl_n20, U_refctl_n19, U_refctl_n18, U_refctl_n17, U_refctl_n16,
         U_refctl_n15, U_refctl_n14, U_refctl_n12, U_refctl_n11, U_refctl_n10,
         U_refctl_n9, U_refctl_n8, U_refctl_n7, U_refctl_n6, U_refctl_n5,
         U_refctl_n4, U_refctl_n3, U_refctl_n2, U_refctl_n1, U_refctl_N31,
         U_refctl_N30, U_refctl_N29, U_refctl_N28, U_refctl_N27, U_refctl_N26,
         U_refctl_N25, U_refctl_N24, U_refctl_N23, U_refctl_N22, U_refctl_N21,
         U_refctl_N20, U_refctl_N19, U_refctl_N18, U_refctl_N17, U_refctl_N16,
         U_refctl_next_state_0_, U_refctl_ref_req_next, U_refctl_count_next_0_,
         U_refctl_count_next_1_, U_refctl_count_next_2_,
         U_refctl_count_next_3_, U_refctl_count_next_4_,
         U_refctl_count_next_5_, U_refctl_count_next_7_,
         U_refctl_count_next_9_, U_refctl_count_next_11_,
         U_refctl_count_next_13_, U_refctl_count_next_14_,
         U_refctl_count_next_15_, U_refctl_count_0_, U_refctl_count_1_,
         U_refctl_count_2_, U_refctl_count_3_, U_refctl_count_4_,
         U_refctl_count_5_, U_refctl_count_6_, U_refctl_count_7_,
         U_refctl_count_8_, U_refctl_count_9_, U_refctl_count_10_,
         U_refctl_count_11_, U_refctl_count_12_, U_refctl_count_13_,
         U_refctl_count_14_, U_refctl_count_15_, U_refctl_current_state_0_,
         U_refctl_current_state_1_, U_dmc_n70, U_dmc_n69, U_dmc_n68, U_dmc_n67,
         U_dmc_n66, U_dmc_n65, U_dmc_n64, U_dmc_n63, U_dmc_n62, U_dmc_n61,
         U_dmc_n60, U_dmc_n59, U_dmc_n58, U_dmc_n55, U_dmc_n54, U_dmc_n53,
         U_dmc_n52, U_dmc_n51, U_dmc_n50, U_dmc_n49, U_dmc_n48, U_dmc_n47,
         U_dmc_n46, U_dmc_n45, U_dmc_n44, U_dmc_n43, U_dmc_n42, U_dmc_n41,
         U_dmc_n40, U_dmc_n39, U_dmc_n35, U_dmc_n34, U_dmc_n33, U_dmc_n32,
         U_dmc_n31, U_dmc_n30, U_dmc_n29, U_dmc_n28, U_dmc_n27, U_dmc_n26,
         U_dmc_n25, U_dmc_n24, U_dmc_n23, U_dmc_n22, U_dmc_n21, U_dmc_n20,
         U_dmc_n19, U_dmc_n18, U_dmc_n16, U_dmc_n15, U_dmc_n11, U_dmc_n10,
         U_dmc_n8, U_dmc_n7, U_dmc_n6, U_dmc_n5, U_dmc_n4, U_dmc_n3, U_dmc_n2,
         U_dmc_n1, U_dmc_n14, U_dmc_n13, U_dmc_n12, U_dmc_N24, U_dmc_N23,
         U_dmc_terminate, U_dmc_data_cnt_0_, U_dmc_data_cnt_1_,
         U_dmc_data_cnt_2_, U_dmc_data_cnt_3_, U_dmc_data_cnt_4_,
         U_dmc_data_cnt_5_, U_dmc_dmc_cs_0_, U_dmc_dmc_cs_1_, U_dmc_dmc_cs_2_,
         U_dsdc_U_minmax1_dwbb_n34, U_dsdc_U_minmax1_dwbb_n33,
         U_dsdc_U_minmax1_dwbb_n32, U_dsdc_U_minmax1_dwbb_n31,
         U_dsdc_U_minmax1_dwbb_n30, U_dsdc_U_minmax1_dwbb_n29,
         U_dsdc_U_minmax1_dwbb_n26, U_dsdc_U_minmax1_dwbb_n24,
         U_dsdc_U_minmax1_dwbb_n22, U_dsdc_U_minmax1_dwbb_n21,
         U_dsdc_U_minmax1_dwbb_n20, U_dsdc_U_minmax1_dwbb_n19,
         U_dsdc_U_minmax1_dwbb_n15, U_dsdc_U_minmax1_dwbb_n12,
         U_dsdc_U_minmax1_dwbb_n11, U_dsdc_U_minmax1_dwbb_n9,
         U_dsdc_U_minmax1_dwbb_n6, U_dsdc_U_minmax1_dwbb_n5,
         U_dsdc_U_minmax1_dwbb_n4, U_dsdc_U_minmax1_dwbb_n2,
         U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_GT_4_,
         U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_PI_1_,
         U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_0_,
         U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_1_,
         U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_,
         U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96;
  wire   [23:26] n;
  wire   [31:0] miu_rd_data_reg;
  wire   [31:0] cr_reg_data_out;
  wire   [3:0] pre_dqm;
  wire   [3:0] ad_data_mask;
  wire   [3:0] cr_row_addr_width;
  wire   [4:0] cr_num_open_banks;
  wire   [12:0] cr_exn_mode_value;
  wire   [3:0] cr_t_ras_min;
  wire   [2:0] cr_t_rcd;
  wire   [2:0] cr_t_rp;
  wire   [3:1] cr_t_rc;
  wire   [1:0] cr_t_wr;
  wire   [1:0] cr_t_wtr;
  wire   [3:0] cr_t_rcar;
  wire   [8:0] cr_t_xsr;
  wire   [15:0] cr_t_init;
  wire   [3:0] cr_num_init_ref;
  wire   [3:0] ad_cr_data_mask;
  wire   [1:0] cr_bank_addr_width;
  wire   [7:5] cr_block_size1;
  wire   [15:0] cr_t_ref;
  wire   [15:2] U_dsdc_num_row;
  wire   [14:4] U_dsdc_i_col_addr_nxt;
  wire   [5:0] U_dsdc_cas_cnt_nxt;
  wire   [2:0] U_dsdc_num_init_ref_cnt_nxt;
  wire   [4:0] U_dsdc_term_cnt_nxt;
  wire   [2:0] U_dsdc_wtr_cnt_nxt;
  wire   [2:0] U_dsdc_wr_cnt_nxt;
  wire   [2:0] U_dsdc_rp_cnt2_nxt;
  wire   [2:0] U_dsdc_rp_cnt1_nxt;
  wire   [3:0] U_dsdc_rcar_cnt2_nxt;
  wire   [3:0] U_dsdc_rcar_cnt1_nxt;
  wire   [15:13] U_dsdc_s_addr_nxt_a;
  wire   [3:0] U_dsdc_r_bm_open_bank;
  wire   [3:0] U_dsdc_r_data_mask;
  wire   [2088:2092] U_dsdc_n;
  wire   [1:0] U_ddrwr_ddr_dqm;
  wire   [15:0] U_ddrwr_ddr_wr_data;
  wire   [1:0] U_ddrwr_i2_dqs;
  wire   [31:24] U_cr_srefr;
  wire   [15:11] U_addrdec_row_addr_mask;
  wire   [5:0] U_dmc_data_cnt_nxt;

  DFFS_X2 cr_push_reg_n_reg ( .D(cr_push_n), .CK(hclk), .SN(hresetn), .Q(
        cr_push_reg_n) );
  DFFR_X1 miu_rd_data_reg_reg_31_ ( .D(cr_reg_data_out[31]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[31]) );
  DFFR_X1 miu_rd_data_reg_reg_30_ ( .D(cr_reg_data_out[30]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[30]) );
  DFFR_X1 miu_rd_data_reg_reg_29_ ( .D(cr_reg_data_out[29]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[29]) );
  DFFR_X1 miu_rd_data_reg_reg_28_ ( .D(cr_reg_data_out[28]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[28]) );
  DFFR_X1 miu_rd_data_reg_reg_27_ ( .D(cr_reg_data_out[27]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[27]) );
  DFFR_X1 miu_rd_data_reg_reg_26_ ( .D(cr_reg_data_out[26]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[26]) );
  DFFR_X1 miu_rd_data_reg_reg_25_ ( .D(cr_reg_data_out[25]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[25]) );
  DFFR_X1 miu_rd_data_reg_reg_24_ ( .D(cr_reg_data_out[24]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[24]) );
  DFFR_X1 miu_rd_data_reg_reg_23_ ( .D(cr_reg_data_out[23]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[23]) );
  DFFR_X1 miu_rd_data_reg_reg_22_ ( .D(cr_reg_data_out[22]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[22]) );
  DFFR_X1 miu_rd_data_reg_reg_21_ ( .D(cr_reg_data_out[21]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[21]) );
  DFFR_X1 miu_rd_data_reg_reg_20_ ( .D(cr_reg_data_out[20]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[20]) );
  DFFR_X1 miu_rd_data_reg_reg_19_ ( .D(cr_reg_data_out[19]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[19]) );
  DFFR_X1 miu_rd_data_reg_reg_18_ ( .D(cr_reg_data_out[18]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[18]) );
  DFFR_X1 miu_rd_data_reg_reg_17_ ( .D(cr_reg_data_out[17]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[17]) );
  DFFR_X1 miu_rd_data_reg_reg_16_ ( .D(cr_reg_data_out[16]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[16]) );
  DFFR_X1 miu_rd_data_reg_reg_15_ ( .D(cr_reg_data_out[15]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[15]) );
  DFFR_X1 miu_rd_data_reg_reg_14_ ( .D(cr_reg_data_out[14]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[14]) );
  DFFR_X1 miu_rd_data_reg_reg_13_ ( .D(cr_reg_data_out[13]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[13]) );
  DFFR_X1 miu_rd_data_reg_reg_12_ ( .D(cr_reg_data_out[12]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[12]) );
  DFFR_X1 miu_rd_data_reg_reg_11_ ( .D(cr_reg_data_out[11]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[11]) );
  DFFR_X1 miu_rd_data_reg_reg_10_ ( .D(cr_reg_data_out[10]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[10]) );
  DFFR_X1 miu_rd_data_reg_reg_9_ ( .D(cr_reg_data_out[9]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[9]) );
  DFFR_X1 miu_rd_data_reg_reg_8_ ( .D(cr_reg_data_out[8]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[8]) );
  DFFR_X1 miu_rd_data_reg_reg_7_ ( .D(cr_reg_data_out[7]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[7]) );
  DFFR_X1 miu_rd_data_reg_reg_6_ ( .D(cr_reg_data_out[6]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[6]) );
  DFFR_X1 miu_rd_data_reg_reg_5_ ( .D(cr_reg_data_out[5]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[5]) );
  DFFR_X1 miu_rd_data_reg_reg_4_ ( .D(cr_reg_data_out[4]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[4]) );
  DFFR_X1 miu_rd_data_reg_reg_3_ ( .D(cr_reg_data_out[3]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[3]) );
  DFFR_X1 miu_rd_data_reg_reg_2_ ( .D(cr_reg_data_out[2]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[2]) );
  DFFR_X1 miu_rd_data_reg_reg_1_ ( .D(cr_reg_data_out[1]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[1]) );
  DFFR_X1 miu_rd_data_reg_reg_0_ ( .D(cr_reg_data_out[0]), .CK(hclk), .RN(
        hresetn), .Q(miu_rd_data_reg[0]) );
  AOI22_X1 U3 ( .A1(s_rd_data[2]), .A2(n82), .B1(n17), .B2(miu_rd_data_reg[2]), 
        .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(miu_rd_data_out[2]) );
  AOI22_X1 U5 ( .A1(s_rd_data[8]), .A2(n82), .B1(n17), .B2(miu_rd_data_reg[8]), 
        .ZN(n2) );
  INV_X1 U6 ( .A(n2), .ZN(miu_rd_data_out[8]) );
  AOI22_X1 U7 ( .A1(s_rd_data[4]), .A2(n82), .B1(n17), .B2(miu_rd_data_reg[4]), 
        .ZN(n3) );
  INV_X1 U8 ( .A(n3), .ZN(miu_rd_data_out[4]) );
  AOI22_X1 U9 ( .A1(s_rd_data[11]), .A2(n82), .B1(n17), .B2(
        miu_rd_data_reg[11]), .ZN(n4) );
  INV_X1 U10 ( .A(n4), .ZN(miu_rd_data_out[11]) );
  AOI22_X1 U11 ( .A1(s_rd_data[14]), .A2(n82), .B1(n17), .B2(
        miu_rd_data_reg[14]), .ZN(n5) );
  INV_X1 U12 ( .A(n5), .ZN(miu_rd_data_out[14]) );
  AOI22_X1 U13 ( .A1(s_rd_data[13]), .A2(n82), .B1(n17), .B2(
        miu_rd_data_reg[13]), .ZN(n6) );
  INV_X1 U14 ( .A(n6), .ZN(miu_rd_data_out[13]) );
  AOI22_X1 U15 ( .A1(s_rd_data[15]), .A2(n82), .B1(n16), .B2(
        miu_rd_data_reg[15]), .ZN(n7) );
  INV_X1 U16 ( .A(n7), .ZN(miu_rd_data_out[15]) );
  AND3_X4 U18 ( .A1(dmc_push_n), .A2(cr_push_reg_n), .A3(n17), .ZN(miu_push_n)
         );
  INV_X8 U19 ( .A(n18), .ZN(n17) );
  NAND2_X1 U20 ( .A1(n21), .A2(hiu_mem_req), .ZN(n19) );
  INV_X1 U21 ( .A(sdram_req_i), .ZN(n21) );
  NAND2_X2 U24 ( .A1(ad_sdram_type_0_), .A2(ctl_chip_select_0_), .ZN(
        s_sel_n[0]) );
  OAI22_X2 U25 ( .A1(n21), .A2(U_cr_n39), .B1(ad_static_mem_req), .B2(n19), 
        .ZN(N28) );
  INV_X4 U26 ( .A(n44), .ZN(n14) );
  INV_X4 U27 ( .A(ctl_push_n), .ZN(n18) );
  MUX2_X2 U29 ( .A(s_rd_data[22]), .B(miu_rd_data_reg[22]), .S(n16), .Z(
        miu_rd_data_out[22]) );
  MUX2_X2 U30 ( .A(s_rd_data[30]), .B(miu_rd_data_reg[30]), .S(n17), .Z(
        miu_rd_data_out[30]) );
  MUX2_X2 U31 ( .A(s_rd_data[20]), .B(miu_rd_data_reg[20]), .S(n17), .Z(
        miu_rd_data_out[20]) );
  MUX2_X2 U32 ( .A(s_rd_data[31]), .B(miu_rd_data_reg[31]), .S(n16), .Z(
        miu_rd_data_out[31]) );
  MUX2_X2 U33 ( .A(s_rd_data[24]), .B(miu_rd_data_reg[24]), .S(n17), .Z(
        miu_rd_data_out[24]) );
  MUX2_X2 U34 ( .A(s_rd_data[28]), .B(miu_rd_data_reg[28]), .S(n16), .Z(
        miu_rd_data_out[28]) );
  MUX2_X2 U35 ( .A(s_rd_data[27]), .B(miu_rd_data_reg[27]), .S(n17), .Z(
        miu_rd_data_out[27]) );
  MUX2_X2 U36 ( .A(s_rd_data[18]), .B(miu_rd_data_reg[18]), .S(n16), .Z(
        miu_rd_data_out[18]) );
  MUX2_X2 U37 ( .A(s_rd_data[16]), .B(miu_rd_data_reg[16]), .S(n17), .Z(
        miu_rd_data_out[16]) );
  MUX2_X2 U38 ( .A(s_rd_data[23]), .B(miu_rd_data_reg[23]), .S(n16), .Z(
        miu_rd_data_out[23]) );
  MUX2_X2 U39 ( .A(s_rd_data[21]), .B(miu_rd_data_reg[21]), .S(n17), .Z(
        miu_rd_data_out[21]) );
  MUX2_X2 U40 ( .A(s_rd_data[19]), .B(miu_rd_data_reg[19]), .S(n16), .Z(
        miu_rd_data_out[19]) );
  MUX2_X2 U41 ( .A(s_rd_data[17]), .B(miu_rd_data_reg[17]), .S(n16), .Z(
        miu_rd_data_out[17]) );
  MUX2_X2 U42 ( .A(s_rd_data[25]), .B(miu_rd_data_reg[25]), .S(n17), .Z(
        miu_rd_data_out[25]) );
  MUX2_X2 U43 ( .A(s_rd_data[26]), .B(miu_rd_data_reg[26]), .S(n17), .Z(
        miu_rd_data_out[26]) );
  MUX2_X2 U44 ( .A(s_rd_data[29]), .B(miu_rd_data_reg[29]), .S(n16), .Z(
        miu_rd_data_out[29]) );
  AND3_X4 U45 ( .A1(cr_pop_n), .A2(ctl_pop_n), .A3(dmc_pop_n), .ZN(miu_pop_n)
         );
  MUX2_X2 U48 ( .A(s_rd_data[0]), .B(miu_rd_data_reg[0]), .S(n16), .Z(
        miu_rd_data_out[0]) );
  MUX2_X2 U49 ( .A(s_rd_data[10]), .B(miu_rd_data_reg[10]), .S(n16), .Z(
        miu_rd_data_out[10]) );
  MUX2_X2 U50 ( .A(s_rd_data[12]), .B(miu_rd_data_reg[12]), .S(n16), .Z(
        miu_rd_data_out[12]) );
  MUX2_X2 U51 ( .A(s_rd_data[1]), .B(miu_rd_data_reg[1]), .S(n16), .Z(
        miu_rd_data_out[1]) );
  MUX2_X2 U52 ( .A(s_rd_data[3]), .B(miu_rd_data_reg[3]), .S(n16), .Z(
        miu_rd_data_out[3]) );
  MUX2_X2 U53 ( .A(s_rd_data[5]), .B(miu_rd_data_reg[5]), .S(n16), .Z(
        miu_rd_data_out[5]) );
  MUX2_X2 U54 ( .A(s_rd_data[6]), .B(miu_rd_data_reg[6]), .S(n16), .Z(
        miu_rd_data_out[6]) );
  MUX2_X2 U55 ( .A(s_rd_data[7]), .B(miu_rd_data_reg[7]), .S(n16), .Z(
        miu_rd_data_out[7]) );
  MUX2_X2 U56 ( .A(s_rd_data[9]), .B(miu_rd_data_reg[9]), .S(n16), .Z(
        miu_rd_data_out[9]) );
  OAI211_X1 U_dsdc_U2200 ( .C1(U_dsdc_init_cnt_14_), .C2(U_dsdc_n482), .A(
        U_dsdc_init_cnt_15_), .B(U_dsdc_n1676), .ZN(U_dsdc_n1673) );
  OAI211_X1 U_dsdc_U2198 ( .C1(U_dsdc_r_wrapped_burst), .C2(U_dsdc_n166), .A(
        U_dsdc_r_burst_size_0_), .B(U_dsdc_n299), .ZN(U_dsdc_n1559) );
  NOR4_X1 U_dsdc_U2197 ( .A1(U_dsdc_operation_cs_3_), .A2(U_dsdc_n432), .A3(
        U_dsdc_n341), .A4(U_dsdc_n1506), .ZN(U_dsdc_n1479) );
  AOI21_X1 U_dsdc_U2196 ( .B1(U_dsdc_n1450), .B2(U_dsdc_n1522), .A(U_dsdc_n432), .ZN(U_dsdc_n1486) );
  XNOR2_X2 U_dsdc_U2195 ( .A(cr_t_wr[1]), .B(cr_t_wr[0]), .ZN(U_dsdc_n1306) );
  XOR2_X2 U_dsdc_U2194 ( .A(U_dsdc_n1276), .B(U_dsdc_n1278), .Z(U_dsdc_n1277)
         );
  XOR2_X2 U_dsdc_U2193 ( .A(U_dsdc_n1272), .B(U_dsdc_n1267), .Z(U_dsdc_n1271)
         );
  XNOR2_X2 U_dsdc_U2192 ( .A(cr_t_wtr[1]), .B(cr_t_wtr[0]), .ZN(U_dsdc_n1247)
         );
  MUX2_X2 U_dsdc_U2191 ( .A(cr_t_ras_min[3]), .B(U_dsdc_n1245), .S(U_dsdc_n313), .Z(U_dsdc_N4463) );
  MUX2_X2 U_dsdc_U2190 ( .A(cr_t_rc[3]), .B(U_dsdc_n1235), .S(U_dsdc_n313), 
        .Z(U_dsdc_N4476) );
  MUX2_X2 U_dsdc_U2189 ( .A(U_dsdc_n1225), .B(U_dsdc_bm_row_addr_3__0_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4477) );
  MUX2_X2 U_dsdc_U2188 ( .A(U_dsdc_n1224), .B(U_dsdc_bm_row_addr_3__1_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4478) );
  MUX2_X2 U_dsdc_U2187 ( .A(U_dsdc_n1223), .B(U_dsdc_bm_row_addr_3__2_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4479) );
  MUX2_X2 U_dsdc_U2186 ( .A(U_dsdc_n1222), .B(U_dsdc_bm_row_addr_3__3_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4480) );
  MUX2_X2 U_dsdc_U2185 ( .A(U_dsdc_n1221), .B(U_dsdc_bm_row_addr_3__4_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4481) );
  MUX2_X2 U_dsdc_U2184 ( .A(U_dsdc_n1220), .B(U_dsdc_bm_row_addr_3__5_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4482) );
  MUX2_X2 U_dsdc_U2183 ( .A(U_dsdc_n1219), .B(U_dsdc_bm_row_addr_3__6_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4483) );
  MUX2_X2 U_dsdc_U2182 ( .A(U_dsdc_n1218), .B(U_dsdc_bm_row_addr_3__13_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4490) );
  MUX2_X2 U_dsdc_U2181 ( .A(U_dsdc_n1217), .B(U_dsdc_bm_row_addr_3__14_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4491) );
  MUX2_X2 U_dsdc_U2180 ( .A(U_dsdc_n1216), .B(U_dsdc_bm_row_addr_3__15_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4492) );
  MUX2_X2 U_dsdc_U2179 ( .A(cr_t_ras_min[3]), .B(U_dsdc_n1215), .S(U_dsdc_n310), .Z(U_dsdc_N4416) );
  MUX2_X2 U_dsdc_U2178 ( .A(cr_t_rc[3]), .B(U_dsdc_n1208), .S(U_dsdc_n310), 
        .Z(U_dsdc_N4429) );
  MUX2_X2 U_dsdc_U2177 ( .A(U_dsdc_n1225), .B(U_dsdc_bm_row_addr_2__0_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4430) );
  MUX2_X2 U_dsdc_U2176 ( .A(U_dsdc_n1224), .B(U_dsdc_bm_row_addr_2__1_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4431) );
  MUX2_X2 U_dsdc_U2175 ( .A(U_dsdc_n1223), .B(U_dsdc_bm_row_addr_2__2_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4432) );
  MUX2_X2 U_dsdc_U2174 ( .A(U_dsdc_n1222), .B(U_dsdc_bm_row_addr_2__3_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4433) );
  MUX2_X2 U_dsdc_U2173 ( .A(U_dsdc_n1221), .B(U_dsdc_bm_row_addr_2__4_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4434) );
  MUX2_X2 U_dsdc_U2172 ( .A(U_dsdc_n1220), .B(U_dsdc_bm_row_addr_2__5_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4435) );
  MUX2_X2 U_dsdc_U2171 ( .A(U_dsdc_n1219), .B(U_dsdc_bm_row_addr_2__6_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4436) );
  MUX2_X2 U_dsdc_U2170 ( .A(U_dsdc_n1218), .B(U_dsdc_bm_row_addr_2__13_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4443) );
  MUX2_X2 U_dsdc_U2169 ( .A(U_dsdc_n1217), .B(U_dsdc_bm_row_addr_2__14_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4444) );
  MUX2_X2 U_dsdc_U2168 ( .A(U_dsdc_n1216), .B(U_dsdc_bm_row_addr_2__15_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4445) );
  MUX2_X2 U_dsdc_U2167 ( .A(cr_t_ras_min[3]), .B(U_dsdc_n1201), .S(U_dsdc_n620), .Z(U_dsdc_N4369) );
  MUX2_X2 U_dsdc_U2166 ( .A(cr_t_rc[3]), .B(U_dsdc_n1194), .S(U_dsdc_n620), 
        .Z(U_dsdc_N4382) );
  MUX2_X2 U_dsdc_U2165 ( .A(U_dsdc_n1225), .B(U_dsdc_bm_row_addr_1__0_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4383) );
  MUX2_X2 U_dsdc_U2164 ( .A(U_dsdc_n1224), .B(U_dsdc_bm_row_addr_1__1_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4384) );
  MUX2_X2 U_dsdc_U2163 ( .A(U_dsdc_n1223), .B(U_dsdc_bm_row_addr_1__2_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4385) );
  MUX2_X2 U_dsdc_U2162 ( .A(U_dsdc_n1222), .B(U_dsdc_bm_row_addr_1__3_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4386) );
  MUX2_X2 U_dsdc_U2161 ( .A(U_dsdc_n1221), .B(U_dsdc_bm_row_addr_1__4_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4387) );
  MUX2_X2 U_dsdc_U2160 ( .A(U_dsdc_n1220), .B(U_dsdc_bm_row_addr_1__5_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4388) );
  MUX2_X2 U_dsdc_U2159 ( .A(U_dsdc_n1219), .B(U_dsdc_bm_row_addr_1__6_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4389) );
  MUX2_X2 U_dsdc_U2158 ( .A(U_dsdc_n1218), .B(U_dsdc_bm_row_addr_1__13_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4396) );
  MUX2_X2 U_dsdc_U2157 ( .A(U_dsdc_n1217), .B(U_dsdc_bm_row_addr_1__14_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4397) );
  MUX2_X2 U_dsdc_U2156 ( .A(U_dsdc_n1216), .B(U_dsdc_bm_row_addr_1__15_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4398) );
  MUX2_X2 U_dsdc_U2155 ( .A(cr_t_ras_min[3]), .B(U_dsdc_n1187), .S(n83), .Z(
        U_dsdc_N4322) );
  MUX2_X2 U_dsdc_U2154 ( .A(cr_t_rc[3]), .B(U_dsdc_n1180), .S(n83), .Z(
        U_dsdc_N4335) );
  MUX2_X2 U_dsdc_U2152 ( .A(U_dsdc_n1225), .B(U_dsdc_bm_row_addr_0__0_), .S(
        n83), .Z(U_dsdc_N4336) );
  MUX2_X2 U_dsdc_U2151 ( .A(U_dsdc_n1224), .B(U_dsdc_bm_row_addr_0__1_), .S(
        n83), .Z(U_dsdc_N4337) );
  MUX2_X2 U_dsdc_U2150 ( .A(U_dsdc_n1223), .B(U_dsdc_bm_row_addr_0__2_), .S(
        n83), .Z(U_dsdc_N4338) );
  MUX2_X2 U_dsdc_U2149 ( .A(U_dsdc_n1222), .B(U_dsdc_bm_row_addr_0__3_), .S(
        n83), .Z(U_dsdc_N4339) );
  MUX2_X2 U_dsdc_U2148 ( .A(U_dsdc_n1221), .B(U_dsdc_bm_row_addr_0__4_), .S(
        n83), .Z(U_dsdc_N4340) );
  MUX2_X2 U_dsdc_U2147 ( .A(U_dsdc_n1220), .B(U_dsdc_bm_row_addr_0__5_), .S(
        n83), .Z(U_dsdc_N4341) );
  MUX2_X2 U_dsdc_U2146 ( .A(U_dsdc_n1219), .B(U_dsdc_bm_row_addr_0__6_), .S(
        n83), .Z(U_dsdc_N4342) );
  MUX2_X2 U_dsdc_U2145 ( .A(U_dsdc_n1218), .B(U_dsdc_bm_row_addr_0__13_), .S(
        n83), .Z(U_dsdc_N4349) );
  MUX2_X2 U_dsdc_U2144 ( .A(U_dsdc_n1217), .B(U_dsdc_bm_row_addr_0__14_), .S(
        n83), .Z(U_dsdc_N4350) );
  MUX2_X2 U_dsdc_U2143 ( .A(U_dsdc_n1216), .B(U_dsdc_bm_row_addr_0__15_), .S(
        n83), .Z(U_dsdc_N4351) );
  MUX2_X2 U_dsdc_U2142 ( .A(U_dsdc_n1164), .B(cr_t_rcd[0]), .S(U_dsdc_n1166), 
        .Z(U_dsdc_N4139) );
  MUX2_X2 U_dsdc_U2141 ( .A(U_dsdc_n1162), .B(cr_t_rcd[1]), .S(U_dsdc_n1166), 
        .Z(U_dsdc_N4140) );
  MUX2_X2 U_dsdc_U2140 ( .A(U_dsdc_n1156), .B(U_cr_n120), .S(U_dsdc_n1166), 
        .Z(U_dsdc_n1157) );
  MUX2_X2 U_dsdc_U2139 ( .A(U_dsdc_n1154), .B(U_cr_n128), .S(U_dsdc_n1166), 
        .Z(U_dsdc_n1155) );
  MUX2_X2 U_dsdc_U2137 ( .A(U_dsdc_n1151), .B(U_dsdc_bm_row_addr_3__7_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4484) );
  MUX2_X2 U_dsdc_U2136 ( .A(U_dsdc_n1151), .B(U_dsdc_bm_row_addr_2__7_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4437) );
  MUX2_X2 U_dsdc_U2135 ( .A(U_dsdc_n1151), .B(U_dsdc_bm_row_addr_1__7_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4390) );
  MUX2_X2 U_dsdc_U2134 ( .A(U_dsdc_n1151), .B(U_dsdc_bm_row_addr_0__7_), .S(
        n83), .Z(U_dsdc_N4343) );
  MUX2_X2 U_dsdc_U2133 ( .A(U_dsdc_n1149), .B(U_dsdc_bm_row_addr_3__8_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4485) );
  MUX2_X2 U_dsdc_U2132 ( .A(U_dsdc_n1149), .B(U_dsdc_bm_row_addr_2__8_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4438) );
  MUX2_X2 U_dsdc_U2131 ( .A(U_dsdc_n1149), .B(U_dsdc_bm_row_addr_1__8_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4391) );
  MUX2_X2 U_dsdc_U2130 ( .A(U_dsdc_n1149), .B(U_dsdc_bm_row_addr_0__8_), .S(
        n83), .Z(U_dsdc_N4344) );
  MUX2_X2 U_dsdc_U2129 ( .A(U_dsdc_n1148), .B(U_dsdc_bm_row_addr_3__9_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4486) );
  MUX2_X2 U_dsdc_U2128 ( .A(U_dsdc_n1148), .B(U_dsdc_bm_row_addr_2__9_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4439) );
  MUX2_X2 U_dsdc_U2127 ( .A(U_dsdc_n1148), .B(U_dsdc_bm_row_addr_1__9_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4392) );
  MUX2_X2 U_dsdc_U2126 ( .A(U_dsdc_n1148), .B(U_dsdc_bm_row_addr_0__9_), .S(
        n83), .Z(U_dsdc_N4345) );
  MUX2_X2 U_dsdc_U2125 ( .A(U_dsdc_n1146), .B(U_dsdc_bm_row_addr_3__10_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4487) );
  MUX2_X2 U_dsdc_U2124 ( .A(U_dsdc_n1146), .B(U_dsdc_bm_row_addr_2__10_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4440) );
  MUX2_X2 U_dsdc_U2123 ( .A(U_dsdc_n1146), .B(U_dsdc_bm_row_addr_1__10_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4393) );
  MUX2_X2 U_dsdc_U2122 ( .A(U_dsdc_n1146), .B(U_dsdc_bm_row_addr_0__10_), .S(
        n83), .Z(U_dsdc_N4346) );
  MUX2_X2 U_dsdc_U2121 ( .A(U_dsdc_n1145), .B(U_dsdc_bm_row_addr_3__11_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4488) );
  MUX2_X2 U_dsdc_U2120 ( .A(U_dsdc_n1145), .B(U_dsdc_bm_row_addr_2__11_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4441) );
  MUX2_X2 U_dsdc_U2119 ( .A(U_dsdc_n1145), .B(U_dsdc_bm_row_addr_1__11_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4394) );
  MUX2_X2 U_dsdc_U2118 ( .A(U_dsdc_n1145), .B(U_dsdc_bm_row_addr_0__11_), .S(
        n83), .Z(U_dsdc_N4347) );
  MUX2_X2 U_dsdc_U2117 ( .A(U_dsdc_n1143), .B(U_dsdc_bm_row_addr_3__12_), .S(
        U_dsdc_n313), .Z(U_dsdc_N4489) );
  MUX2_X2 U_dsdc_U2116 ( .A(U_dsdc_n1143), .B(U_dsdc_bm_row_addr_2__12_), .S(
        U_dsdc_n310), .Z(U_dsdc_N4442) );
  MUX2_X2 U_dsdc_U2115 ( .A(U_dsdc_n1143), .B(U_dsdc_bm_row_addr_1__12_), .S(
        U_dsdc_n620), .Z(U_dsdc_N4395) );
  MUX2_X2 U_dsdc_U2114 ( .A(U_dsdc_n1143), .B(U_dsdc_bm_row_addr_0__12_), .S(
        n83), .Z(U_dsdc_N4348) );
  XNOR2_X2 U_dsdc_U2113 ( .A(U_dsdc_n1093), .B(U_dsdc_n1091), .ZN(
        U_dsdc_cas_latency_2_) );
  INV_X4 U_dsdc_U2112 ( .A(U_dsdc_n1121), .ZN(U_dsdc_n1142) );
  MUX2_X2 U_dsdc_U2111 ( .A(U_dsdc_n1166), .B(U_dsdc_n1326), .S(
        U_dsdc_bm_num_open_bank_3_), .Z(U_dsdc_n1023) );
  MUX2_X2 U_dsdc_U2110 ( .A(U_dsdc_n1159), .B(U_dsdc_n1290), .S(
        U_dsdc_bm_num_open_bank_2_), .Z(U_dsdc_n1015) );
  MUX2_X2 U_dsdc_U2109 ( .A(U_dsdc_n1166), .B(U_dsdc_n1326), .S(
        U_dsdc_bm_num_open_bank_1_), .Z(U_dsdc_n1010) );
  MUX2_X2 U_dsdc_U2108 ( .A(U_dsdc_n1290), .B(U_dsdc_n1159), .S(U_dsdc_n340), 
        .Z(U_dsdc_n1007) );
  XNOR2_X2 U_dsdc_U2107 ( .A(ad_sdram_chip_select_0_), .B(U_dsdc_n361), .ZN(
        U_dsdc_n827) );
  XOR2_X2 U_dsdc_U2106 ( .A(U_dsdc_n697), .B(U_dsdc_i_col_addr_8_), .Z(
        U_dsdc_n1401) );
  XNOR2_X2 U_dsdc_U2105 ( .A(U_dsdc_n681), .B(U_dsdc_i_col_addr_6_), .ZN(
        U_dsdc_n1404) );
  XOR2_X2 U_dsdc_U2104 ( .A(U_dsdc_n699), .B(U_dsdc_i_col_addr_4_), .Z(
        U_dsdc_n1406) );
  XNOR2_X2 U_dsdc_U2103 ( .A(U_dsdc_n679), .B(U_dsdc_i_col_addr_14_), .ZN(
        U_dsdc_n1990) );
  XNOR2_X2 U_dsdc_U2102 ( .A(U_dsdc_n678), .B(U_dsdc_i_col_addr_13_), .ZN(
        U_dsdc_n1407) );
  NAND2_X2 U_dsdc_U2101 ( .A1(U_dsdc_n1418), .A2(U_dsdc_n1163), .ZN(
        U_dsdc_n1258) );
  INV_X4 U_dsdc_U2100 ( .A(U_dsdc_n2041), .ZN(U_dsdc_n1817) );
  XNOR2_X2 U_dsdc_U2099 ( .A(U_dsdc_n700), .B(U_dsdc_i_col_addr_12_), .ZN(
        U_dsdc_n1408) );
  NAND2_X2 U_dsdc_U2098 ( .A1(U_dsdc_n891), .A2(U_dsdc_n1411), .ZN(
        U_dsdc_n2013) );
  INV_X4 U_dsdc_U2097 ( .A(U_dsdc_n1413), .ZN(U_dsdc_n759) );
  INV_X4 U_dsdc_U2096 ( .A(U_dsdc_n2014), .ZN(U_dsdc_n1038) );
  INV_X4 U_dsdc_U2095 ( .A(U_dsdc_n966), .ZN(U_dsdc_n964) );
  NAND2_X2 U_dsdc_U2094 ( .A1(U_dsdc_n1979), .A2(U_dsdc_n1978), .ZN(
        U_dsdc_n2008) );
  NOR2_X2 U_dsdc_U2093 ( .A1(U_dsdc_n1577), .A2(U_dsdc_n1574), .ZN(
        U_dsdc_n1800) );
  NOR2_X4 U_dsdc_U2092 ( .A1(debug_ad_bank_addr[1]), .A2(U_dsdc_n1127), .ZN(
        U_dsdc_n604) );
  OAI21_X1 U_dsdc_U2091 ( .B1(U_dsdc_n1326), .B2(U_dsdc_n1166), .A(U_dsdc_n340), .ZN(U_dsdc_n1005) );
  AOI221_X2 U_dsdc_U2090 ( .B1(U_dsdc_n2066), .B2(U_dsdc_n2059), .C1(U_cr_n39), 
        .C2(U_dsdc_n2059), .A(U_dsdc_n1478), .ZN(U_dsdc_n1576) );
  NAND4_X1 U_dsdc_U2089 ( .A1(U_dsdc_n820), .A2(U_dsdc_n914), .A3(U_dsdc_n1483), .A4(U_dsdc_n825), .ZN(U_dsdc_n850) );
  AOI222_X1 U_dsdc_U2088 ( .A1(U_dsdc_RSOP_1683_C2_CONTROL1), .A2(
        U_dsdc_data_cnt_3_), .B1(U_dsdc_n751), .B2(U_dsdc_r_burst_size_3_), 
        .C1(U_dsdc_n983), .C2(hiu_burst_size[3]), .ZN(U_dsdc_n749) );
  AOI222_X1 U_dsdc_U2087 ( .A1(U_dsdc_RSOP_1683_C2_CONTROL1), .A2(
        U_dsdc_data_cnt_5_), .B1(U_dsdc_n751), .B2(U_dsdc_r_burst_size_5_), 
        .C1(U_dsdc_n983), .C2(hiu_burst_size[5]), .ZN(U_dsdc_n747) );
  OAI211_X1 U_dsdc_U2086 ( .C1(U_dsdc_n1300), .C2(U_dsdc_n1558), .A(
        U_dsdc_n1415), .B(U_dsdc_n354), .ZN(U_dsdc_n859) );
  AOI21_X1 U_dsdc_U2085 ( .B1(U_dsdc_n1312), .B2(U_dsdc_n1558), .A(U_dsdc_n181), .ZN(U_dsdc_n1316) );
  INV_X4 U_dsdc_U2084 ( .A(U_dsdc_n1112), .ZN(U_dsdc_n1388) );
  XNOR2_X2 U_dsdc_U2083 ( .A(U_dsdc_n565), .B(debug_ad_row_addr[2]), .ZN(
        U_dsdc_n566) );
  XNOR2_X2 U_dsdc_U2082 ( .A(debug_ad_row_addr[0]), .B(U_dsdc_n561), .ZN(
        U_dsdc_n567) );
  XNOR2_X2 U_dsdc_U2081 ( .A(U_dsdc_n557), .B(debug_ad_row_addr[4]), .ZN(
        U_dsdc_n568) );
  XNOR2_X2 U_dsdc_U2080 ( .A(U_dsdc_n548), .B(debug_ad_row_addr[14]), .ZN(
        U_dsdc_n549) );
  XNOR2_X2 U_dsdc_U2079 ( .A(U_dsdc_n546), .B(debug_ad_row_addr[10]), .ZN(
        U_dsdc_n550) );
  XNOR2_X2 U_dsdc_U2078 ( .A(U_dsdc_n519), .B(U_addrdec_n241), .ZN(U_dsdc_n539) );
  XNOR2_X2 U_dsdc_U2077 ( .A(U_dsdc_n510), .B(debug_ad_row_addr[8]), .ZN(
        U_dsdc_n511) );
  XNOR2_X2 U_dsdc_U2076 ( .A(U_dsdc_n504), .B(debug_ad_row_addr[6]), .ZN(
        U_dsdc_n512) );
  OR2_X4 U_dsdc_U2075 ( .A1(U_dsdc_n1660), .A2(U_dsdc_n1661), .ZN(U_dsdc_n399)
         );
  AND2_X4 U_dsdc_U2074 ( .A1(U_dsdc_n1425), .A2(U_dsdc_n166), .ZN(U_dsdc_n360)
         );
  OR2_X4 U_dsdc_U2073 ( .A1(U_dsdc_n1658), .A2(U_dsdc_n1655), .ZN(U_dsdc_n346)
         );
  OR2_X4 U_dsdc_U2072 ( .A1(U_dsdc_n1660), .A2(U_dsdc_n1655), .ZN(U_dsdc_n345)
         );
  AND2_X4 U_dsdc_U2071 ( .A1(U_dsdc_n159), .A2(U_dsdc_bm_row_addr_2__2_), .ZN(
        U_dsdc_n330) );
  AND2_X4 U_dsdc_U2070 ( .A1(U_dsdc_n998), .A2(U_dsdc_bm_row_addr_0__8_), .ZN(
        U_dsdc_n314) );
  AND2_X4 U_dsdc_U2069 ( .A1(U_dsdc_n998), .A2(U_dsdc_bm_row_addr_0__10_), 
        .ZN(U_dsdc_n312) );
  AND2_X4 U_dsdc_U2067 ( .A1(U_dsdc_n1415), .A2(U_dsdc_n703), .ZN(U_dsdc_n305)
         );
  NAND2_X2 U_dsdc_U2066 ( .A1(debug_ad_bank_addr[1]), .A2(U_dsdc_n1127), .ZN(
        U_dsdc_n599) );
  AND2_X4 U_dsdc_U2064 ( .A1(U_dsdc_n725), .A2(U_dsdc_n1258), .ZN(U_dsdc_n184)
         );
  INV_X4 U_dsdc_U2062 ( .A(U_dsdc_n1546), .ZN(U_dsdc_n983) );
  AND3_X4 U_dsdc_U2061 ( .A1(U_dsdc_n791), .A2(U_dsdc_n790), .A3(U_dsdc_n789), 
        .ZN(U_dsdc_n810) );
  AND3_X4 U_dsdc_U2060 ( .A1(U_dsdc_n788), .A2(U_dsdc_n787), .A3(U_dsdc_n786), 
        .ZN(U_dsdc_n802) );
  AND3_X4 U_dsdc_U2059 ( .A1(U_dsdc_n794), .A2(U_dsdc_n793), .A3(U_dsdc_n792), 
        .ZN(U_dsdc_n808) );
  AND3_X4 U_dsdc_U2058 ( .A1(U_dsdc_n784), .A2(U_dsdc_n783), .A3(U_dsdc_n782), 
        .ZN(U_dsdc_n805) );
  NOR2_X2 U_dsdc_U2057 ( .A1(U_dsdc_n1447), .A2(U_dsdc_n354), .ZN(U_dsdc_n1980) );
  NOR2_X2 U_dsdc_U2056 ( .A1(U_dsdc_n184), .A2(U_dsdc_n166), .ZN(U_dsdc_n1364)
         );
  AND2_X4 U_dsdc_U2055 ( .A1(U_dsdc_n292), .A2(U_dsdc_r_close_bank_addr_1_), 
        .ZN(U_dsdc_n1840) );
  INV_X4 U_dsdc_U2054 ( .A(U_dsdc_n1411), .ZN(U_dsdc_n1309) );
  NOR2_X2 U_dsdc_U2053 ( .A1(U_dsdc_n712), .A2(U_dsdc_n667), .ZN(U_dsdc_n1425)
         );
  INV_X1 U_dsdc_U2052 ( .A(U_dsdc_n663), .ZN(U_dsdc_n1561) );
  NOR2_X1 U_dsdc_U2051 ( .A1(U_dsdc_n1427), .A2(U_dsdc_n167), .ZN(U_dsdc_n691)
         );
  NOR2_X1 U_dsdc_U2050 ( .A1(U_dsdc_n692), .A2(U_dsdc_n355), .ZN(U_dsdc_n866)
         );
  AND4_X4 U_dsdc_U2049 ( .A1(U_dsdc_n885), .A2(sdram_req_i), .A3(U_dsdc_n988), 
        .A4(U_dsdc_n1438), .ZN(U_dsdc_n886) );
  NOR2_X2 U_dsdc_U2048 ( .A1(U_dsdc_n880), .A2(U_dsdc_n165), .ZN(U_dsdc_n1299)
         );
  NOR2_X2 U_dsdc_U2047 ( .A1(U_dsdc_n1455), .A2(U_dsdc_n1521), .ZN(
        U_dsdc_n1499) );
  NOR3_X2 U_dsdc_U2046 ( .A1(U_dsdc_rcar_cnt1_2_), .A2(U_dsdc_rcar_cnt1_1_), 
        .A3(U_dsdc_rcar_cnt1_0_), .ZN(U_dsdc_n1584) );
  NOR3_X2 U_dsdc_U2045 ( .A1(U_dsdc_xsr_cnt_8_), .A2(U_dsdc_xsr_cnt_7_), .A3(
        U_dsdc_n1727), .ZN(U_dsdc_n1728) );
  NAND2_X1 U_dsdc_U2043 ( .A1(U_dsdc_n1296), .A2(U_dsdc_access_cs_0_), .ZN(
        U_dsdc_n867) );
  INV_X4 U_dsdc_U2042 ( .A(U_dsdc_n1577), .ZN(U_dsdc_n2063) );
  AND3_X4 U_dsdc_U2041 ( .A1(U_dsdc_n1728), .A2(U_dsdc_n1430), .A3(
        U_dsdc_n1489), .ZN(ctl_init_done) );
  NAND3_X1 U_dsdc_U2039 ( .A1(U_dsdc_n1427), .A2(U_dsdc_access_cs_4_), .A3(
        U_dsdc_n170), .ZN(U_dsdc_n653) );
  AOI22_X1 U_dsdc_U2038 ( .A1(U_dsdc_n1424), .A2(U_dsdc_n1425), .B1(
        U_dsdc_n1412), .B2(U_dsdc_n165), .ZN(U_dsdc_n729) );
  XOR2_X2 U_dsdc_U2037 ( .A(U_dsdc_N4241), .B(U_dsdc_n612), .Z(
        U_dsdc_num_row[3]) );
  OAI21_X1 U_dsdc_U2036 ( .B1(U_dsdc_n1356), .B2(U_dsdc_access_cs_0_), .A(
        U_dsdc_n1355), .ZN(U_dsdc_n1370) );
  XNOR2_X2 U_dsdc_U2035 ( .A(cr_row_addr_width[2]), .B(U_dsdc_n1662), .ZN(
        U_dsdc_n1657) );
  XOR2_X2 U_dsdc_U2034 ( .A(U_dsdc_N4253), .B(U_dsdc_n611), .Z(
        U_dsdc_num_row[15]) );
  NAND3_X1 U_dsdc_U2033 ( .A1(hiu_rw), .A2(U_dsdc_n1284), .A3(n84), .ZN(
        U_dsdc_n969) );
  XOR2_X2 U_dsdc_U2032 ( .A(U_dsdc_N4240), .B(U_dsdc_n598), .Z(
        U_dsdc_num_row[2]) );
  XNOR2_X2 U_dsdc_U2031 ( .A(U_dsdc_n616), .B(U_dsdc_n346), .ZN(
        U_dsdc_num_row[7]) );
  XNOR2_X2 U_dsdc_U2030 ( .A(U_dsdc_n609), .B(U_dsdc_n399), .ZN(
        U_dsdc_num_row[13]) );
  XNOR2_X2 U_dsdc_U2029 ( .A(U_dsdc_n614), .B(U_dsdc_n345), .ZN(
        U_dsdc_num_row[5]) );
  XNOR2_X2 U_dsdc_U2028 ( .A(U_dsdc_N4248), .B(U_dsdc_n606), .ZN(
        U_dsdc_num_row[10]) );
  XNOR2_X2 U_dsdc_U2027 ( .A(U_dsdc_N4244), .B(U_dsdc_n615), .ZN(
        U_dsdc_num_row[6]) );
  XNOR2_X2 U_dsdc_U2026 ( .A(U_dsdc_N4246), .B(U_dsdc_n617), .ZN(
        U_dsdc_num_row[8]) );
  XNOR2_X2 U_dsdc_U2025 ( .A(U_dsdc_N4242), .B(U_dsdc_n613), .ZN(
        U_dsdc_num_row[4]) );
  XNOR2_X2 U_dsdc_U2024 ( .A(U_dsdc_N4252), .B(U_dsdc_n610), .ZN(
        U_dsdc_num_row[14]) );
  XNOR2_X2 U_dsdc_U2023 ( .A(U_dsdc_N4250), .B(U_dsdc_n608), .ZN(
        U_dsdc_num_row[12]) );
  AOI222_X1 U_dsdc_U2022 ( .A1(U_dsdc_n1268), .A2(U_dsdc_cas_cnt_5_), .B1(
        U_dsdc_r_burst_size_5_), .B2(U_dsdc_n1269), .C1(U_dsdc_n1270), .C2(
        hiu_burst_size[5]), .ZN(U_dsdc_n1267) );
  OR3_X4 U_dsdc_U2021 ( .A1(U_dsdc_n2073), .A2(U_dsdc_n1876), .A3(U_dsdc_n1875), .ZN(U_dsdc_n1881) );
  MUX2_X2 U_dsdc_U2020 ( .A(U_dsdc_n1880), .B(U_dsdc_n1879), .S(
        U_dsdc_delta_delay_1_), .Z(U_dsdc_n215) );
  NAND3_X1 U_dsdc_U2019 ( .A1(U_dsdc_n1345), .A2(ad_sdram_chip_select_0_), 
        .A3(U_dsdc_n1395), .ZN(U_dsdc_n1347) );
  NAND3_X2 U_dsdc_U2018 ( .A1(U_dsdc_n1409), .A2(U_dsdc_n1546), .A3(
        U_dsdc_n2013), .ZN(U_dsdc_n1815) );
  INV_X4 U_dsdc_U2017 ( .A(U_dsdc_n1815), .ZN(U_dsdc_n1819) );
  NOR2_X2 U_dsdc_U2016 ( .A1(U_dsdc_n1728), .A2(U_dsdc_n1754), .ZN(
        U_dsdc_n1750) );
  OR3_X4 U_dsdc_U2015 ( .A1(U_dsdc_n1425), .A2(U_dsdc_n1415), .A3(U_dsdc_n2074), .ZN(U_dsdc_n2079) );
  NOR2_X2 U_dsdc_U2014 ( .A1(U_dsdc_r_burst_size_2_), .A2(
        U_dsdc_r_burst_size_1_), .ZN(U_dsdc_n687) );
  NOR2_X2 U_dsdc_U2011 ( .A1(U_dsdc_n660), .A2(U_dsdc_n690), .ZN(U_dsdc_n1415)
         );
  NOR2_X2 U_dsdc_U2010 ( .A1(U_dsdc_cas_latency_cnt_0_), .A2(
        U_dsdc_cas_latency_cnt_1_), .ZN(U_dsdc_n1082) );
  NOR2_X2 U_dsdc_U2008 ( .A1(U_dsdc_n1165), .A2(U_dsdc_rcd_cnt_2_), .ZN(
        U_dsdc_n1163) );
  NAND2_X2 U_dsdc_U2007 ( .A1(U_dsdc_n1312), .A2(U_dsdc_r_wrapped_burst), .ZN(
        U_dsdc_n904) );
  NOR2_X2 U_dsdc_U2006 ( .A1(U_dsdc_n1297), .A2(U_dsdc_wr_cnt_2_), .ZN(
        U_dsdc_n1296) );
  NOR2_X2 U_dsdc_U2005 ( .A1(power_down), .A2(cr_do_power_down), .ZN(
        U_dsdc_n1436) );
  NOR2_X2 U_dsdc_U2004 ( .A1(U_dsdc_bm_ras_cnt_max_0_), .A2(
        U_dsdc_bm_ras_cnt_max_1_), .ZN(U_dsdc_n1153) );
  NOR2_X2 U_dsdc_U2003 ( .A1(U_dsdc_n1161), .A2(U_dsdc_bm_ras_cnt_max_3_), 
        .ZN(U_dsdc_n1437) );
  OAI21_X2 U_dsdc_U2002 ( .B1(U_dsdc_n1294), .B2(U_dsdc_n1292), .A(
        U_dsdc_n1978), .ZN(U_dsdc_n1336) );
  NOR2_X2 U_dsdc_U2001 ( .A1(U_dsdc_n1325), .A2(U_dsdc_n1336), .ZN(
        U_dsdc_n1394) );
  NAND2_X2 U_dsdc_U2000 ( .A1(U_dsdc_n964), .A2(U_dsdc_access_cs_4_), .ZN(
        U_dsdc_n725) );
  NOR2_X2 U_dsdc_U1999 ( .A1(U_dsdc_n904), .A2(U_dsdc_n1309), .ZN(U_dsdc_n1410) );
  NOR2_X2 U_dsdc_U1998 ( .A1(U_dsdc_n1309), .A2(U_dsdc_n1312), .ZN(U_dsdc_n881) );
  NAND2_X2 U_dsdc_U1997 ( .A1(U_dsdc_i_col_addr_1_), .A2(U_dsdc_n433), .ZN(
        U_dsdc_n1040) );
  NOR2_X2 U_dsdc_U1996 ( .A1(U_dsdc_n641), .A2(U_dsdc_n341), .ZN(U_dsdc_n1434)
         );
  NOR2_X2 U_dsdc_U1995 ( .A1(U_dsdc_n1258), .A2(U_dsdc_n1300), .ZN(
        U_dsdc_n1269) );
  NOR3_X2 U_dsdc_U1994 ( .A1(U_dsdc_n1270), .A2(U_dsdc_n1269), .A3(
        U_dsdc_n1268), .ZN(U_dsdc_n1340) );
  NAND3_X2 U_dsdc_U1993 ( .A1(sdram_req_i), .A2(U_dsdc_n1428), .A3(n84), .ZN(
        U_dsdc_n1975) );
  INV_X4 U_dsdc_U1992 ( .A(U_dsdc_n1975), .ZN(U_dsdc_n670) );
  NAND2_X2 U_dsdc_U1991 ( .A1(U_dsdc_n1312), .A2(U_dsdc_n328), .ZN(U_dsdc_n903) );
  NOR2_X2 U_dsdc_U1990 ( .A1(U_dsdc_cas_cnt_2_), .A2(U_dsdc_n1446), .ZN(
        U_dsdc_n663) );
  NAND2_X2 U_dsdc_U1989 ( .A1(U_dsdc_n1061), .A2(U_dsdc_n305), .ZN(U_dsdc_n991) );
  NAND2_X2 U_dsdc_U1988 ( .A1(U_dsdc_n1082), .A2(U_dsdc_n331), .ZN(
        U_dsdc_n1094) );
  NOR2_X2 U_dsdc_U1987 ( .A1(U_dsdc_n1094), .A2(U_dsdc_cas_latency_cnt_3_), 
        .ZN(U_dsdc_n1414) );
  NAND2_X2 U_dsdc_U1986 ( .A1(U_dsdc_n1344), .A2(U_dsdc_n735), .ZN(U_dsdc_n746) );
  INV_X4 U_dsdc_U1985 ( .A(U_dsdc_n1415), .ZN(U_dsdc_n2071) );
  NOR2_X2 U_dsdc_U1984 ( .A1(U_dsdc_n2071), .A2(U_dsdc_n703), .ZN(U_dsdc_n936)
         );
  NAND2_X2 U_dsdc_U1983 ( .A1(U_dsdc_n654), .A2(U_dsdc_access_cs_2_), .ZN(
        U_dsdc_n741) );
  NOR2_X2 U_dsdc_U1982 ( .A1(U_dsdc_early_term_flag), .A2(U_dsdc_data_flag), 
        .ZN(U_dsdc_n1419) );
  NAND2_X2 U_dsdc_U1981 ( .A1(U_dsdc_n738), .A2(U_dsdc_n737), .ZN(U_dsdc_n756)
         );
  NAND2_X2 U_dsdc_U1980 ( .A1(U_dsdc_n756), .A2(U_dsdc_n1079), .ZN(U_dsdc_n745) );
  INV_X4 U_dsdc_U1979 ( .A(U_dsdc_n1412), .ZN(U_dsdc_n934) );
  NAND3_X2 U_dsdc_U1976 ( .A1(U_dsdc_n746), .A2(U_dsdc_n745), .A3(U_dsdc_n744), 
        .ZN(U_dsdc_RSOP_1683_C2_CONTROL1) );
  NOR2_X2 U_dsdc_U1975 ( .A1(U_dsdc_n660), .A2(U_dsdc_n711), .ZN(U_dsdc_n1418)
         );
  NAND2_X2 U_dsdc_U1974 ( .A1(U_dsdc_n326), .A2(U_dsdc_n174), .ZN(U_dsdc_n1165) );
  NAND2_X2 U_dsdc_U1973 ( .A1(cr_s_ready_valid), .A2(U_dsdc_n1484), .ZN(
        U_dsdc_n1637) );
  INV_X4 U_dsdc_U1972 ( .A(U_dsdc_n1637), .ZN(U_dsdc_n1444) );
  NAND2_X2 U_dsdc_U1971 ( .A1(U_dsdc_n1444), .A2(U_dsdc_n1414), .ZN(
        U_dsdc_n1876) );
  NAND2_X2 U_dsdc_U1970 ( .A1(U_dsdc_n668), .A2(U_dsdc_n305), .ZN(U_dsdc_n760)
         );
  NOR2_X2 U_dsdc_U1969 ( .A1(U_dsdc_n1876), .A2(U_dsdc_n760), .ZN(
        U_dsdc_DP_OP_1642_126_2028_I4) );
  NAND4_X2 U_dsdc_U1968 ( .A1(U_dsdc_n1546), .A2(U_dsdc_n601), .A3(
        U_dsdc_n1258), .A4(U_dsdc_n755), .ZN(U_dsdc_n1380) );
  NAND2_X2 U_dsdc_U1967 ( .A1(U_dsdc_n1546), .A2(U_dsdc_n1258), .ZN(
        U_dsdc_n753) );
  NAND2_X2 U_dsdc_U1966 ( .A1(U_dsdc_n754), .A2(U_dsdc_n601), .ZN(
        U_dsdc_DP_OP_1642_126_2028_I6) );
  AOI22_X2 U_dsdc_U1965 ( .A1(U_dsdc_DP_OP_1642_126_2028_n85), .A2(
        U_dsdc_data_cnt_2_), .B1(U_dsdc_n751), .B2(U_dsdc_r_burst_size_2_), 
        .ZN(U_dsdc_n750) );
  INV_X4 U_dsdc_U1964 ( .A(U_dsdc_n752), .ZN(U_dsdc_DP_OP_1642_126_2028_I5_1_)
         );
  OAI211_X2 U_dsdc_U1963 ( .C1(U_dsdc_n754), .C2(U_dsdc_n342), .A(U_dsdc_n601), 
        .B(U_dsdc_n755), .ZN(U_dsdc_DP_OP_1642_126_2028_n86) );
  NOR2_X2 U_dsdc_U1962 ( .A1(U_dsdc_n1444), .A2(U_dsdc_data_cnt_0_), .ZN(
        U_dsdc_n1825) );
  NAND2_X2 U_dsdc_U1961 ( .A1(U_dsdc_n1825), .A2(U_dsdc_n436), .ZN(
        U_dsdc_n1823) );
  NOR2_X2 U_dsdc_U1960 ( .A1(U_dsdc_data_cnt_2_), .A2(U_dsdc_n1823), .ZN(
        U_dsdc_n1822) );
  NAND2_X2 U_dsdc_U1959 ( .A1(U_dsdc_n1822), .A2(U_dsdc_n437), .ZN(
        U_dsdc_n1820) );
  NOR2_X2 U_dsdc_U1958 ( .A1(U_dsdc_n1820), .A2(U_dsdc_data_cnt_4_), .ZN(
        U_dsdc_n762) );
  AOI21_X2 U_dsdc_U1957 ( .B1(U_dsdc_n1344), .B2(U_cr_n58), .A(U_dsdc_n756), 
        .ZN(U_dsdc_n757) );
  NOR2_X2 U_dsdc_U1956 ( .A1(U_dsdc_n757), .A2(U_dsdc_n1079), .ZN(U_dsdc_n764)
         );
  NAND2_X2 U_dsdc_U1955 ( .A1(U_dsdc_n668), .A2(U_dsdc_n1412), .ZN(U_dsdc_n758) );
  OAI22_X2 U_dsdc_U1954 ( .A1(U_dsdc_n761), .A2(U_dsdc_n760), .B1(U_dsdc_n759), 
        .B2(U_dsdc_n758), .ZN(U_dsdc_n1381) );
  INV_X4 U_dsdc_U1953 ( .A(debug_ad_row_addr[1]), .ZN(U_dsdc_n814) );
  NAND2_X2 U_dsdc_U1951 ( .A1(U_dsdc_n159), .A2(U_dsdc_bm_row_addr_2__1_), 
        .ZN(U_dsdc_n799) );
  INV_X4 U_dsdc_U1950 ( .A(U_dsdc_n813), .ZN(U_dsdc_n815) );
  NAND2_X2 U_dsdc_U1948 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__11_), 
        .ZN(U_dsdc_n791) );
  NAND2_X2 U_dsdc_U1947 ( .A1(U_dsdc_n159), .A2(U_dsdc_bm_row_addr_2__11_), 
        .ZN(U_dsdc_n790) );
  INV_X4 U_dsdc_U1946 ( .A(U_dsdc_n810), .ZN(U_dsdc_n812) );
  INV_X4 U_dsdc_U1943 ( .A(debug_ad_row_addr[9]), .ZN(U_dsdc_n803) );
  NAND2_X2 U_dsdc_U1942 ( .A1(U_dsdc_n159), .A2(U_dsdc_bm_row_addr_2__9_), 
        .ZN(U_dsdc_n787) );
  INV_X4 U_dsdc_U1941 ( .A(U_dsdc_n802), .ZN(U_dsdc_n804) );
  NOR3_X2 U_dsdc_U1940 ( .A1(U_dsdc_bm_row_addr_0__9_), .A2(U_dsdc_n803), .A3(
        U_dsdc_n804), .ZN(U_dsdc_n524) );
  NAND2_X2 U_dsdc_U1939 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__5_), 
        .ZN(U_dsdc_n794) );
  NAND2_X2 U_dsdc_U1938 ( .A1(U_dsdc_n159), .A2(U_dsdc_bm_row_addr_2__5_), 
        .ZN(U_dsdc_n793) );
  NAND2_X2 U_dsdc_U1937 ( .A1(debug_ad_row_addr[5]), .A2(U_dsdc_n808), .ZN(
        U_dsdc_n522) );
  NOR2_X2 U_dsdc_U1936 ( .A1(U_dsdc_bm_row_addr_0__5_), .A2(U_dsdc_n522), .ZN(
        U_dsdc_n523) );
  NOR2_X2 U_dsdc_U1935 ( .A1(U_dsdc_n524), .A2(U_dsdc_n523), .ZN(U_dsdc_n535)
         );
  NAND2_X2 U_dsdc_U1934 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__15_), 
        .ZN(U_dsdc_n784) );
  NAND2_X2 U_dsdc_U1933 ( .A1(U_dsdc_n159), .A2(U_dsdc_bm_row_addr_2__15_), 
        .ZN(U_dsdc_n783) );
  INV_X4 U_dsdc_U1932 ( .A(U_dsdc_n805), .ZN(U_dsdc_n807) );
  NAND2_X2 U_dsdc_U1931 ( .A1(U_dsdc_n807), .A2(U_dsdc_n806), .ZN(U_dsdc_n527)
         );
  NAND2_X2 U_dsdc_U1930 ( .A1(U_dsdc_n815), .A2(U_dsdc_n814), .ZN(U_dsdc_n526)
         );
  NAND2_X2 U_dsdc_U1929 ( .A1(U_addrdec_n231), .A2(U_dsdc_n812), .ZN(
        U_dsdc_n525) );
  NAND3_X2 U_dsdc_U1928 ( .A1(U_dsdc_n527), .A2(U_dsdc_n526), .A3(U_dsdc_n525), 
        .ZN(U_dsdc_n528) );
  INV_X4 U_dsdc_U1927 ( .A(U_dsdc_n528), .ZN(U_dsdc_n531) );
  NAND2_X2 U_dsdc_U1926 ( .A1(U_dsdc_n803), .A2(U_dsdc_n804), .ZN(U_dsdc_n530)
         );
  INV_X4 U_dsdc_U1925 ( .A(debug_ad_row_addr[5]), .ZN(U_dsdc_n1104) );
  NAND2_X2 U_dsdc_U1924 ( .A1(U_dsdc_n1104), .A2(U_dsdc_n809), .ZN(U_dsdc_n529) );
  NAND3_X2 U_dsdc_U1923 ( .A1(U_dsdc_n531), .A2(U_dsdc_n530), .A3(U_dsdc_n529), 
        .ZN(U_dsdc_n532) );
  NOR2_X2 U_dsdc_U1922 ( .A1(U_dsdc_n806), .A2(U_dsdc_n807), .ZN(U_dsdc_n533)
         );
  NOR2_X2 U_dsdc_U1921 ( .A1(U_dsdc_n532), .A2(U_dsdc_n177), .ZN(U_dsdc_n534)
         );
  NAND3_X2 U_dsdc_U1920 ( .A1(U_dsdc_n536), .A2(U_dsdc_n535), .A3(U_dsdc_n534), 
        .ZN(U_dsdc_n537) );
  NAND3_X2 U_dsdc_U1919 ( .A1(U_dsdc_n778), .A2(U_dsdc_n777), .A3(U_dsdc_n776), 
        .ZN(U_dsdc_n785) );
  NAND3_X2 U_dsdc_U1917 ( .A1(U_dsdc_n797), .A2(U_dsdc_n796), .A3(U_dsdc_n795), 
        .ZN(U_dsdc_n602) );
  INV_X4 U_dsdc_U1916 ( .A(debug_ad_row_addr[7]), .ZN(U_dsdc_n816) );
  NAND2_X2 U_dsdc_U1915 ( .A1(U_dsdc_n602), .A2(U_dsdc_n816), .ZN(U_dsdc_n540)
         );
  NAND2_X2 U_dsdc_U1914 ( .A1(U_dsdc_n516), .A2(U_dsdc_n515), .ZN(U_dsdc_n517)
         );
  AOI21_X2 U_dsdc_U1913 ( .B1(U_dsdc_n159), .B2(U_dsdc_bm_row_addr_2__12_), 
        .A(U_dsdc_n517), .ZN(U_dsdc_n519) );
  NAND3_X2 U_dsdc_U1912 ( .A1(U_dsdc_n538), .A2(U_dsdc_n540), .A3(U_dsdc_n539), 
        .ZN(U_dsdc_n541) );
  INV_X4 U_dsdc_U1911 ( .A(U_dsdc_n541), .ZN(U_dsdc_n487) );
  INV_X4 U_dsdc_U1909 ( .A(debug_ad_row_addr[3]), .ZN(U_dsdc_n801) );
  NAND2_X2 U_dsdc_U1908 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__6_), 
        .ZN(U_dsdc_n502) );
  NAND3_X2 U_dsdc_U1907 ( .A1(U_dsdc_n502), .A2(U_dsdc_n501), .A3(U_dsdc_n500), 
        .ZN(U_dsdc_n503) );
  AOI21_X2 U_dsdc_U1906 ( .B1(U_dsdc_n159), .B2(U_dsdc_bm_row_addr_2__6_), .A(
        U_dsdc_n503), .ZN(U_dsdc_n504) );
  NAND2_X2 U_dsdc_U1905 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__8_), 
        .ZN(U_dsdc_n508) );
  INV_X4 U_dsdc_U1904 ( .A(U_dsdc_n604), .ZN(U_dsdc_n600) );
  NOR2_X2 U_dsdc_U1901 ( .A1(n86), .A2(U_dsdc_n314), .ZN(U_dsdc_n507) );
  NAND2_X2 U_dsdc_U1900 ( .A1(U_dsdc_n508), .A2(U_dsdc_n507), .ZN(U_dsdc_n509)
         );
  AOI21_X2 U_dsdc_U1899 ( .B1(U_dsdc_n159), .B2(U_dsdc_bm_row_addr_2__8_), .A(
        U_dsdc_n509), .ZN(U_dsdc_n510) );
  NOR2_X2 U_dsdc_U1898 ( .A1(U_dsdc_n512), .A2(U_dsdc_n511), .ZN(U_dsdc_n513)
         );
  NAND3_X2 U_dsdc_U1897 ( .A1(U_dsdc_n332), .A2(U_dsdc_n514), .A3(U_dsdc_n513), 
        .ZN(U_dsdc_n542) );
  NAND2_X2 U_dsdc_U1896 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__4_), 
        .ZN(U_dsdc_n555) );
  NOR2_X2 U_dsdc_U1895 ( .A1(U_dsdc_n339), .A2(U_dsdc_n600), .ZN(U_dsdc_n552)
         );
  AOI21_X2 U_dsdc_U1894 ( .B1(U_dsdc_n998), .B2(U_dsdc_bm_row_addr_0__4_), .A(
        U_dsdc_n552), .ZN(U_dsdc_n553) );
  NAND2_X2 U_dsdc_U1893 ( .A1(U_dsdc_n555), .A2(U_dsdc_n553), .ZN(U_dsdc_n556)
         );
  AOI21_X2 U_dsdc_U1892 ( .B1(U_dsdc_n159), .B2(U_dsdc_bm_row_addr_2__4_), .A(
        U_dsdc_n556), .ZN(U_dsdc_n557) );
  NAND2_X2 U_dsdc_U1891 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__0_), 
        .ZN(U_dsdc_n559) );
  NAND2_X2 U_dsdc_U1889 ( .A1(U_dsdc_n559), .A2(U_dsdc_n558), .ZN(U_dsdc_n560)
         );
  NAND2_X2 U_dsdc_U1887 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__2_), 
        .ZN(U_dsdc_n563) );
  NAND2_X2 U_dsdc_U1886 ( .A1(U_dsdc_n563), .A2(U_dsdc_n562), .ZN(U_dsdc_n564)
         );
  NOR2_X2 U_dsdc_U1885 ( .A1(U_dsdc_n564), .A2(U_dsdc_n330), .ZN(U_dsdc_n565)
         );
  NOR3_X2 U_dsdc_U1884 ( .A1(U_dsdc_n568), .A2(U_dsdc_n567), .A3(U_dsdc_n566), 
        .ZN(U_dsdc_n569) );
  NOR3_X2 U_dsdc_U1883 ( .A1(U_dsdc_n798), .A2(U_dsdc_n801), .A3(
        U_dsdc_bm_row_addr_0__3_), .ZN(U_dsdc_n551) );
  NAND2_X2 U_dsdc_U1882 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__10_), 
        .ZN(U_dsdc_n544) );
  NOR2_X2 U_dsdc_U1881 ( .A1(U_dsdc_n176), .A2(U_dsdc_n312), .ZN(U_dsdc_n543)
         );
  NAND2_X2 U_dsdc_U1880 ( .A1(U_dsdc_n544), .A2(U_dsdc_n543), .ZN(U_dsdc_n545)
         );
  AOI21_X2 U_dsdc_U1879 ( .B1(U_dsdc_n159), .B2(U_dsdc_bm_row_addr_2__10_), 
        .A(U_dsdc_n545), .ZN(U_dsdc_n546) );
  NAND2_X2 U_dsdc_U1878 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__14_), 
        .ZN(U_dsdc_n547) );
  NOR3_X2 U_dsdc_U1877 ( .A1(U_dsdc_n551), .A2(U_dsdc_n550), .A3(U_dsdc_n549), 
        .ZN(U_dsdc_n570) );
  NAND2_X2 U_dsdc_U1876 ( .A1(U_dsdc_n569), .A2(U_dsdc_n570), .ZN(U_dsdc_n486)
         );
  NOR2_X2 U_dsdc_U1875 ( .A1(U_dsdc_n542), .A2(U_dsdc_n486), .ZN(U_dsdc_n485)
         );
  NAND2_X2 U_dsdc_U1874 ( .A1(U_dsdc_n808), .A2(debug_ad_row_addr[5]), .ZN(
        U_dsdc_n488) );
  NOR2_X2 U_dsdc_U1872 ( .A1(U_dsdc_n798), .A2(U_dsdc_n801), .ZN(U_dsdc_n491)
         );
  NOR3_X2 U_dsdc_U1871 ( .A1(U_dsdc_n492), .A2(U_dsdc_n318), .A3(U_dsdc_n491), 
        .ZN(U_dsdc_n498) );
  NAND2_X2 U_dsdc_U1870 ( .A1(U_dsdc_bm_row_addr_0__5_), .A2(U_dsdc_n1104), 
        .ZN(U_dsdc_n493) );
  NOR3_X2 U_dsdc_U1869 ( .A1(U_dsdc_n496), .A2(U_dsdc_n495), .A3(U_dsdc_n494), 
        .ZN(U_dsdc_n497) );
  AOI21_X2 U_dsdc_U1868 ( .B1(U_dsdc_n499), .B2(U_dsdc_n498), .A(U_dsdc_n497), 
        .ZN(U_dsdc_n571) );
  INV_X4 U_dsdc_U1867 ( .A(U_dsdc_n571), .ZN(U_dsdc_n484) );
  NAND3_X2 U_dsdc_U1866 ( .A1(U_dsdc_n487), .A2(U_dsdc_n485), .A3(U_dsdc_n484), 
        .ZN(U_dsdc_n483) );
  NOR2_X2 U_dsdc_U1865 ( .A1(U_dsdc_n884), .A2(U_dsdc_n827), .ZN(U_dsdc_n818)
         );
  NAND2_X2 U_dsdc_U1864 ( .A1(U_dsdc_n186), .A2(U_dsdc_n420), .ZN(U_dsdc_n1196) );
  NOR2_X2 U_dsdc_U1863 ( .A1(U_dsdc_n1196), .A2(U_dsdc_bm_ras_cnt_1__2_), .ZN(
        U_dsdc_n1200) );
  NAND2_X2 U_dsdc_U1862 ( .A1(U_dsdc_n1200), .A2(U_dsdc_n364), .ZN(
        U_dsdc_n1195) );
  NAND2_X2 U_dsdc_U1861 ( .A1(U_dsdc_n195), .A2(U_dsdc_n397), .ZN(U_dsdc_n1297) );
  INV_X4 U_dsdc_U1860 ( .A(U_dsdc_n1296), .ZN(U_dsdc_n1294) );
  NAND2_X2 U_dsdc_U1859 ( .A1(U_dsdc_n187), .A2(U_dsdc_n421), .ZN(U_dsdc_n1238) );
  NOR2_X2 U_dsdc_U1858 ( .A1(U_dsdc_n1238), .A2(U_dsdc_bm_ras_cnt_3__2_), .ZN(
        U_dsdc_n1244) );
  NAND2_X2 U_dsdc_U1857 ( .A1(U_dsdc_n1244), .A2(U_dsdc_n382), .ZN(
        U_dsdc_n1237) );
  NAND2_X2 U_dsdc_U1856 ( .A1(U_dsdc_n188), .A2(U_dsdc_n422), .ZN(U_dsdc_n1210) );
  NOR2_X2 U_dsdc_U1855 ( .A1(U_dsdc_n1210), .A2(U_dsdc_bm_ras_cnt_2__2_), .ZN(
        U_dsdc_n1214) );
  NAND2_X2 U_dsdc_U1854 ( .A1(U_dsdc_n1214), .A2(U_dsdc_n365), .ZN(
        U_dsdc_n1209) );
  NAND2_X2 U_dsdc_U1853 ( .A1(U_dsdc_n189), .A2(U_dsdc_n424), .ZN(U_dsdc_n1182) );
  NOR2_X2 U_dsdc_U1852 ( .A1(U_dsdc_n1182), .A2(U_dsdc_bm_ras_cnt_0__2_), .ZN(
        U_dsdc_n1186) );
  NAND2_X2 U_dsdc_U1851 ( .A1(U_dsdc_n1186), .A2(U_dsdc_n363), .ZN(
        U_dsdc_n1181) );
  NOR2_X2 U_dsdc_U1850 ( .A1(U_dsdc_n979), .A2(U_dsdc_n1546), .ZN(U_dsdc_n980)
         );
  INV_X4 U_dsdc_U1849 ( .A(U_dsdc_oldest_bank_0_), .ZN(U_dsdc_n999) );
  NOR2_X2 U_dsdc_U1848 ( .A1(U_dsdc_n999), .A2(U_dsdc_n837), .ZN(U_dsdc_n840)
         );
  NOR2_X2 U_dsdc_U1847 ( .A1(U_dsdc_oldest_bank_0_), .A2(U_dsdc_n838), .ZN(
        U_dsdc_n839) );
  OAI21_X2 U_dsdc_U1846 ( .B1(U_dsdc_n840), .B2(U_dsdc_n839), .A(U_dsdc_n1000), 
        .ZN(U_dsdc_n846) );
  NOR2_X2 U_dsdc_U1845 ( .A1(U_dsdc_n999), .A2(U_dsdc_n841), .ZN(U_dsdc_n844)
         );
  NOR2_X2 U_dsdc_U1844 ( .A1(U_dsdc_oldest_bank_0_), .A2(U_dsdc_n842), .ZN(
        U_dsdc_n843) );
  OAI21_X2 U_dsdc_U1843 ( .B1(U_dsdc_n844), .B2(U_dsdc_n843), .A(
        U_dsdc_oldest_bank_1_), .ZN(U_dsdc_n845) );
  NAND3_X2 U_dsdc_U1842 ( .A1(U_dsdc_n846), .A2(U_dsdc_n845), .A3(U_dsdc_n1296), .ZN(U_dsdc_n986) );
  INV_X4 U_dsdc_U1841 ( .A(U_dsdc_n1483), .ZN(U_dsdc_n940) );
  NOR2_X2 U_dsdc_U1840 ( .A1(U_dsdc_n827), .A2(U_dsdc_n940), .ZN(U_dsdc_n819)
         );
  NAND2_X2 U_dsdc_U1839 ( .A1(U_dsdc_n884), .A2(U_dsdc_n819), .ZN(U_dsdc_n825)
         );
  INV_X4 U_dsdc_U1838 ( .A(U_dsdc_n825), .ZN(U_dsdc_n984) );
  NOR2_X2 U_dsdc_U1837 ( .A1(U_dsdc_n986), .A2(U_dsdc_n985), .ZN(U_dsdc_n1003)
         );
  INV_X4 U_dsdc_U1836 ( .A(U_dsdc_n1003), .ZN(U_dsdc_n1004) );
  NAND3_X2 U_dsdc_U1835 ( .A1(U_dsdc_n1326), .A2(U_dsdc_n180), .A3(U_dsdc_n340), .ZN(U_dsdc_n1017) );
  NOR3_X2 U_dsdc_U1834 ( .A1(U_dsdc_n1017), .A2(U_dsdc_bm_num_open_bank_3_), 
        .A3(U_dsdc_bm_num_open_bank_2_), .ZN(U_dsdc_n1022) );
  NAND2_X2 U_dsdc_U1833 ( .A1(U_dsdc_n984), .A2(U_dsdc_n826), .ZN(U_dsdc_n975)
         );
  NAND2_X2 U_dsdc_U1832 ( .A1(U_dsdc_n975), .A2(U_dsdc_n1483), .ZN(
        U_dsdc_n1345) );
  OAI21_X2 U_dsdc_U1831 ( .B1(U_dsdc_bm_rc_cnt_0__2_), .B2(
        U_dsdc_bm_rc_cnt_0__3_), .A(U_dsdc_n998), .ZN(U_dsdc_n829) );
  NAND2_X2 U_dsdc_U1830 ( .A1(U_dsdc_n400), .A2(U_dsdc_n190), .ZN(U_dsdc_n1228) );
  NAND2_X2 U_dsdc_U1829 ( .A1(U_dsdc_n401), .A2(U_dsdc_n191), .ZN(U_dsdc_n1203) );
  AOI22_X2 U_dsdc_U1828 ( .A1(U_dsdc_n978), .A2(U_dsdc_n1228), .B1(U_dsdc_n159), .B2(U_dsdc_n1203), .ZN(U_dsdc_n834) );
  NAND2_X2 U_dsdc_U1827 ( .A1(U_dsdc_n402), .A2(U_dsdc_n192), .ZN(U_dsdc_n1175) );
  NAND2_X2 U_dsdc_U1826 ( .A1(U_dsdc_n419), .A2(U_dsdc_n193), .ZN(U_dsdc_n1189) );
  AOI22_X2 U_dsdc_U1825 ( .A1(U_dsdc_n998), .A2(U_dsdc_n1175), .B1(U_dsdc_n604), .B2(U_dsdc_n1189), .ZN(U_dsdc_n833) );
  NAND3_X2 U_dsdc_U1824 ( .A1(U_dsdc_n835), .A2(U_dsdc_n834), .A3(U_dsdc_n833), 
        .ZN(U_dsdc_n976) );
  INV_X4 U_dsdc_U1823 ( .A(U_dsdc_n827), .ZN(U_dsdc_n988) );
  NAND2_X2 U_dsdc_U1822 ( .A1(U_dsdc_n1616), .A2(U_dsdc_n430), .ZN(
        U_dsdc_n1362) );
  INV_X4 U_dsdc_U1821 ( .A(U_dsdc_n1362), .ZN(U_dsdc_n1422) );
  NOR2_X2 U_dsdc_U1820 ( .A1(U_dsdc_n658), .A2(U_dsdc_n712), .ZN(U_dsdc_n1384)
         );
  NAND3_X2 U_dsdc_U1819 ( .A1(U_dsdc_n1166), .A2(U_dsdc_bm_num_open_bank_1_), 
        .A3(U_dsdc_bm_num_open_bank_0_), .ZN(U_dsdc_n1020) );
  NOR2_X2 U_dsdc_U1818 ( .A1(U_dsdc_n1022), .A2(U_dsdc_n1021), .ZN(
        U_dsdc_n1026) );
  INV_X4 U_dsdc_U1817 ( .A(U_dsdc_n1326), .ZN(U_dsdc_n1290) );
  NAND2_X2 U_dsdc_U1816 ( .A1(U_dsdc_n1449), .A2(U_dsdc_n1465), .ZN(
        U_dsdc_n2056) );
  OAI21_X2 U_dsdc_U1815 ( .B1(U_dsdc_n1546), .B2(U_dsdc_n988), .A(U_dsdc_n1354), .ZN(U_dsdc_n990) );
  NAND2_X2 U_dsdc_U1814 ( .A1(U_dsdc_n1153), .A2(U_dsdc_n428), .ZN(
        U_dsdc_n1161) );
  NAND2_X2 U_dsdc_U1813 ( .A1(U_dsdc_n1437), .A2(U_dsdc_n1296), .ZN(
        U_dsdc_n1496) );
  NOR2_X2 U_dsdc_U1812 ( .A1(U_dsdc_n1496), .A2(U_dsdc_n940), .ZN(U_dsdc_n989)
         );
  NAND2_X2 U_dsdc_U1811 ( .A1(U_dsdc_n990), .A2(U_dsdc_n989), .ZN(U_dsdc_n1283) );
  NAND2_X2 U_dsdc_U1810 ( .A1(U_dsdc_n1416), .A2(U_dsdc_n1437), .ZN(
        U_dsdc_n1342) );
  AOI21_X2 U_dsdc_U1809 ( .B1(U_dsdc_n1386), .B2(U_dsdc_n994), .A(U_dsdc_n993), 
        .ZN(U_dsdc_n995) );
  NAND2_X2 U_dsdc_U1808 ( .A1(U_dsdc_n1283), .A2(U_dsdc_n995), .ZN(
        U_dsdc_n1325) );
  NAND2_X2 U_dsdc_U1807 ( .A1(U_dsdc_n1300), .A2(U_dsdc_n1412), .ZN(
        U_dsdc_n1064) );
  NOR2_X2 U_dsdc_U1806 ( .A1(U_dsdc_n1064), .A2(U_dsdc_n165), .ZN(U_dsdc_n715)
         );
  NAND2_X2 U_dsdc_U1805 ( .A1(U_dsdc_n1980), .A2(U_dsdc_n715), .ZN(
        U_dsdc_n1978) );
  NAND3_X2 U_dsdc_U1804 ( .A1(U_dsdc_n1290), .A2(U_dsdc_n1159), .A3(
        U_dsdc_n1394), .ZN(U_dsdc_n1006) );
  NAND2_X2 U_dsdc_U1803 ( .A1(U_dsdc_n1007), .A2(U_dsdc_n1006), .ZN(
        U_dsdc_n1011) );
  NOR2_X2 U_dsdc_U1802 ( .A1(U_dsdc_n1011), .A2(U_dsdc_n1010), .ZN(
        U_dsdc_n1016) );
  NAND2_X2 U_dsdc_U1801 ( .A1(U_dsdc_n1016), .A2(U_dsdc_n1015), .ZN(
        U_dsdc_n1024) );
  NAND2_X2 U_dsdc_U1800 ( .A1(U_dsdc_n603), .A2(U_dsdc_n1025), .ZN(U_dsdc_n297) );
  INV_X4 U_dsdc_U1799 ( .A(U_dsdc_n914), .ZN(U_dsdc_n900) );
  INV_X4 U_dsdc_U1798 ( .A(hiu_wrapped_burst), .ZN(U_dsdc_n821) );
  NOR2_X2 U_dsdc_U1797 ( .A1(hiu_burst_size[4]), .A2(U_dsdc_n1448), .ZN(
        U_dsdc_n1254) );
  NAND2_X2 U_dsdc_U1796 ( .A1(U_dsdc_n1254), .A2(hiu_burst_size[0]), .ZN(
        U_dsdc_n1557) );
  NOR2_X2 U_dsdc_U1795 ( .A1(U_dsdc_n821), .A2(U_dsdc_n1557), .ZN(U_dsdc_n1053) );
  NAND2_X2 U_dsdc_U1794 ( .A1(U_dsdc_n194), .A2(U_dsdc_n398), .ZN(U_dsdc_n1248) );
  NOR2_X2 U_dsdc_U1793 ( .A1(U_dsdc_n1248), .A2(U_dsdc_wtr_cnt_2_), .ZN(
        U_dsdc_n1284) );
  NAND2_X2 U_dsdc_U1792 ( .A1(U_dsdc_n1393), .A2(U_dsdc_n1079), .ZN(
        U_dsdc_n1090) );
  NOR2_X2 U_dsdc_U1791 ( .A1(s_cas_latency[1]), .A2(n90), .ZN(U_dsdc_n1464) );
  OAI221_X2 U_dsdc_U1790 ( .B1(n91), .B2(U_dsdc_n1461), .C1(s_cas_latency[2]), 
        .C2(U_dsdc_n1464), .A(U_dsdc_n1460), .ZN(U_dsdc_n1462) );
  NOR2_X2 U_dsdc_U1789 ( .A1(U_dsdc_n1088), .A2(U_cr_n40), .ZN(U_dsdc_n1084)
         );
  NOR2_X2 U_dsdc_U1788 ( .A1(U_dsdc_n1464), .A2(U_dsdc_n1081), .ZN(
        U_dsdc_n1092) );
  NAND4_X2 U_dsdc_U1787 ( .A1(U_dsdc_n168), .A2(U_dsdc_n356), .A3(U_dsdc_n185), 
        .A4(U_dsdc_n164), .ZN(U_dsdc_n2082) );
  NOR2_X2 U_dsdc_U1786 ( .A1(U_dsdc_r_bm_close_all), .A2(U_dsdc_n2082), .ZN(
        U_dsdc_n1826) );
  NAND2_X2 U_dsdc_U1785 ( .A1(U_dsdc_n1826), .A2(U_dsdc_n1846), .ZN(
        U_dsdc_n1942) );
  NOR3_X2 U_dsdc_U1784 ( .A1(U_dsdc_r_bm_close_bank_2_), .A2(U_dsdc_n395), 
        .A3(U_dsdc_n1942), .ZN(U_dsdc_n1867) );
  INV_X4 U_dsdc_U1783 ( .A(U_dsdc_n2082), .ZN(U_dsdc_n1941) );
  NOR2_X2 U_dsdc_U1782 ( .A1(U_dsdc_n395), .A2(U_dsdc_n1941), .ZN(U_dsdc_n1850) );
  NAND2_X2 U_dsdc_U1781 ( .A1(U_dsdc_n164), .A2(U_dsdc_n1850), .ZN(
        U_dsdc_n1860) );
  INV_X4 U_dsdc_U1780 ( .A(U_dsdc_n1867), .ZN(U_dsdc_n1859) );
  NOR2_X2 U_dsdc_U1779 ( .A1(U_dsdc_r_close_bank_addr_0_), .A2(
        U_dsdc_r_close_bank_addr_1_), .ZN(U_dsdc_n1842) );
  NAND2_X2 U_dsdc_U1778 ( .A1(U_dsdc_r_close_bank_addr_0_), .A2(
        U_dsdc_r_close_bank_addr_1_), .ZN(U_dsdc_n1841) );
  NOR2_X2 U_dsdc_U1777 ( .A1(U_dsdc_r_close_bank_addr_1_), .A2(U_dsdc_n292), 
        .ZN(U_dsdc_n1839) );
  AOI22_X2 U_dsdc_U1776 ( .A1(U_dsdc_bm_bank_age_2__3_), .A2(U_dsdc_n1840), 
        .B1(U_dsdc_n1839), .B2(U_dsdc_bm_bank_age_1__3_), .ZN(U_dsdc_n1827) );
  OAI21_X2 U_dsdc_U1775 ( .B1(U_dsdc_n1841), .B2(U_dsdc_n284), .A(U_dsdc_n1827), .ZN(U_dsdc_n1828) );
  AOI21_X2 U_dsdc_U1774 ( .B1(U_dsdc_n1842), .B2(U_dsdc_bm_bank_age_0__3_), 
        .A(U_dsdc_n1828), .ZN(U_dsdc_n1953) );
  AOI22_X2 U_dsdc_U1773 ( .A1(U_dsdc_bm_bank_age_2__1_), .A2(U_dsdc_n1840), 
        .B1(U_dsdc_n1839), .B2(U_dsdc_bm_bank_age_1__1_), .ZN(U_dsdc_n1829) );
  AOI21_X2 U_dsdc_U1772 ( .B1(U_dsdc_n1842), .B2(U_dsdc_bm_bank_age_0__1_), 
        .A(U_dsdc_n1830), .ZN(U_dsdc_n1944) );
  AOI22_X2 U_dsdc_U1771 ( .A1(U_dsdc_bm_bank_age_2__0_), .A2(U_dsdc_n1840), 
        .B1(U_dsdc_n1839), .B2(U_dsdc_bm_bank_age_1__0_), .ZN(U_dsdc_n1831) );
  AOI21_X2 U_dsdc_U1770 ( .B1(U_dsdc_n1842), .B2(U_dsdc_bm_bank_age_0__0_), 
        .A(U_dsdc_n1832), .ZN(U_dsdc_n1833) );
  NOR2_X2 U_dsdc_U1769 ( .A1(U_dsdc_n1944), .A2(U_dsdc_n1833), .ZN(
        U_dsdc_n1945) );
  NOR2_X2 U_dsdc_U1768 ( .A1(U_dsdc_n477), .A2(U_dsdc_n308), .ZN(U_dsdc_n1911)
         );
  NAND2_X2 U_dsdc_U1767 ( .A1(U_dsdc_n1944), .A2(U_dsdc_n1833), .ZN(
        U_dsdc_n1943) );
  AOI22_X2 U_dsdc_U1766 ( .A1(U_dsdc_n336), .A2(U_dsdc_n1951), .B1(U_dsdc_n178), .B2(U_dsdc_n1943), .ZN(U_dsdc_n1834) );
  OAI221_X2 U_dsdc_U1765 ( .B1(U_dsdc_bm_bank_age_2__0_), .B2(
        U_dsdc_bm_bank_age_2__1_), .C1(U_dsdc_bm_bank_age_2__0_), .C2(
        U_dsdc_n1944), .A(U_dsdc_n1834), .ZN(U_dsdc_n1836) );
  AOI22_X2 U_dsdc_U1762 ( .A1(U_dsdc_bm_bank_age_2__4_), .A2(U_dsdc_n1840), 
        .B1(U_dsdc_n1839), .B2(U_dsdc_bm_bank_age_1__4_), .ZN(U_dsdc_n1844) );
  AOI22_X2 U_dsdc_U1761 ( .A1(U_dsdc_bm_bank_age_0__4_), .A2(U_dsdc_n1842), 
        .B1(U_dsdc_n476), .B2(U_dsdc_bm_bank_age_3__4_), .ZN(U_dsdc_n1843) );
  NAND2_X2 U_dsdc_U1760 ( .A1(U_dsdc_n1844), .A2(U_dsdc_n1843), .ZN(
        U_dsdc_n1954) );
  NAND3_X2 U_dsdc_U1759 ( .A1(U_dsdc_n178), .A2(U_dsdc_n353), .A3(U_dsdc_n1849), .ZN(U_dsdc_n1856) );
  NOR3_X2 U_dsdc_U1758 ( .A1(U_dsdc_r_bm_close_all), .A2(U_dsdc_n1846), .A3(
        U_dsdc_n2082), .ZN(U_dsdc_n1961) );
  AOI21_X2 U_dsdc_U1757 ( .B1(U_dsdc_bm_bank_age_2__1_), .B2(
        U_dsdc_bm_bank_age_2__0_), .A(U_dsdc_n1860), .ZN(U_dsdc_n1855) );
  AOI211_X2 U_dsdc_U1756 ( .C1(U_dsdc_n1867), .C2(U_dsdc_n1856), .A(
        U_dsdc_n1961), .B(U_dsdc_n1855), .ZN(U_dsdc_n1858) );
  OAI221_X2 U_dsdc_U1755 ( .B1(U_dsdc_bm_bank_age_2__2_), .B2(U_dsdc_n1860), 
        .C1(U_dsdc_n336), .C2(U_dsdc_n1859), .A(U_dsdc_n1858), .ZN(
        U_dsdc_n1865) );
  AOI221_X2 U_dsdc_U1754 ( .B1(U_dsdc_n1867), .B2(U_dsdc_bm_bank_age_2__3_), 
        .C1(U_dsdc_n1866), .C2(U_dsdc_n459), .A(U_dsdc_n1865), .ZN(
        U_dsdc_n1870) );
  NOR2_X2 U_dsdc_U1753 ( .A1(U_dsdc_n336), .A2(U_dsdc_n1861), .ZN(U_dsdc_n1868) );
  OAI21_X2 U_dsdc_U1752 ( .B1(U_dsdc_n1870), .B2(U_dsdc_n350), .A(U_dsdc_n1869), .ZN(U_dsdc_n213) );
  AOI211_X2 U_dsdc_U1751 ( .C1(U_dsdc_n1024), .C2(U_dsdc_bm_num_open_bank_3_), 
        .A(U_dsdc_n1018), .B(U_dsdc_n1022), .ZN(U_dsdc_n1019) );
  INV_X4 U_dsdc_U1750 ( .A(U_dsdc_n1019), .ZN(U_dsdc_n296) );
  NOR3_X2 U_dsdc_U1749 ( .A1(U_dsdc_r_bm_close_bank_1_), .A2(U_dsdc_n383), 
        .A3(U_dsdc_n1942), .ZN(U_dsdc_n1937) );
  NOR3_X2 U_dsdc_U1748 ( .A1(U_dsdc_r_bm_open_bank[1]), .A2(U_dsdc_n1941), 
        .A3(U_dsdc_n383), .ZN(U_dsdc_n1936) );
  INV_X4 U_dsdc_U1747 ( .A(U_dsdc_n1936), .ZN(U_dsdc_n1930) );
  INV_X4 U_dsdc_U1746 ( .A(U_dsdc_n1937), .ZN(U_dsdc_n1929) );
  AOI22_X2 U_dsdc_U1745 ( .A1(U_dsdc_n335), .A2(U_dsdc_n1943), .B1(U_dsdc_n337), .B2(U_dsdc_n1951), .ZN(U_dsdc_n1912) );
  OAI221_X2 U_dsdc_U1744 ( .B1(U_dsdc_bm_bank_age_1__0_), .B2(
        U_dsdc_bm_bank_age_1__1_), .C1(U_dsdc_bm_bank_age_1__0_), .C2(
        U_dsdc_n1944), .A(U_dsdc_n1912), .ZN(U_dsdc_n1914) );
  AOI221_X2 U_dsdc_U1743 ( .B1(U_dsdc_n1945), .B2(U_dsdc_n1915), .C1(
        U_dsdc_n1914), .C2(U_dsdc_n1915), .A(U_dsdc_n1913), .ZN(U_dsdc_n1916)
         );
  AOI21_X2 U_dsdc_U1742 ( .B1(U_dsdc_bm_bank_age_1__3_), .B2(U_dsdc_n1953), 
        .A(U_dsdc_n1916), .ZN(U_dsdc_n1917) );
  NAND3_X2 U_dsdc_U1741 ( .A1(U_dsdc_n335), .A2(U_dsdc_n352), .A3(U_dsdc_n1920), .ZN(U_dsdc_n1926) );
  AOI21_X2 U_dsdc_U1740 ( .B1(U_dsdc_bm_bank_age_1__1_), .B2(
        U_dsdc_bm_bank_age_1__0_), .A(U_dsdc_n1930), .ZN(U_dsdc_n1925) );
  AOI211_X2 U_dsdc_U1739 ( .C1(U_dsdc_n1937), .C2(U_dsdc_n1926), .A(
        U_dsdc_n1961), .B(U_dsdc_n1925), .ZN(U_dsdc_n1928) );
  OAI221_X2 U_dsdc_U1738 ( .B1(U_dsdc_bm_bank_age_1__2_), .B2(U_dsdc_n1930), 
        .C1(U_dsdc_n337), .C2(U_dsdc_n1929), .A(U_dsdc_n1928), .ZN(
        U_dsdc_n1935) );
  AOI221_X2 U_dsdc_U1737 ( .B1(U_dsdc_n1937), .B2(U_dsdc_bm_bank_age_1__3_), 
        .C1(U_dsdc_n1936), .C2(U_dsdc_n460), .A(U_dsdc_n1935), .ZN(
        U_dsdc_n1940) );
  NAND3_X2 U_dsdc_U1736 ( .A1(U_dsdc_bm_bank_age_1__1_), .A2(
        U_dsdc_bm_bank_age_1__0_), .A3(U_dsdc_n1936), .ZN(U_dsdc_n1931) );
  NOR2_X2 U_dsdc_U1735 ( .A1(U_dsdc_n337), .A2(U_dsdc_n1931), .ZN(U_dsdc_n1938) );
  OAI21_X2 U_dsdc_U1734 ( .B1(U_dsdc_n1940), .B2(U_dsdc_n349), .A(U_dsdc_n1939), .ZN(U_dsdc_n227) );
  NOR2_X2 U_dsdc_U1733 ( .A1(U_dsdc_n903), .A2(U_dsdc_n1309), .ZN(U_dsdc_n879)
         );
  NAND2_X2 U_dsdc_U1732 ( .A1(U_dsdc_n682), .A2(U_dsdc_n758), .ZN(U_dsdc_n724)
         );
  NAND2_X2 U_dsdc_U1731 ( .A1(U_dsdc_n457), .A2(U_dsdc_n200), .ZN(U_dsdc_n650)
         );
  NOR2_X2 U_dsdc_U1730 ( .A1(U_dsdc_term_cnt_0_), .A2(U_dsdc_term_cnt_1_), 
        .ZN(U_dsdc_n1638) );
  INV_X4 U_dsdc_U1729 ( .A(U_dsdc_n1638), .ZN(U_dsdc_n1640) );
  NOR3_X2 U_dsdc_U1728 ( .A1(U_dsdc_n650), .A2(U_dsdc_term_cnt_3_), .A3(
        U_dsdc_n1640), .ZN(U_dsdc_n1424) );
  NAND2_X2 U_dsdc_U1727 ( .A1(U_dsdc_n171), .A2(U_dsdc_n309), .ZN(U_dsdc_n1329) );
  NOR2_X2 U_dsdc_U1726 ( .A1(U_dsdc_n1329), .A2(U_dsdc_rp_cnt2_2_), .ZN(
        U_dsdc_n1426) );
  NAND2_X2 U_dsdc_U1725 ( .A1(U_dsdc_n1424), .A2(U_dsdc_n1426), .ZN(
        U_dsdc_n1871) );
  INV_X4 U_dsdc_U1724 ( .A(U_dsdc_n1871), .ZN(U_dsdc_n1423) );
  NAND3_X2 U_dsdc_U1723 ( .A1(U_dsdc_n1423), .A2(U_dsdc_r_rw), .A3(
        U_dsdc_n1425), .ZN(U_dsdc_n1627) );
  INV_X4 U_dsdc_U1722 ( .A(U_dsdc_n1627), .ZN(U_dsdc_n722) );
  NOR2_X2 U_dsdc_U1721 ( .A1(U_dsdc_n692), .A2(U_dsdc_n690), .ZN(U_dsdc_n1293)
         );
  INV_X4 U_dsdc_U1720 ( .A(U_dsdc_n1410), .ZN(U_dsdc_n1556) );
  INV_X4 U_dsdc_U1719 ( .A(U_dsdc_n936), .ZN(U_dsdc_n673) );
  NOR2_X2 U_dsdc_U1718 ( .A1(U_dsdc_n673), .A2(U_dsdc_n904), .ZN(U_dsdc_n683)
         );
  AOI21_X2 U_dsdc_U1717 ( .B1(U_dsdc_n1060), .B2(U_dsdc_n724), .A(U_dsdc_n683), 
        .ZN(U_dsdc_n1403) );
  NAND2_X2 U_dsdc_U1716 ( .A1(U_dsdc_n736), .A2(U_dsdc_access_cs_0_), .ZN(
        U_dsdc_n1629) );
  NOR2_X2 U_dsdc_U1715 ( .A1(U_dsdc_n684), .A2(U_dsdc_n1633), .ZN(U_dsdc_n728)
         );
  AOI21_X2 U_dsdc_U1714 ( .B1(U_dsdc_n685), .B2(U_dsdc_n1423), .A(U_dsdc_n728), 
        .ZN(U_dsdc_n686) );
  NOR2_X2 U_dsdc_U1713 ( .A1(U_dsdc_n686), .A2(U_dsdc_n1419), .ZN(U_dsdc_n1625) );
  NOR3_X2 U_dsdc_U1712 ( .A1(U_dsdc_n1559), .A2(U_dsdc_n1258), .A3(U_dsdc_n688), .ZN(U_dsdc_n689) );
  AOI211_X2 U_dsdc_U1711 ( .C1(U_dsdc_n865), .C2(U_dsdc_wrapped_pop_flag), .A(
        U_dsdc_n1625), .B(U_dsdc_n689), .ZN(U_dsdc_n1560) );
  OAI221_X2 U_dsdc_U1710 ( .B1(U_dsdc_n1561), .B2(U_dsdc_n1403), .C1(
        U_dsdc_n1561), .C2(U_dsdc_n1651), .A(U_dsdc_n1560), .ZN(U_dsdc_n1562)
         );
  NOR3_X2 U_dsdc_U1709 ( .A1(U_dsdc_n1293), .A2(U_dsdc_n1563), .A3(
        U_dsdc_n1562), .ZN(U_dsdc_n726) );
  OAI211_X2 U_dsdc_U1708 ( .C1(U_dsdc_n727), .C2(U_dsdc_n181), .A(U_dsdc_n726), 
        .B(U_dsdc_n725), .ZN(ctl_burst_done) );
  NOR2_X2 U_dsdc_U1707 ( .A1(U_dsdc_n1175), .A2(U_dsdc_bm_rc_cnt_0__2_), .ZN(
        U_dsdc_n1179) );
  NOR2_X2 U_dsdc_U1706 ( .A1(U_dsdc_n1179), .A2(U_dsdc_n441), .ZN(U_dsdc_n1180) );
  AOI21_X2 U_dsdc_U1705 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[13]), .A(
        U_dsdc_n1132), .ZN(U_dsdc_n1169) );
  INV_X4 U_dsdc_U1704 ( .A(U_dsdc_n1169), .ZN(U_dsdc_n1218) );
  AOI21_X2 U_dsdc_U1703 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[3]), .A(
        U_dsdc_n1115), .ZN(U_dsdc_n1170) );
  INV_X4 U_dsdc_U1702 ( .A(U_dsdc_n1170), .ZN(U_dsdc_n1222) );
  AOI21_X2 U_dsdc_U1701 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[9]), .A(
        U_dsdc_n1073), .ZN(U_dsdc_n1147) );
  INV_X4 U_dsdc_U1700 ( .A(U_dsdc_n1147), .ZN(U_dsdc_n1148) );
  AOI21_X2 U_dsdc_U1699 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[2]), .A(
        U_dsdc_n1116), .ZN(U_dsdc_n1171) );
  INV_X4 U_dsdc_U1698 ( .A(U_dsdc_n1171), .ZN(U_dsdc_n1223) );
  NAND2_X2 U_dsdc_U1697 ( .A1(U_dsdc_n1109), .A2(U_dsdc_r_row_addr_10_), .ZN(
        U_dsdc_n1027) );
  OAI21_X2 U_dsdc_U1696 ( .B1(U_dsdc_n1112), .B2(U_dsdc_n1028), .A(
        U_dsdc_n1027), .ZN(U_dsdc_n1146) );
  NAND2_X2 U_dsdc_U1695 ( .A1(U_dsdc_n1109), .A2(U_dsdc_r_row_addr_4_), .ZN(
        U_dsdc_n1110) );
  OAI21_X2 U_dsdc_U1694 ( .B1(U_dsdc_n1112), .B2(U_dsdc_n1111), .A(
        U_dsdc_n1110), .ZN(U_dsdc_n1221) );
  AOI21_X2 U_dsdc_U1693 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[11]), .A(
        U_dsdc_n1069), .ZN(U_dsdc_n1144) );
  INV_X4 U_dsdc_U1692 ( .A(U_dsdc_n1144), .ZN(U_dsdc_n1145) );
  AOI21_X2 U_dsdc_U1691 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[1]), .A(
        U_dsdc_n1117), .ZN(U_dsdc_n1172) );
  INV_X4 U_dsdc_U1690 ( .A(U_dsdc_n1172), .ZN(U_dsdc_n1224) );
  NAND2_X2 U_dsdc_U1689 ( .A1(U_dsdc_n1109), .A2(U_dsdc_r_row_addr_8_), .ZN(
        U_dsdc_n1075) );
  OAI21_X2 U_dsdc_U1688 ( .B1(U_dsdc_n1112), .B2(U_dsdc_n1076), .A(
        U_dsdc_n1075), .ZN(U_dsdc_n1149) );
  AOI21_X2 U_dsdc_U1687 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[7]), .A(
        U_dsdc_n1095), .ZN(U_dsdc_n1150) );
  INV_X4 U_dsdc_U1686 ( .A(U_dsdc_n1150), .ZN(U_dsdc_n1151) );
  NAND2_X2 U_dsdc_U1685 ( .A1(U_dsdc_n1109), .A2(U_dsdc_r_row_addr_5_), .ZN(
        U_dsdc_n1103) );
  OAI21_X2 U_dsdc_U1684 ( .B1(U_dsdc_n1112), .B2(U_dsdc_n1104), .A(
        U_dsdc_n1103), .ZN(U_dsdc_n1220) );
  NAND2_X2 U_dsdc_U1683 ( .A1(U_dsdc_n1109), .A2(U_dsdc_r_row_addr_6_), .ZN(
        U_dsdc_n1097) );
  OAI21_X2 U_dsdc_U1682 ( .B1(U_dsdc_n1112), .B2(U_dsdc_n1098), .A(
        U_dsdc_n1097), .ZN(U_dsdc_n1219) );
  NAND2_X2 U_dsdc_U1681 ( .A1(U_dsdc_n1109), .A2(U_dsdc_r_row_addr_12_), .ZN(
        U_dsdc_n1058) );
  OAI21_X2 U_dsdc_U1680 ( .B1(U_dsdc_n1112), .B2(U_addrdec_n241), .A(
        U_dsdc_n1058), .ZN(U_dsdc_n1143) );
  AOI21_X2 U_dsdc_U1679 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[14]), .A(
        U_dsdc_n1134), .ZN(U_dsdc_n1168) );
  INV_X4 U_dsdc_U1678 ( .A(U_dsdc_n1168), .ZN(U_dsdc_n1217) );
  AOI21_X2 U_dsdc_U1677 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[0]), .A(
        U_dsdc_n1122), .ZN(U_dsdc_n1173) );
  INV_X4 U_dsdc_U1676 ( .A(U_dsdc_n1173), .ZN(U_dsdc_n1225) );
  AOI21_X2 U_dsdc_U1675 ( .B1(U_dsdc_n1388), .B2(debug_ad_row_addr[15]), .A(
        U_dsdc_n1137), .ZN(U_dsdc_n1167) );
  INV_X4 U_dsdc_U1674 ( .A(U_dsdc_n1167), .ZN(U_dsdc_n1216) );
  NOR2_X2 U_dsdc_U1673 ( .A1(U_dsdc_n1228), .A2(U_dsdc_bm_rc_cnt_3__2_), .ZN(
        U_dsdc_n1234) );
  NOR2_X2 U_dsdc_U1672 ( .A1(U_dsdc_n1234), .A2(U_dsdc_n442), .ZN(U_dsdc_n1235) );
  OAI21_X2 U_dsdc_U1671 ( .B1(U_dsdc_n1013), .B2(U_dsdc_n1012), .A(U_dsdc_n338), .ZN(U_dsdc_n1014) );
  OAI21_X2 U_dsdc_U1670 ( .B1(U_dsdc_n1016), .B2(U_dsdc_n338), .A(U_dsdc_n1014), .ZN(U_dsdc_n295) );
  NOR3_X2 U_dsdc_U1669 ( .A1(U_dsdc_n1053), .A2(U_dsdc_n883), .A3(U_dsdc_n822), 
        .ZN(U_dsdc_n932) );
  AOI21_X2 U_dsdc_U1668 ( .B1(U_dsdc_n858), .B2(U_dsdc_n1426), .A(U_dsdc_n857), 
        .ZN(U_dsdc_n907) );
  NOR2_X2 U_dsdc_U1667 ( .A1(U_dsdc_n710), .A2(U_dsdc_n1163), .ZN(U_dsdc_n967)
         );
  NOR2_X2 U_dsdc_U1666 ( .A1(U_dsdc_n907), .A2(U_dsdc_n967), .ZN(U_dsdc_n944)
         );
  NOR2_X2 U_dsdc_U1665 ( .A1(U_dsdc_n691), .A2(U_dsdc_n1293), .ZN(U_dsdc_n1358) );
  NOR2_X2 U_dsdc_U1664 ( .A1(U_dsdc_n866), .A2(U_dsdc_n871), .ZN(U_dsdc_n693)
         );
  NAND2_X2 U_dsdc_U1663 ( .A1(U_dsdc_n1358), .A2(U_dsdc_n693), .ZN(
        U_dsdc_n1802) );
  NAND2_X2 U_dsdc_U1662 ( .A1(U_dsdc_n741), .A2(U_dsdc_n1633), .ZN(
        U_dsdc_n1349) );
  NOR2_X2 U_dsdc_U1661 ( .A1(U_dsdc_n914), .A2(n21), .ZN(U_dsdc_n1041) );
  AOI21_X2 U_dsdc_U1660 ( .B1(U_dsdc_n1348), .B2(U_dsdc_n712), .A(U_dsdc_n711), 
        .ZN(U_dsdc_n945) );
  AOI211_X2 U_dsdc_U1659 ( .C1(U_dsdc_n983), .C2(U_dsdc_n948), .A(U_dsdc_n947), 
        .B(U_dsdc_n946), .ZN(U_dsdc_n955) );
  NAND2_X2 U_dsdc_U1658 ( .A1(U_dsdc_n1437), .A2(U_dsdc_n714), .ZN(U_dsdc_n880) );
  NAND2_X2 U_dsdc_U1657 ( .A1(U_dsdc_n1041), .A2(U_dsdc_n883), .ZN(
        U_dsdc_n1033) );
  NOR2_X2 U_dsdc_U1656 ( .A1(U_dsdc_n1033), .A2(U_dsdc_n2013), .ZN(U_dsdc_n960) );
  NAND2_X2 U_dsdc_U1655 ( .A1(U_dsdc_n887), .A2(U_dsdc_n886), .ZN(U_dsdc_n890)
         );
  NAND2_X2 U_dsdc_U1654 ( .A1(U_dsdc_n1436), .A2(U_cr_n56), .ZN(U_dsdc_n896)
         );
  NAND2_X2 U_dsdc_U1653 ( .A1(U_cr_n39), .A2(n84), .ZN(U_dsdc_n889) );
  NOR2_X2 U_dsdc_U1652 ( .A1(U_dsdc_n896), .A2(U_dsdc_n889), .ZN(U_dsdc_n1032)
         );
  INV_X4 U_dsdc_U1651 ( .A(U_dsdc_n1032), .ZN(U_dsdc_n892) );
  NOR2_X2 U_dsdc_U1650 ( .A1(U_dsdc_n892), .A2(U_dsdc_n1031), .ZN(U_dsdc_n1042) );
  AOI21_X2 U_dsdc_U1649 ( .B1(U_dsdc_n890), .B2(U_dsdc_n1042), .A(U_dsdc_n165), 
        .ZN(U_dsdc_n1310) );
  NAND2_X2 U_dsdc_U1648 ( .A1(U_dsdc_n892), .A2(U_dsdc_n891), .ZN(U_dsdc_n893)
         );
  NAND2_X2 U_dsdc_U1647 ( .A1(U_dsdc_n1310), .A2(U_dsdc_n893), .ZN(
        U_dsdc_n1298) );
  NAND2_X2 U_dsdc_U1646 ( .A1(U_dsdc_n1298), .A2(U_dsdc_n1411), .ZN(
        U_dsdc_n1252) );
  NAND2_X2 U_dsdc_U1645 ( .A1(U_dsdc_n1299), .A2(U_dsdc_n881), .ZN(
        U_dsdc_n1979) );
  NAND3_X2 U_dsdc_U1644 ( .A1(U_dsdc_n894), .A2(U_dsdc_n1252), .A3(
        U_dsdc_n1979), .ZN(U_dsdc_n1374) );
  AOI21_X2 U_dsdc_U1643 ( .B1(U_dsdc_n354), .B2(U_dsdc_n895), .A(U_dsdc_n1374), 
        .ZN(U_dsdc_n954) );
  NOR2_X2 U_dsdc_U1642 ( .A1(U_dsdc_row_cnt_14_), .A2(U_dsdc_row_cnt_12_), 
        .ZN(U_dsdc_n596) );
  NAND3_X2 U_dsdc_U1641 ( .A1(U_dsdc_n596), .A2(U_dsdc_n197), .A3(U_dsdc_n426), 
        .ZN(U_dsdc_n597) );
  NOR2_X2 U_dsdc_U1640 ( .A1(U_dsdc_n1485), .A2(U_dsdc_n1490), .ZN(
        U_dsdc_n1468) );
  INV_X4 U_dsdc_U1639 ( .A(U_dsdc_n1435), .ZN(U_dsdc_n1506) );
  NOR2_X2 U_dsdc_U1638 ( .A1(U_dsdc_n1506), .A2(U_dsdc_n1451), .ZN(
        U_dsdc_n1467) );
  AOI22_X2 U_dsdc_U1637 ( .A1(U_dsdc_n1478), .A2(U_dsdc_n1468), .B1(
        U_dsdc_n1467), .B2(U_cr_n39), .ZN(U_dsdc_n1492) );
  NOR2_X2 U_dsdc_U1636 ( .A1(U_dsdc_n1451), .A2(U_dsdc_n1490), .ZN(
        U_dsdc_n1489) );
  INV_X4 U_dsdc_U1635 ( .A(U_dsdc_n1512), .ZN(U_dsdc_n1521) );
  NOR2_X2 U_dsdc_U1634 ( .A1(U_dsdc_operation_cs_1_), .A2(U_dsdc_n1521), .ZN(
        U_dsdc_n1519) );
  NOR2_X2 U_dsdc_U1633 ( .A1(U_dsdc_operation_cs_3_), .A2(
        U_dsdc_operation_cs_2_), .ZN(U_dsdc_n1450) );
  NAND2_X2 U_dsdc_U1632 ( .A1(U_dsdc_n1450), .A2(U_dsdc_n432), .ZN(
        U_dsdc_n1454) );
  NOR2_X2 U_dsdc_U1631 ( .A1(U_dsdc_n1490), .A2(U_dsdc_n1454), .ZN(
        U_dsdc_n1498) );
  NOR4_X2 U_dsdc_U1630 ( .A1(U_dsdc_n1489), .A2(U_dsdc_n1519), .A3(
        U_dsdc_n1498), .A4(U_dsdc_n1486), .ZN(U_dsdc_n2054) );
  NOR2_X2 U_dsdc_U1629 ( .A1(U_dsdc_n1506), .A2(U_dsdc_n1485), .ZN(
        U_dsdc_n1534) );
  NOR2_X2 U_dsdc_U1628 ( .A1(U_dsdc_n1451), .A2(U_dsdc_n1455), .ZN(
        ctl_sd_in_sf_mode) );
  NOR2_X2 U_dsdc_U1627 ( .A1(U_dsdc_n1534), .A2(ctl_sd_in_sf_mode), .ZN(
        U_dsdc_n2060) );
  NOR2_X2 U_dsdc_U1626 ( .A1(U_dsdc_n1485), .A2(U_dsdc_n1522), .ZN(
        U_dsdc_n2064) );
  NOR2_X2 U_dsdc_U1625 ( .A1(U_dsdc_n1454), .A2(U_dsdc_n1506), .ZN(
        U_dsdc_n1526) );
  INV_X4 U_dsdc_U1624 ( .A(U_dsdc_n1584), .ZN(U_dsdc_n1587) );
  NOR2_X2 U_dsdc_U1623 ( .A1(U_dsdc_rcar_cnt1_3_), .A2(U_dsdc_n1587), .ZN(
        U_dsdc_n1577) );
  NOR2_X2 U_dsdc_U1622 ( .A1(U_dsdc_n1467), .A2(U_dsdc_n1468), .ZN(
        U_dsdc_n1574) );
  NAND2_X2 U_dsdc_U1621 ( .A1(U_dsdc_n1434), .A2(U_dsdc_n642), .ZN(
        U_dsdc_n2051) );
  NOR2_X2 U_dsdc_U1620 ( .A1(U_dsdc_n1577), .A2(U_dsdc_n2051), .ZN(
        U_dsdc_n1565) );
  NOR2_X2 U_dsdc_U1619 ( .A1(U_dsdc_n1454), .A2(U_dsdc_n1522), .ZN(
        U_dsdc_n1432) );
  NAND2_X2 U_dsdc_U1618 ( .A1(U_dsdc_n661), .A2(U_dsdc_n1434), .ZN(
        U_dsdc_n1510) );
  NOR2_X2 U_dsdc_U1617 ( .A1(U_dsdc_n1432), .A2(U_dsdc_n1524), .ZN(
        U_dsdc_n1535) );
  NAND3_X2 U_dsdc_U1616 ( .A1(U_dsdc_n198), .A2(U_dsdc_n427), .A3(U_dsdc_n169), 
        .ZN(U_dsdc_n1509) );
  NOR2_X2 U_dsdc_U1615 ( .A1(U_dsdc_n1535), .A2(U_dsdc_n1431), .ZN(
        U_dsdc_n1617) );
  NOR4_X2 U_dsdc_U1614 ( .A1(U_dsdc_xsr_cnt_0_), .A2(U_dsdc_xsr_cnt_1_), .A3(
        U_dsdc_xsr_cnt_3_), .A4(U_dsdc_xsr_cnt_2_), .ZN(U_dsdc_n1740) );
  INV_X4 U_dsdc_U1613 ( .A(U_dsdc_n1740), .ZN(U_dsdc_n1737) );
  NOR3_X2 U_dsdc_U1612 ( .A1(U_dsdc_xsr_cnt_4_), .A2(U_dsdc_xsr_cnt_5_), .A3(
        U_dsdc_n1737), .ZN(U_dsdc_n1736) );
  NAND2_X2 U_dsdc_U1611 ( .A1(U_dsdc_n1736), .A2(U_dsdc_n359), .ZN(
        U_dsdc_n1727) );
  NOR2_X2 U_dsdc_U1610 ( .A1(U_dsdc_n1451), .A2(U_dsdc_n1522), .ZN(
        U_dsdc_n1536) );
  NOR2_X2 U_dsdc_U1609 ( .A1(U_dsdc_n1728), .A2(U_dsdc_n1452), .ZN(
        U_dsdc_n1500) );
  NOR4_X2 U_dsdc_U1608 ( .A1(U_dsdc_n1800), .A2(U_dsdc_n1565), .A3(
        U_dsdc_n1617), .A4(U_dsdc_n1500), .ZN(U_dsdc_n1453) );
  NAND3_X2 U_dsdc_U1607 ( .A1(U_dsdc_n1492), .A2(U_dsdc_n930), .A3(
        U_dsdc_n1453), .ZN(U_dsdc_n952) );
  NAND2_X2 U_dsdc_U1606 ( .A1(U_dsdc_n199), .A2(U_dsdc_n429), .ZN(U_dsdc_n1491) );
  INV_X4 U_dsdc_U1605 ( .A(U_dsdc_n1491), .ZN(U_dsdc_n1430) );
  NOR3_X2 U_dsdc_U1604 ( .A1(U_dsdc_n1490), .A2(U_dsdc_n1430), .A3(U_dsdc_n949), .ZN(U_dsdc_n951) );
  NAND2_X2 U_dsdc_U1603 ( .A1(U_dsdc_n662), .A2(U_dsdc_n661), .ZN(U_dsdc_n2058) );
  NOR4_X2 U_dsdc_U1602 ( .A1(U_dsdc_n952), .A2(U_dsdc_n951), .A3(U_dsdc_n1511), 
        .A4(U_dsdc_n950), .ZN(U_dsdc_n953) );
  AOI21_X2 U_dsdc_U1601 ( .B1(U_dsdc_n955), .B2(U_dsdc_n954), .A(U_dsdc_n953), 
        .ZN(U_dsdc_N403) );
  NAND3_X2 U_dsdc_U1599 ( .A1(U_dsdc_n913), .A2(U_dsdc_n848), .A3(U_dsdc_n847), 
        .ZN(U_dsdc_n899) );
  NOR2_X2 U_dsdc_U1598 ( .A1(U_dsdc_n851), .A2(U_dsdc_n1546), .ZN(U_dsdc_n878)
         );
  OAI211_X2 U_dsdc_U1597 ( .C1(U_dsdc_n1353), .C2(U_dsdc_n939), .A(
        U_dsdc_n1352), .B(U_dsdc_n854), .ZN(U_dsdc_n908) );
  NOR2_X2 U_dsdc_U1596 ( .A1(U_dsdc_n165), .A2(U_dsdc_n1980), .ZN(U_dsdc_n1456) );
  NAND2_X2 U_dsdc_U1595 ( .A1(U_dsdc_n1300), .A2(U_dsdc_n1456), .ZN(
        U_dsdc_n902) );
  AOI211_X2 U_dsdc_U1594 ( .C1(U_dsdc_n916), .C2(U_dsdc_n864), .A(U_dsdc_n863), 
        .B(U_dsdc_n862), .ZN(U_dsdc_n875) );
  AOI211_X2 U_dsdc_U1593 ( .C1(U_dsdc_n1416), .C2(U_dsdc_n1152), .A(
        U_dsdc_n870), .B(U_dsdc_n1350), .ZN(U_dsdc_n922) );
  NAND4_X2 U_dsdc_U1592 ( .A1(U_dsdc_n2069), .A2(U_dsdc_n2071), .A3(
        U_dsdc_n1309), .A4(U_dsdc_n872), .ZN(U_dsdc_n873) );
  NAND2_X2 U_dsdc_U1591 ( .A1(U_dsdc_n725), .A2(U_dsdc_n710), .ZN(U_dsdc_n1974) );
  NOR4_X2 U_dsdc_U1590 ( .A1(U_dsdc_n878), .A2(U_dsdc_n908), .A3(U_dsdc_n877), 
        .A4(U_dsdc_n876), .ZN(U_dsdc_n898) );
  NOR2_X2 U_dsdc_U1589 ( .A1(U_dsdc_n952), .A2(U_dsdc_n897), .ZN(U_dsdc_n909)
         );
  AOI21_X2 U_dsdc_U1588 ( .B1(U_dsdc_n898), .B2(U_dsdc_n954), .A(U_dsdc_n909), 
        .ZN(U_dsdc_N401) );
  NAND2_X2 U_dsdc_U1587 ( .A1(U_dsdc_n1557), .A2(U_dsdc_n1438), .ZN(
        U_dsdc_n1372) );
  INV_X4 U_dsdc_U1586 ( .A(U_dsdc_n1372), .ZN(U_dsdc_n1043) );
  AOI21_X2 U_dsdc_U1585 ( .B1(U_dsdc_n1061), .B2(U_dsdc_n703), .A(U_dsdc_n2071), .ZN(U_dsdc_n1367) );
  AOI21_X2 U_dsdc_U1584 ( .B1(U_dsdc_access_cs_2_), .B2(U_dsdc_n915), .A(
        U_dsdc_n1367), .ZN(U_dsdc_n919) );
  AOI21_X2 U_dsdc_U1583 ( .B1(U_dsdc_n903), .B2(U_dsdc_n181), .A(U_dsdc_n934), 
        .ZN(U_dsdc_n917) );
  OAI21_X2 U_dsdc_U1582 ( .B1(U_dsdc_n917), .B2(U_dsdc_n1415), .A(U_dsdc_n916), 
        .ZN(U_dsdc_n918) );
  OAI21_X2 U_dsdc_U1581 ( .B1(U_dsdc_r_rw), .B2(U_dsdc_n967), .A(U_dsdc_n1974), 
        .ZN(U_dsdc_n958) );
  AOI211_X2 U_dsdc_U1580 ( .C1(U_dsdc_n925), .C2(U_dsdc_n983), .A(U_dsdc_n924), 
        .B(U_dsdc_n923), .ZN(U_dsdc_n931) );
  NOR4_X2 U_dsdc_U1579 ( .A1(U_dsdc_num_init_ref_cnt_0_), .A2(
        U_dsdc_num_init_ref_cnt_1_), .A3(U_dsdc_num_init_ref_cnt_2_), .A4(
        U_dsdc_num_init_ref_cnt_3_), .ZN(U_dsdc_n1564) );
  INV_X4 U_dsdc_U1578 ( .A(U_dsdc_n2051), .ZN(U_dsdc_n1433) );
  NOR2_X2 U_dsdc_U1577 ( .A1(cr_do_initialize), .A2(U_dsdc_n1470), .ZN(
        U_dsdc_n1466) );
  NAND2_X2 U_dsdc_U1576 ( .A1(U_dsdc_n1436), .A2(U_dsdc_n1466), .ZN(
        U_dsdc_n2052) );
  NOR2_X2 U_dsdc_U1575 ( .A1(U_dsdc_n2052), .A2(U_cr_n39), .ZN(U_dsdc_n1758)
         );
  NAND2_X2 U_dsdc_U1574 ( .A1(U_dsdc_n1432), .A2(U_dsdc_n1509), .ZN(
        U_dsdc_n1501) );
  NOR2_X2 U_dsdc_U1573 ( .A1(U_dsdc_n1485), .A2(U_dsdc_n1455), .ZN(
        U_dsdc_n1581) );
  NOR4_X2 U_dsdc_U1572 ( .A1(U_dsdc_n362), .A2(U_dsdc_n1758), .A3(U_dsdc_n928), 
        .A4(U_dsdc_n927), .ZN(U_dsdc_n929) );
  AOI22_X2 U_dsdc_U1571 ( .A1(U_dsdc_n954), .A2(U_dsdc_n931), .B1(U_dsdc_n930), 
        .B2(U_dsdc_n929), .ZN(U_dsdc_N404) );
  NAND2_X2 U_dsdc_U1570 ( .A1(U_dsdc_n2071), .A2(U_dsdc_n934), .ZN(U_dsdc_n956) );
  NOR4_X2 U_dsdc_U1569 ( .A1(U_dsdc_n1802), .A2(U_dsdc_n956), .A3(U_dsdc_n1349), .A4(U_dsdc_n1425), .ZN(U_dsdc_n959) );
  NAND4_X2 U_dsdc_U1568 ( .A1(U_dsdc_n972), .A2(U_dsdc_n959), .A3(U_dsdc_n958), 
        .A4(U_dsdc_n957), .ZN(U_dsdc_n963) );
  NOR3_X2 U_dsdc_U1567 ( .A1(U_dsdc_r_bm_close_bank_3_), .A2(U_dsdc_n396), 
        .A3(U_dsdc_n1942), .ZN(U_dsdc_n1907) );
  NOR3_X2 U_dsdc_U1566 ( .A1(U_dsdc_r_bm_open_bank[3]), .A2(U_dsdc_n1941), 
        .A3(U_dsdc_n396), .ZN(U_dsdc_n1906) );
  INV_X4 U_dsdc_U1565 ( .A(U_dsdc_n1906), .ZN(U_dsdc_n1900) );
  INV_X4 U_dsdc_U1564 ( .A(U_dsdc_n1907), .ZN(U_dsdc_n1899) );
  AOI22_X2 U_dsdc_U1563 ( .A1(U_dsdc_n302), .A2(U_dsdc_n1943), .B1(U_dsdc_n303), .B2(U_dsdc_n1951), .ZN(U_dsdc_n1882) );
  OAI221_X2 U_dsdc_U1562 ( .B1(U_dsdc_bm_bank_age_3__0_), .B2(
        U_dsdc_bm_bank_age_3__1_), .C1(U_dsdc_bm_bank_age_3__0_), .C2(
        U_dsdc_n1944), .A(U_dsdc_n1882), .ZN(U_dsdc_n1884) );
  AOI221_X2 U_dsdc_U1561 ( .B1(U_dsdc_n1945), .B2(U_dsdc_n1885), .C1(
        U_dsdc_n1884), .C2(U_dsdc_n1885), .A(U_dsdc_n1883), .ZN(U_dsdc_n1886)
         );
  AOI21_X2 U_dsdc_U1560 ( .B1(U_dsdc_bm_bank_age_3__3_), .B2(U_dsdc_n1953), 
        .A(U_dsdc_n1886), .ZN(U_dsdc_n1887) );
  AOI222_X2 U_dsdc_U1559 ( .A1(U_dsdc_n1887), .A2(U_dsdc_n351), .B1(
        U_dsdc_n1887), .B2(U_dsdc_n1954), .C1(U_dsdc_n351), .C2(U_dsdc_n1954), 
        .ZN(U_dsdc_n1890) );
  NAND3_X2 U_dsdc_U1558 ( .A1(U_dsdc_n302), .A2(U_dsdc_n304), .A3(U_dsdc_n1890), .ZN(U_dsdc_n1896) );
  AOI21_X2 U_dsdc_U1557 ( .B1(U_dsdc_bm_bank_age_3__1_), .B2(
        U_dsdc_bm_bank_age_3__0_), .A(U_dsdc_n1900), .ZN(U_dsdc_n1895) );
  AOI211_X2 U_dsdc_U1556 ( .C1(U_dsdc_n1907), .C2(U_dsdc_n1896), .A(
        U_dsdc_n1961), .B(U_dsdc_n1895), .ZN(U_dsdc_n1898) );
  OAI221_X2 U_dsdc_U1555 ( .B1(U_dsdc_bm_bank_age_3__2_), .B2(U_dsdc_n1900), 
        .C1(U_dsdc_n303), .C2(U_dsdc_n1899), .A(U_dsdc_n1898), .ZN(
        U_dsdc_n1905) );
  AOI221_X2 U_dsdc_U1554 ( .B1(U_dsdc_n1907), .B2(U_dsdc_bm_bank_age_3__3_), 
        .C1(U_dsdc_n1906), .C2(U_dsdc_n284), .A(U_dsdc_n1905), .ZN(
        U_dsdc_n1910) );
  NOR2_X2 U_dsdc_U1553 ( .A1(U_dsdc_n303), .A2(U_dsdc_n1901), .ZN(U_dsdc_n1908) );
  AOI22_X2 U_dsdc_U1552 ( .A1(U_dsdc_bm_bank_age_3__4_), .A2(U_dsdc_n1910), 
        .B1(U_dsdc_n1909), .B2(U_dsdc_n351), .ZN(U_dsdc_n222) );
  NOR2_X2 U_dsdc_U1551 ( .A1(U_dsdc_n1203), .A2(U_dsdc_bm_rc_cnt_2__2_), .ZN(
        U_dsdc_n1207) );
  NOR2_X2 U_dsdc_U1550 ( .A1(U_dsdc_n1207), .A2(U_dsdc_n439), .ZN(U_dsdc_n1208) );
  NOR2_X2 U_dsdc_U1549 ( .A1(U_dsdc_n1189), .A2(U_dsdc_bm_rc_cnt_1__2_), .ZN(
        U_dsdc_n1193) );
  NOR2_X2 U_dsdc_U1548 ( .A1(U_dsdc_n1193), .A2(U_dsdc_n438), .ZN(U_dsdc_n1194) );
  NAND2_X2 U_dsdc_U1547 ( .A1(U_dsdc_n1166), .A2(U_dsdc_n604), .ZN(U_dsdc_n307) );
  INV_X4 U_dsdc_U1546 ( .A(U_dsdc_n307), .ZN(U_dsdc_n621) );
  AOI211_X2 U_dsdc_U1545 ( .C1(U_dsdc_n964), .C2(U_dsdc_pre_amble_mute), .A(
        U_dsdc_n1411), .B(U_dsdc_n963), .ZN(U_dsdc_n965) );
  INV_X4 U_dsdc_U1544 ( .A(U_dsdc_n965), .ZN(U_dsdc_pre_amble_nxt) );
  INV_X4 U_dsdc_U1543 ( .A(U_dsdc_n1011), .ZN(U_dsdc_n1009) );
  OAI211_X2 U_dsdc_U1542 ( .C1(U_dsdc_n1009), .C2(U_dsdc_n180), .A(
        U_dsdc_n1017), .B(U_dsdc_n1008), .ZN(U_dsdc_n294) );
  NAND2_X2 U_dsdc_U1541 ( .A1(U_dsdc_n960), .A2(U_dsdc_n1032), .ZN(
        U_dsdc_n1289) );
  NAND2_X2 U_dsdc_U1540 ( .A1(U_dsdc_n1289), .A2(U_dsdc_n1252), .ZN(
        U_dsdc_n1039) );
  AOI22_X2 U_dsdc_U1539 ( .A1(hiu_terminate), .A2(U_dsdc_n166), .B1(
        U_dsdc_n1040), .B2(U_dsdc_n1039), .ZN(U_dsdc_n1050) );
  NAND2_X2 U_dsdc_U1538 ( .A1(U_dsdc_n1320), .A2(U_dsdc_n1044), .ZN(
        U_dsdc_n1051) );
  NAND2_X2 U_dsdc_U1537 ( .A1(U_dsdc_n619), .A2(U_dsdc_n166), .ZN(U_dsdc_n1314) );
  INV_X4 U_dsdc_U1536 ( .A(U_dsdc_n1314), .ZN(U_dsdc_n1048) );
  AOI22_X2 U_dsdc_U1535 ( .A1(U_dsdc_n1051), .A2(ad_data_mask[1]), .B1(
        U_dsdc_r_data_mask[1]), .B2(U_dsdc_n1048), .ZN(U_dsdc_n1046) );
  NAND2_X2 U_dsdc_U1534 ( .A1(U_dsdc_n1050), .A2(U_dsdc_n1046), .ZN(
        U_dsdc_N426) );
  AOI22_X2 U_dsdc_U1533 ( .A1(U_dsdc_n1051), .A2(ad_data_mask[0]), .B1(
        U_dsdc_r_data_mask[0]), .B2(U_dsdc_n1048), .ZN(U_dsdc_n1045) );
  NAND2_X2 U_dsdc_U1532 ( .A1(U_dsdc_n1050), .A2(U_dsdc_n1045), .ZN(
        U_dsdc_N425) );
  AOI22_X2 U_dsdc_U1531 ( .A1(U_dsdc_n1051), .A2(ad_data_mask[3]), .B1(
        U_dsdc_r_data_mask[3]), .B2(U_dsdc_n1048), .ZN(U_dsdc_n1049) );
  NAND2_X2 U_dsdc_U1530 ( .A1(U_dsdc_n1050), .A2(U_dsdc_n1049), .ZN(
        U_dsdc_N428) );
  AOI22_X2 U_dsdc_U1529 ( .A1(U_dsdc_n1051), .A2(ad_data_mask[2]), .B1(
        U_dsdc_r_data_mask[2]), .B2(U_dsdc_n1048), .ZN(U_dsdc_n1047) );
  NAND2_X2 U_dsdc_U1528 ( .A1(U_dsdc_n1050), .A2(U_dsdc_n1047), .ZN(
        U_dsdc_N427) );
  AOI21_X2 U_dsdc_U1527 ( .B1(U_dsdc_n1413), .B2(U_dsdc_n672), .A(U_dsdc_n669), 
        .ZN(U_dsdc_n1409) );
  NOR2_X2 U_dsdc_U1526 ( .A1(U_dsdc_n1124), .A2(U_dsdc_n1056), .ZN(
        U_dsdc_n1057) );
  INV_X4 U_dsdc_U1525 ( .A(U_dsdc_n1268), .ZN(U_dsdc_n1260) );
  OAI22_X2 U_dsdc_U1524 ( .A1(U_dsdc_n1064), .A2(U_dsdc_n1457), .B1(
        U_dsdc_n2071), .B2(U_dsdc_n1312), .ZN(U_dsdc_n1067) );
  NOR2_X2 U_dsdc_U1523 ( .A1(U_dsdc_n1067), .A2(U_dsdc_n1066), .ZN(
        U_dsdc_n1068) );
  NAND2_X2 U_dsdc_U1522 ( .A1(U_dsdc_i_col_addr_1_), .A2(U_dsdc_i_col_addr_2_), 
        .ZN(U_dsdc_n1810) );
  NOR2_X2 U_dsdc_U1521 ( .A1(U_dsdc_n1810), .A2(U_dsdc_n443), .ZN(U_dsdc_n699)
         );
  NAND2_X2 U_dsdc_U1520 ( .A1(U_dsdc_i_col_addr_6_), .A2(U_dsdc_i_col_addr_7_), 
        .ZN(U_dsdc_n671) );
  NOR2_X2 U_dsdc_U1519 ( .A1(U_dsdc_n681), .A2(U_dsdc_n671), .ZN(U_dsdc_n697)
         );
  NAND3_X2 U_dsdc_U1518 ( .A1(U_dsdc_n697), .A2(U_dsdc_i_col_addr_9_), .A3(
        U_dsdc_i_col_addr_8_), .ZN(U_dsdc_n702) );
  NOR2_X2 U_dsdc_U1517 ( .A1(U_dsdc_n702), .A2(U_dsdc_n444), .ZN(U_dsdc_n701)
         );
  NAND2_X2 U_dsdc_U1516 ( .A1(U_dsdc_n701), .A2(U_dsdc_i_col_addr_11_), .ZN(
        U_dsdc_n700) );
  NAND2_X2 U_dsdc_U1515 ( .A1(U_dsdc_n677), .A2(U_dsdc_i_col_addr_12_), .ZN(
        U_dsdc_n678) );
  OAI211_X2 U_dsdc_U1514 ( .C1(U_dsdc_n1142), .C2(debug_ad_col_addr_13_), .A(
        U_dsdc_n1168), .B(U_dsdc_n1135), .ZN(U_dsdc_s_addr_nxt_a[14]) );
  NOR2_X2 U_dsdc_U1513 ( .A1(U_dsdc_t_xp_cnt_1_), .A2(U_dsdc_t_xp_cnt_0_), 
        .ZN(U_dsdc_n1482) );
  INV_X4 U_dsdc_U1512 ( .A(U_dsdc_n1534), .ZN(U_dsdc_n2057) );
  AOI21_X2 U_dsdc_U1511 ( .B1(U_dsdc_n1466), .B2(U_dsdc_n1465), .A(
        U_dsdc_n1581), .ZN(U_dsdc_n1540) );
  INV_X4 U_dsdc_U1510 ( .A(U_dsdc_n1467), .ZN(U_dsdc_n2066) );
  INV_X4 U_dsdc_U1509 ( .A(U_dsdc_n1468), .ZN(U_dsdc_n2059) );
  OAI22_X2 U_dsdc_U1508 ( .A1(U_dsdc_n1482), .A2(U_dsdc_n1471), .B1(
        U_dsdc_n1470), .B2(U_dsdc_n1469), .ZN(U_dsdc_n1472) );
  NOR4_X2 U_dsdc_U1507 ( .A1(U_dsdc_n1800), .A2(U_dsdc_n1576), .A3(U_dsdc_n362), .A4(U_dsdc_n1472), .ZN(U_dsdc_n1503) );
  NOR4_X2 U_dsdc_U1506 ( .A1(U_dsdc_init_cnt_0_), .A2(U_dsdc_init_cnt_1_), 
        .A3(U_dsdc_init_cnt_2_), .A4(U_dsdc_init_cnt_3_), .ZN(U_dsdc_n1708) );
  NOR3_X2 U_dsdc_U1505 ( .A1(U_dsdc_init_cnt_5_), .A2(U_dsdc_init_cnt_4_), 
        .A3(U_dsdc_n1704), .ZN(U_dsdc_n1701) );
  NOR3_X2 U_dsdc_U1504 ( .A1(U_dsdc_init_cnt_7_), .A2(U_dsdc_init_cnt_6_), 
        .A3(U_dsdc_n1697), .ZN(U_dsdc_n1694) );
  NOR3_X2 U_dsdc_U1503 ( .A1(U_dsdc_init_cnt_9_), .A2(U_dsdc_init_cnt_8_), 
        .A3(U_dsdc_n1690), .ZN(U_dsdc_n1687) );
  NOR3_X2 U_dsdc_U1502 ( .A1(U_dsdc_init_cnt_11_), .A2(U_dsdc_init_cnt_10_), 
        .A3(U_dsdc_n1683), .ZN(U_dsdc_n1679) );
  NOR2_X2 U_dsdc_U1501 ( .A1(U_dsdc_init_cnt_13_), .A2(U_dsdc_init_cnt_12_), 
        .ZN(U_dsdc_n481) );
  NAND2_X2 U_dsdc_U1500 ( .A1(U_dsdc_n1679), .A2(U_dsdc_n481), .ZN(U_dsdc_n482) );
  AOI211_X2 U_dsdc_U1499 ( .C1(U_dsdc_n1474), .C2(U_dsdc_n1473), .A(
        U_dsdc_n1521), .B(U_dsdc_n1522), .ZN(U_dsdc_n1475) );
  AOI211_X2 U_dsdc_U1498 ( .C1(U_dsdc_n1526), .C2(U_dsdc_n1675), .A(
        U_dsdc_n2064), .B(U_dsdc_n1475), .ZN(U_dsdc_n1504) );
  AOI21_X2 U_dsdc_U1497 ( .B1(U_dsdc_n1489), .B2(U_dsdc_n1476), .A(
        U_dsdc_n1536), .ZN(U_dsdc_n1477) );
  NAND3_X2 U_dsdc_U1496 ( .A1(U_dsdc_n1503), .A2(U_dsdc_n1504), .A3(
        U_dsdc_n1477), .ZN(U_dsdc_n1533) );
  INV_X4 U_dsdc_U1495 ( .A(ctl_sd_in_sf_mode), .ZN(U_dsdc_n1532) );
  OAI21_X2 U_dsdc_U1494 ( .B1(U_dsdc_n2057), .B2(U_dsdc_n2056), .A(
        U_dsdc_n1532), .ZN(U_dsdc_n1523) );
  NAND2_X2 U_dsdc_U1493 ( .A1(U_dsdc_n1479), .A2(U_dsdc_n1482), .ZN(
        U_dsdc_n1537) );
  OAI22_X2 U_dsdc_U1492 ( .A1(U_dsdc_n2066), .A2(U_dsdc_n2062), .B1(n84), .B2(
        U_dsdc_n1537), .ZN(U_dsdc_n1525) );
  AOI221_X2 U_dsdc_U1491 ( .B1(U_dsdc_n1533), .B2(U_dsdc_operation_cs_3_), 
        .C1(U_dsdc_n1523), .C2(U_dsdc_operation_cs_3_), .A(U_dsdc_n1525), .ZN(
        U_dsdc_n1481) );
  NAND2_X2 U_dsdc_U1490 ( .A1(U_dsdc_n644), .A2(U_dsdc_n1433), .ZN(
        U_dsdc_n1480) );
  NAND4_X2 U_dsdc_U1489 ( .A1(U_dsdc_n1540), .A2(U_dsdc_n1481), .A3(
        U_dsdc_n1579), .A4(U_dsdc_n1480), .ZN(U_dsdc_n2094) );
  OAI22_X2 U_dsdc_U1488 ( .A1(U_dsdc_t_xp_cnt_0_), .A2(U_dsdc_n1482), .B1(
        U_dsdc_n2057), .B2(U_dsdc_n2094), .ZN(U_dsdc_N4228) );
  NAND3_X2 U_dsdc_U1487 ( .A1(U_dsdc_n1503), .A2(U_dsdc_n1502), .A3(
        U_dsdc_n1501), .ZN(U_dsdc_n1518) );
  AOI211_X2 U_dsdc_U1486 ( .C1(U_dsdc_n2064), .C2(U_dsdc_n2063), .A(
        U_dsdc_n1519), .B(U_dsdc_n1518), .ZN(U_dsdc_n1520) );
  OAI21_X2 U_dsdc_U1485 ( .B1(U_dsdc_n1522), .B2(U_dsdc_n1521), .A(
        U_dsdc_n1520), .ZN(U_dsdc_n1542) );
  NOR3_X2 U_dsdc_U1484 ( .A1(U_dsdc_n1524), .A2(U_dsdc_n1523), .A3(
        U_dsdc_n1542), .ZN(U_dsdc_n1530) );
  NOR2_X2 U_dsdc_U1483 ( .A1(U_dsdc_n2065), .A2(U_dsdc_n1675), .ZN(
        U_dsdc_n2061) );
  OAI21_X2 U_dsdc_U1482 ( .B1(U_dsdc_n1491), .B2(U_dsdc_n1505), .A(
        U_dsdc_n2058), .ZN(U_dsdc_n1618) );
  AOI211_X2 U_dsdc_U1481 ( .C1(U_dsdc_n1430), .C2(U_dsdc_n1519), .A(
        ctl_init_done), .B(U_dsdc_n1493), .ZN(U_dsdc_n1507) );
  NOR4_X2 U_dsdc_U1480 ( .A1(U_dsdc_n1581), .A2(U_dsdc_n2061), .A3(
        U_dsdc_n1618), .A4(U_dsdc_n1527), .ZN(U_dsdc_n1528) );
  OAI211_X2 U_dsdc_U1479 ( .C1(U_dsdc_n1530), .C2(U_dsdc_n343), .A(
        U_dsdc_n1529), .B(U_dsdc_n1528), .ZN(U_dsdc_n2096) );
  OAI21_X2 U_dsdc_U1478 ( .B1(U_dsdc_n2064), .B2(U_dsdc_n1575), .A(
        U_dsdc_n2063), .ZN(U_dsdc_n1588) );
  NOR2_X2 U_dsdc_U1477 ( .A1(U_dsdc_n1510), .A2(U_dsdc_n1509), .ZN(
        U_dsdc_n1667) );
  NOR3_X2 U_dsdc_U1476 ( .A1(U_dsdc_n1564), .A2(U_dsdc_n2051), .A3(
        U_dsdc_n2063), .ZN(U_dsdc_n1580) );
  INV_X4 U_dsdc_U1475 ( .A(U_dsdc_n1576), .ZN(U_dsdc_n573) );
  NAND2_X2 U_dsdc_U1474 ( .A1(U_dsdc_n1536), .A2(U_dsdc_n1728), .ZN(
        U_dsdc_n1578) );
  OAI22_X2 U_dsdc_U1472 ( .A1(U_dsdc_rcar_cnt1_0_), .A2(U_dsdc_n1588), .B1(
        U_dsdc_n1590), .B2(U_cr_n127), .ZN(U_dsdc_rcar_cnt1_nxt[0]) );
  OAI22_X2 U_dsdc_U1471 ( .A1(U_dsdc_n2057), .A2(U_dsdc_n2094), .B1(
        U_dsdc_n474), .B2(U_dsdc_n239), .ZN(U_dsdc_N4229) );
  NAND3_X2 U_dsdc_U1470 ( .A1(U_dsdc_n645), .A2(U_dsdc_n1430), .A3(
        U_dsdc_n1434), .ZN(U_dsdc_n1497) );
  AOI21_X2 U_dsdc_U1469 ( .B1(U_dsdc_n1499), .B2(cr_do_initialize), .A(
        U_dsdc_n1498), .ZN(U_dsdc_n1676) );
  AOI21_X2 U_dsdc_U1468 ( .B1(U_dsdc_n1534), .B2(U_dsdc_n2056), .A(
        U_dsdc_n1527), .ZN(U_dsdc_n1544) );
  AOI211_X2 U_dsdc_U1467 ( .C1(U_dsdc_n1512), .C2(U_dsdc_n1435), .A(
        U_dsdc_n1511), .B(U_dsdc_n1667), .ZN(U_dsdc_n1514) );
  NOR2_X2 U_dsdc_U1466 ( .A1(U_dsdc_n2052), .A2(cr_do_self_ref_rp), .ZN(
        U_dsdc_n1429) );
  NAND3_X2 U_dsdc_U1465 ( .A1(U_dsdc_n1429), .A2(cr_exn_mode_reg_update), .A3(
        U_cr_n61), .ZN(U_dsdc_n1513) );
  NAND4_X2 U_dsdc_U1464 ( .A1(U_dsdc_n1544), .A2(U_dsdc_n1514), .A3(
        U_dsdc_n1579), .A4(U_dsdc_n1513), .ZN(U_dsdc_n1515) );
  AOI221_X2 U_dsdc_U1463 ( .B1(U_dsdc_n1518), .B2(U_dsdc_operation_cs_0_), 
        .C1(U_dsdc_n1516), .C2(U_dsdc_operation_cs_0_), .A(U_dsdc_n1515), .ZN(
        U_dsdc_n1517) );
  NAND4_X2 U_dsdc_U1462 ( .A1(U_dsdc_n1540), .A2(U_dsdc_n1733), .A3(
        U_dsdc_n1676), .A4(U_dsdc_n1517), .ZN(U_dsdc_n2097) );
  AOI21_X2 U_dsdc_U1461 ( .B1(U_dsdc_rcar_cnt1_0_), .B2(U_dsdc_rcar_cnt1_1_), 
        .A(U_dsdc_n1583), .ZN(U_dsdc_n1582) );
  NOR2_X2 U_dsdc_U1459 ( .A1(U_dsdc_n1326), .A2(U_dsdc_n1325), .ZN(
        U_dsdc_n1328) );
  AOI21_X2 U_dsdc_U1458 ( .B1(U_dsdc_n1327), .B2(cr_t_rp[0]), .A(U_dsdc_n1336), 
        .ZN(U_dsdc_n1333) );
  NOR2_X2 U_dsdc_U1457 ( .A1(U_dsdc_n1328), .A2(cr_t_rp[0]), .ZN(U_dsdc_n1334)
         );
  NOR2_X2 U_dsdc_U1456 ( .A1(U_cr_n148), .A2(cr_t_rp[1]), .ZN(U_dsdc_n1331) );
  NOR2_X2 U_dsdc_U1455 ( .A1(U_dsdc_n1357), .A2(U_dsdc_n1425), .ZN(
        U_dsdc_n1421) );
  AOI21_X2 U_dsdc_U1454 ( .B1(U_dsdc_n1421), .B2(U_dsdc_n1629), .A(
        U_dsdc_n1426), .ZN(U_dsdc_n1335) );
  AOI22_X2 U_dsdc_U1453 ( .A1(U_dsdc_n1334), .A2(U_dsdc_n1331), .B1(
        U_dsdc_n1335), .B2(U_dsdc_n1330), .ZN(U_dsdc_n1332) );
  OAI21_X2 U_dsdc_U1452 ( .B1(U_dsdc_n1333), .B2(U_cr_n147), .A(U_dsdc_n1332), 
        .ZN(U_dsdc_rp_cnt2_nxt[1]) );
  INV_X4 U_dsdc_U1451 ( .A(U_dsdc_n1349), .ZN(U_dsdc_n1397) );
  NAND2_X2 U_dsdc_U1450 ( .A1(U_dsdc_n1637), .A2(U_dsdc_n1414), .ZN(
        U_dsdc_n1805) );
  NAND2_X2 U_dsdc_U1449 ( .A1(U_dsdc_n915), .A2(U_dsdc_n652), .ZN(U_dsdc_n1803) );
  NAND2_X2 U_dsdc_U1448 ( .A1(U_dsdc_n1804), .A2(U_dsdc_n1803), .ZN(
        U_dsdc_n2074) );
  NOR2_X2 U_dsdc_U1447 ( .A1(U_dsdc_n2074), .A2(U_dsdc_n360), .ZN(U_dsdc_n1398) );
  AOI21_X2 U_dsdc_U1446 ( .B1(U_dsdc_n740), .B2(U_dsdc_n736), .A(U_dsdc_n728), 
        .ZN(U_dsdc_n730) );
  OAI21_X2 U_dsdc_U1445 ( .B1(U_dsdc_n730), .B2(U_dsdc_n440), .A(U_dsdc_n729), 
        .ZN(U_dsdc_n731) );
  AOI21_X2 U_dsdc_U1444 ( .B1(U_dsdc_n1805), .B2(U_dsdc_n1415), .A(U_dsdc_n731), .ZN(U_dsdc_n732) );
  OAI211_X2 U_dsdc_U1443 ( .C1(U_dsdc_n1397), .C2(U_dsdc_n733), .A(
        U_dsdc_n1398), .B(U_dsdc_n732), .ZN(U_dsdc_n734) );
  NOR2_X2 U_dsdc_U1442 ( .A1(hiu_terminate), .A2(U_dsdc_n734), .ZN(U_dsdc_n329) );
  OAI211_X2 U_dsdc_U1441 ( .C1(U_dsdc_n1142), .C2(debug_ad_col_addr_12_), .A(
        U_dsdc_n1169), .B(U_dsdc_n1133), .ZN(U_dsdc_s_addr_nxt_a[13]) );
  NAND2_X2 U_dsdc_U1440 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_1_), .ZN(
        U_dsdc_n1812) );
  NAND3_X2 U_dsdc_U1439 ( .A1(U_dsdc_n1480), .A2(U_dsdc_n646), .A3(
        U_dsdc_n1497), .ZN(U_dsdc_n1670) );
  AOI211_X2 U_dsdc_U1438 ( .C1(cr_exn_mode_value[1]), .C2(U_dsdc_n1671), .A(
        U_dsdc_n1118), .B(U_dsdc_n1670), .ZN(U_dsdc_n1119) );
  OAI211_X2 U_dsdc_U1437 ( .C1(U_dsdc_n1142), .C2(U_addrdec_n96), .A(
        U_dsdc_n1172), .B(U_dsdc_n1119), .ZN(U_dsdc_N419) );
  NOR2_X2 U_dsdc_U1436 ( .A1(U_dsdc_n678), .A2(U_dsdc_n446), .ZN(U_dsdc_n679)
         );
  AOI22_X2 U_dsdc_U1435 ( .A1(U_dsdc_n1139), .A2(U_dsdc_n1138), .B1(
        U_dsdc_r_col_addr_14_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1140) );
  OAI211_X2 U_dsdc_U1434 ( .C1(U_dsdc_n1142), .C2(U_dsdc_n1141), .A(
        U_dsdc_n1167), .B(U_dsdc_n1140), .ZN(U_dsdc_s_addr_nxt_a[15]) );
  AOI21_X2 U_dsdc_U1433 ( .B1(U_dsdc_n1295), .B2(U_dsdc_n1294), .A(
        U_dsdc_n1293), .ZN(U_dsdc_n1307) );
  AOI21_X2 U_dsdc_U1432 ( .B1(U_dsdc_wr_cnt_2_), .B2(U_dsdc_n1297), .A(
        U_dsdc_n1296), .ZN(U_dsdc_n1303) );
  AOI21_X2 U_dsdc_U1431 ( .B1(U_dsdc_n1300), .B2(U_dsdc_n1299), .A(
        U_dsdc_n1298), .ZN(U_dsdc_n1301) );
  NOR2_X2 U_dsdc_U1430 ( .A1(U_dsdc_n1301), .A2(U_dsdc_n1309), .ZN(
        U_dsdc_n1304) );
  NAND3_X2 U_dsdc_U1429 ( .A1(U_dsdc_n1304), .A2(cr_t_wr[0]), .A3(cr_t_wr[1]), 
        .ZN(U_dsdc_n1302) );
  OAI21_X2 U_dsdc_U1428 ( .B1(U_dsdc_n1307), .B2(U_dsdc_n1303), .A(
        U_dsdc_n1302), .ZN(U_dsdc_wr_cnt_nxt[2]) );
  NAND2_X2 U_dsdc_U1427 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_4_), .ZN(
        U_dsdc_n1550) );
  OAI211_X2 U_dsdc_U1426 ( .C1(U_dsdc_n1108), .C2(n90), .A(U_dsdc_n1107), .B(
        U_dsdc_n1550), .ZN(U_dsdc_n1113) );
  AOI211_X2 U_dsdc_U1425 ( .C1(U_dsdc_n1138), .C2(U_dsdc_n1406), .A(
        U_dsdc_n1113), .B(U_dsdc_n1221), .ZN(U_dsdc_n1114) );
  OAI21_X2 U_dsdc_U1424 ( .B1(U_dsdc_n1142), .B2(U_addrdec_n97), .A(
        U_dsdc_n1114), .ZN(U_dsdc_N416) );
  OAI211_X2 U_dsdc_U1423 ( .C1(U_dsdc_n184), .C2(U_dsdc_n445), .A(U_dsdc_n1074), .B(U_dsdc_n1497), .ZN(U_dsdc_n1077) );
  AOI211_X2 U_dsdc_U1422 ( .C1(U_dsdc_n1138), .C2(U_dsdc_n1401), .A(
        U_dsdc_n1077), .B(U_dsdc_n1149), .ZN(U_dsdc_n1078) );
  OAI21_X2 U_dsdc_U1421 ( .B1(U_dsdc_n1142), .B2(U_dsdc_n2006), .A(
        U_dsdc_n1078), .ZN(U_dsdc_N412) );
  NAND2_X2 U_dsdc_U1420 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_6_), .ZN(
        U_dsdc_n1554) );
  OAI211_X2 U_dsdc_U1419 ( .C1(U_dsdc_n1108), .C2(n91), .A(U_dsdc_n1096), .B(
        U_dsdc_n1554), .ZN(U_dsdc_n1099) );
  AOI211_X2 U_dsdc_U1418 ( .C1(U_dsdc_n1138), .C2(U_dsdc_n1404), .A(
        U_dsdc_n1099), .B(U_dsdc_n1219), .ZN(U_dsdc_n1100) );
  OAI21_X2 U_dsdc_U1417 ( .B1(U_dsdc_n1142), .B2(U_addrdec_n99), .A(
        U_dsdc_n1100), .ZN(U_dsdc_N414) );
  NOR2_X2 U_dsdc_U1416 ( .A1(U_dsdc_n696), .A2(U_dsdc_n680), .ZN(U_dsdc_n1405)
         );
  NAND2_X2 U_dsdc_U1415 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_5_), .ZN(
        U_dsdc_n1552) );
  OAI211_X2 U_dsdc_U1414 ( .C1(U_dsdc_n1108), .C2(n93), .A(U_dsdc_n1101), .B(
        U_dsdc_n1552), .ZN(U_dsdc_n1105) );
  AOI211_X2 U_dsdc_U1413 ( .C1(U_dsdc_n1138), .C2(U_dsdc_n1405), .A(
        U_dsdc_n1105), .B(U_dsdc_n1220), .ZN(U_dsdc_n1106) );
  OAI21_X2 U_dsdc_U1412 ( .B1(U_dsdc_n1142), .B2(U_addrdec_n98), .A(
        U_dsdc_n1106), .ZN(U_dsdc_N415) );
  OAI211_X2 U_dsdc_U1411 ( .C1(U_dsdc_n605), .C2(U_dsdc_n1984), .A(
        U_dsdc_n1144), .B(U_dsdc_n1070), .ZN(U_dsdc_n1071) );
  AOI21_X2 U_dsdc_U1410 ( .B1(U_dsdc_n1121), .B2(debug_ad_col_addr_10_), .A(
        U_dsdc_n1071), .ZN(U_dsdc_n1072) );
  INV_X4 U_dsdc_U1409 ( .A(U_dsdc_n1072), .ZN(U_dsdc_N409) );
  NOR2_X2 U_dsdc_U1408 ( .A1(U_dsdc_n695), .A2(U_dsdc_n694), .ZN(U_dsdc_n1402)
         );
  OAI211_X2 U_dsdc_U1407 ( .C1(U_dsdc_n962), .C2(U_dsdc_n1040), .A(U_dsdc_n961), .B(U_dsdc_n1979), .ZN(U_dsdc_i_dqs_nxt) );
  OAI21_X2 U_dsdc_U1406 ( .B1(cr_t_rp[1]), .B2(cr_t_rp[2]), .A(U_dsdc_n1334), 
        .ZN(U_dsdc_n1338) );
  AOI22_X2 U_dsdc_U1405 ( .A1(U_dsdc_n1336), .A2(cr_t_rp[0]), .B1(U_dsdc_n1335), .B2(U_dsdc_n171), .ZN(U_dsdc_n1337) );
  NAND2_X2 U_dsdc_U1404 ( .A1(U_dsdc_n1338), .A2(U_dsdc_n1337), .ZN(
        U_dsdc_rp_cnt2_nxt[0]) );
  AOI21_X2 U_dsdc_U1403 ( .B1(U_dsdc_n1810), .B2(U_dsdc_n443), .A(U_dsdc_n699), 
        .ZN(U_dsdc_n1399) );
  NOR2_X2 U_dsdc_U1402 ( .A1(U_dsdc_n698), .A2(U_dsdc_n697), .ZN(U_dsdc_n1400)
         );
  NOR3_X2 U_dsdc_U1401 ( .A1(U_dsdc_n1125), .A2(U_dsdc_n1388), .A3(
        U_dsdc_n1124), .ZN(U_dsdc_n1131) );
  NAND2_X2 U_dsdc_U1400 ( .A1(U_dsdc_n1003), .A2(U_dsdc_oldest_bank_0_), .ZN(
        U_dsdc_n1123) );
  AOI211_X2 U_dsdc_U1399 ( .C1(U_dsdc_r_bank_addr_0_), .C2(U_dsdc_n1128), .A(
        U_dsdc_n1671), .B(U_dsdc_close_bank_addr_0_), .ZN(U_dsdc_n1126) );
  INV_X4 U_dsdc_U1398 ( .A(U_dsdc_n1304), .ZN(U_dsdc_n1308) );
  OAI22_X2 U_dsdc_U1397 ( .A1(U_dsdc_n1308), .A2(U_dsdc_n1306), .B1(
        U_dsdc_n1307), .B2(U_dsdc_n1305), .ZN(U_dsdc_wr_cnt_nxt[1]) );
  OAI22_X2 U_dsdc_U1396 ( .A1(U_dsdc_n1308), .A2(cr_t_wr[0]), .B1(
        U_dsdc_wr_cnt_0_), .B2(U_dsdc_n1307), .ZN(U_dsdc_wr_cnt_nxt[0]) );
  AOI221_X2 U_dsdc_U1395 ( .B1(U_dsdc_row_cnt_0_), .B2(U_dsdc_n1791), .C1(
        U_dsdc_row_cnt_1_), .C2(U_dsdc_n1791), .A(U_dsdc_n1800), .ZN(
        U_dsdc_n1778) );
  NAND2_X2 U_dsdc_U1394 ( .A1(U_dsdc_n1778), .A2(U_dsdc_n577), .ZN(
        U_dsdc_n1774) );
  NOR4_X2 U_dsdc_U1393 ( .A1(cr_row_addr_width[2]), .A2(cr_row_addr_width[0]), 
        .A3(cr_row_addr_width[3]), .A4(U_cr_n42), .ZN(U_dsdc_N4241) );
  NOR4_X2 U_dsdc_U1392 ( .A1(cr_row_addr_width[1]), .A2(cr_row_addr_width[2]), 
        .A3(cr_row_addr_width[3]), .A4(U_cr_n21), .ZN(U_dsdc_N4240) );
  INV_X4 U_dsdc_U1391 ( .A(U_dsdc_n1578), .ZN(U_dsdc_n1757) );
  AOI22_X2 U_dsdc_U1390 ( .A1(U_dsdc_n1758), .A2(cr_ref_all_before_sr), .B1(
        U_dsdc_n1757), .B2(cr_ref_all_after_sr), .ZN(U_dsdc_n1801) );
  INV_X4 U_dsdc_U1389 ( .A(U_dsdc_n1801), .ZN(U_dsdc_n1797) );
  AOI22_X2 U_dsdc_U1388 ( .A1(U_dsdc_n1774), .A2(U_dsdc_row_cnt_3_), .B1(
        U_dsdc_num_row[3]), .B2(U_dsdc_n1797), .ZN(U_dsdc_n1775) );
  NAND2_X2 U_dsdc_U1387 ( .A1(U_dsdc_n1791), .A2(U_dsdc_n574), .ZN(U_dsdc_n582) );
  NAND2_X2 U_dsdc_U1386 ( .A1(U_dsdc_n1775), .A2(U_dsdc_n582), .ZN(U_dsdc_n375) );
  NAND2_X2 U_dsdc_U1385 ( .A1(U_dsdc_n1052), .A2(U_dsdc_n1314), .ZN(
        U_dsdc_write_start_nxt) );
  AOI21_X2 U_dsdc_U1383 ( .B1(U_dsdc_n1629), .B2(U_dsdc_n1633), .A(
        U_dsdc_n1632), .ZN(U_dsdc_n1872) );
  OAI22_X2 U_dsdc_U1382 ( .A1(U_dsdc_n1424), .A2(U_dsdc_n1633), .B1(
        U_dsdc_n1423), .B2(U_dsdc_n1629), .ZN(U_dsdc_n2070) );
  NAND2_X2 U_dsdc_U1381 ( .A1(U_dsdc_n1632), .A2(U_dsdc_n2070), .ZN(
        U_dsdc_n705) );
  AOI21_X2 U_dsdc_U1379 ( .B1(hiu_wrapped_burst), .B2(U_dsdc_n1284), .A(
        U_dsdc_n1438), .ZN(U_dsdc_n1285) );
  AOI211_X2 U_dsdc_U1378 ( .C1(U_dsdc_access_cs_4_), .C2(U_dsdc_n1383), .A(
        U_dsdc_n1288), .B(U_dsdc_n1287), .ZN(U_dsdc_n1291) );
  NAND3_X2 U_dsdc_U1377 ( .A1(U_dsdc_n1291), .A2(U_dsdc_n1290), .A3(
        U_dsdc_n1289), .ZN(U_dsdc_n[2088]) );
  NAND2_X2 U_dsdc_U1376 ( .A1(U_dsdc_n1003), .A2(U_dsdc_oldest_bank_1_), .ZN(
        U_dsdc_n1390) );
  OAI21_X2 U_dsdc_U1375 ( .B1(U_dsdc_n1391), .B2(U_dsdc_n1130), .A(
        U_dsdc_n1390), .ZN(U_dsdc_close_bank_addr_1_) );
  AOI21_X2 U_dsdc_U1374 ( .B1(U_dsdc_r_bank_addr_1_), .B2(U_dsdc_n1128), .A(
        U_dsdc_close_bank_addr_1_), .ZN(U_dsdc_n1129) );
  OAI21_X2 U_dsdc_U1373 ( .B1(U_dsdc_n1131), .B2(U_dsdc_n1130), .A(
        U_dsdc_n1129), .ZN(U_dsdc_s_bank_addr_nxt_a_1_) );
  NAND2_X2 U_dsdc_U1372 ( .A1(U_dsdc_n1152), .A2(U_cr_n58), .ZN(U_dsdc_n766)
         );
  NAND2_X2 U_dsdc_U1371 ( .A1(U_dsdc_n1344), .A2(U_dsdc_n766), .ZN(
        U_dsdc_n1359) );
  NOR4_X2 U_dsdc_U1370 ( .A1(U_dsdc_n1366), .A2(U_dsdc_n1365), .A3(
        U_dsdc_n1364), .A4(U_dsdc_n1363), .ZN(U_dsdc_n1369) );
  NAND2_X2 U_dsdc_U1369 ( .A1(U_dsdc_n767), .A2(U_dsdc_n766), .ZN(U_dsdc_n1368) );
  NAND2_X2 U_dsdc_U1368 ( .A1(U_dsdc_n1805), .A2(U_dsdc_n1367), .ZN(
        U_dsdc_n1387) );
  NAND4_X2 U_dsdc_U1367 ( .A1(U_dsdc_n1370), .A2(U_dsdc_n1369), .A3(
        U_dsdc_n1368), .A4(U_dsdc_n1387), .ZN(U_dsdc_n1371) );
  AOI21_X2 U_dsdc_U1366 ( .B1(U_dsdc_n1373), .B2(U_dsdc_n1372), .A(
        U_dsdc_n1371), .ZN(U_dsdc_n1377) );
  NAND2_X2 U_dsdc_U1365 ( .A1(U_dsdc_n899), .A2(U_dsdc_n983), .ZN(U_dsdc_n1375) );
  NAND3_X2 U_dsdc_U1364 ( .A1(U_dsdc_n1377), .A2(U_dsdc_n1376), .A3(
        U_dsdc_n1375), .ZN(U_dsdc_n[2092]) );
  OAI22_X2 U_dsdc_U1363 ( .A1(U_dsdc_n1391), .A2(U_dsdc_n600), .B1(
        U_dsdc_oldest_bank_1_), .B2(U_dsdc_n1123), .ZN(U_dsdc_bm_close_bank_1_) );
  OAI21_X2 U_dsdc_U1362 ( .B1(U_dsdc_bm_rc_cnt_0__3_), .B2(U_dsdc_n1174), .A(
        n83), .ZN(U_dsdc_n1178) );
  AOI21_X2 U_dsdc_U1361 ( .B1(U_dsdc_bm_rc_cnt_0__0_), .B2(
        U_dsdc_bm_rc_cnt_0__1_), .A(U_dsdc_n1176), .ZN(U_dsdc_n1177) );
  OAI22_X2 U_dsdc_U1359 ( .A1(U_dsdc_n1178), .A2(U_dsdc_n1177), .B1(n83), .B2(
        U_cr_n106), .ZN(U_dsdc_N4333) );
  OAI22_X2 U_dsdc_U1357 ( .A1(U_dsdc_n1178), .A2(U_dsdc_bm_rc_cnt_0__0_), .B1(
        U_cr_n64), .B2(n83), .ZN(U_dsdc_N4332) );
  OAI22_X2 U_dsdc_U1356 ( .A1(U_dsdc_n1090), .A2(U_dsdc_cas_latency_cnt_0_), 
        .B1(U_dsdc_n1393), .B2(U_dsdc_n1089), .ZN(U_dsdc_n300) );
  AOI21_X2 U_dsdc_U1355 ( .B1(U_dsdc_n1038), .B2(U_dsdc_n1037), .A(
        U_dsdc_n1293), .ZN(U_dsdc_n1251) );
  AOI21_X2 U_dsdc_U1354 ( .B1(U_dsdc_n1033), .B2(U_dsdc_n1032), .A(
        U_dsdc_n1031), .ZN(U_dsdc_n1036) );
  OAI211_X2 U_dsdc_U1353 ( .C1(U_dsdc_n1036), .C2(U_dsdc_n1035), .A(
        U_dsdc_n1411), .B(U_dsdc_n1040), .ZN(U_dsdc_n348) );
  OAI21_X2 U_dsdc_U1352 ( .B1(U_dsdc_n1251), .B2(U_dsdc_n466), .A(U_dsdc_n348), 
        .ZN(U_dsdc_n232) );
  AOI21_X2 U_dsdc_U1351 ( .B1(U_dsdc_n1867), .B2(U_dsdc_n1847), .A(
        U_dsdc_n1961), .ZN(U_dsdc_n1851) );
  OAI221_X2 U_dsdc_U1350 ( .B1(U_dsdc_bm_bank_age_2__0_), .B2(U_dsdc_n1860), 
        .C1(U_dsdc_n353), .C2(U_dsdc_n1859), .A(U_dsdc_n1851), .ZN(
        U_dsdc_n1853) );
  OAI21_X2 U_dsdc_U1349 ( .B1(U_dsdc_n178), .B2(U_dsdc_n1853), .A(U_dsdc_n1852), .ZN(U_dsdc_n1854) );
  OAI21_X2 U_dsdc_U1348 ( .B1(U_dsdc_n1859), .B2(U_dsdc_n1856), .A(
        U_dsdc_n1854), .ZN(U_dsdc_n210) );
  OAI21_X2 U_dsdc_U1347 ( .B1(U_dsdc_n1391), .B2(U_dsdc_n572), .A(U_dsdc_n1001), .ZN(U_dsdc_bm_close_bank_0_) );
  OAI21_X2 U_dsdc_U1346 ( .B1(U_dsdc_bm_rc_cnt_3__3_), .B2(U_dsdc_n1227), .A(
        U_dsdc_n313), .ZN(U_dsdc_n1233) );
  AOI21_X2 U_dsdc_U1345 ( .B1(U_dsdc_bm_rc_cnt_3__0_), .B2(
        U_dsdc_bm_rc_cnt_3__1_), .A(U_dsdc_n1229), .ZN(U_dsdc_n1231) );
  OAI22_X2 U_dsdc_U1344 ( .A1(U_dsdc_n1233), .A2(U_dsdc_n1231), .B1(
        U_dsdc_n313), .B2(U_cr_n106), .ZN(U_dsdc_N4474) );
  OAI22_X2 U_dsdc_U1343 ( .A1(U_dsdc_n1233), .A2(U_dsdc_bm_rc_cnt_3__0_), .B1(
        U_cr_n64), .B2(U_dsdc_n313), .ZN(U_dsdc_N4473) );
  INV_X4 U_dsdc_U1342 ( .A(U_dsdc_n763), .ZN(U_dsdc_n289) );
  AOI21_X2 U_dsdc_U1341 ( .B1(U_dsdc_n1791), .B2(U_dsdc_n1788), .A(
        U_dsdc_n1800), .ZN(U_dsdc_n1785) );
  NAND2_X2 U_dsdc_U1340 ( .A1(U_dsdc_n1785), .A2(U_dsdc_n578), .ZN(
        U_dsdc_n1781) );
  NAND2_X2 U_dsdc_U1339 ( .A1(cr_row_addr_width[1]), .A2(cr_row_addr_width[0]), 
        .ZN(U_dsdc_n1662) );
  NAND2_X2 U_dsdc_U1338 ( .A1(U_dsdc_n1652), .A2(cr_row_addr_width[2]), .ZN(
        U_dsdc_n1653) );
  NAND2_X2 U_dsdc_U1336 ( .A1(U_dsdc_n1653), .A2(U_cr_n70), .ZN(U_dsdc_n1656)
         );
  NAND2_X2 U_dsdc_U1335 ( .A1(U_dsdc_n1657), .A2(U_dsdc_n1656), .ZN(
        U_dsdc_n1661) );
  NOR2_X2 U_dsdc_U1334 ( .A1(U_dsdc_n1658), .A2(U_dsdc_n1661), .ZN(
        U_dsdc_N4253) );
  NOR2_X2 U_dsdc_U1333 ( .A1(U_dsdc_n1659), .A2(U_dsdc_n1661), .ZN(
        U_dsdc_N4252) );
  NOR2_X2 U_dsdc_U1332 ( .A1(U_dsdc_n1662), .A2(U_dsdc_n1661), .ZN(
        U_dsdc_N4250) );
  NOR4_X2 U_dsdc_U1331 ( .A1(cr_row_addr_width[1]), .A2(cr_row_addr_width[2]), 
        .A3(U_cr_n21), .A4(U_cr_n70), .ZN(U_dsdc_N4248) );
  NOR2_X2 U_dsdc_U1330 ( .A1(cr_row_addr_width[3]), .A2(U_dsdc_n1653), .ZN(
        U_dsdc_N4246) );
  NAND2_X2 U_dsdc_U1329 ( .A1(U_dsdc_n1657), .A2(U_dsdc_n1654), .ZN(
        U_dsdc_n1655) );
  NOR2_X2 U_dsdc_U1328 ( .A1(U_dsdc_n1659), .A2(U_dsdc_n1655), .ZN(
        U_dsdc_N4244) );
  NOR2_X2 U_dsdc_U1327 ( .A1(U_dsdc_n1662), .A2(U_dsdc_n1656), .ZN(
        U_dsdc_N4242) );
  NOR2_X2 U_dsdc_U1326 ( .A1(U_dsdc_N4242), .A2(U_dsdc_n613), .ZN(U_dsdc_n614)
         );
  NAND2_X2 U_dsdc_U1325 ( .A1(U_cr_n42), .A2(U_cr_n21), .ZN(U_dsdc_n1660) );
  NAND2_X2 U_dsdc_U1324 ( .A1(U_dsdc_n614), .A2(U_dsdc_n345), .ZN(U_dsdc_n615)
         );
  NOR2_X2 U_dsdc_U1323 ( .A1(U_dsdc_N4244), .A2(U_dsdc_n615), .ZN(U_dsdc_n616)
         );
  NAND2_X2 U_dsdc_U1322 ( .A1(U_dsdc_n616), .A2(U_dsdc_n346), .ZN(U_dsdc_n617)
         );
  NOR2_X2 U_dsdc_U1321 ( .A1(U_dsdc_N4246), .A2(U_dsdc_n617), .ZN(U_dsdc_n618)
         );
  NAND2_X2 U_dsdc_U1320 ( .A1(U_dsdc_n618), .A2(U_dsdc_n358), .ZN(U_dsdc_n606)
         );
  NOR2_X2 U_dsdc_U1319 ( .A1(U_dsdc_N4248), .A2(U_dsdc_n606), .ZN(U_dsdc_n607)
         );
  NAND2_X2 U_dsdc_U1318 ( .A1(U_dsdc_n607), .A2(U_dsdc_n357), .ZN(U_dsdc_n608)
         );
  NOR2_X2 U_dsdc_U1317 ( .A1(U_dsdc_N4250), .A2(U_dsdc_n608), .ZN(U_dsdc_n609)
         );
  NAND2_X2 U_dsdc_U1316 ( .A1(U_dsdc_n609), .A2(U_dsdc_n399), .ZN(U_dsdc_n610)
         );
  NOR2_X2 U_dsdc_U1315 ( .A1(U_dsdc_N4252), .A2(U_dsdc_n610), .ZN(U_dsdc_n611)
         );
  AOI22_X2 U_dsdc_U1314 ( .A1(U_dsdc_row_cnt_15_), .A2(U_dsdc_n1781), .B1(
        U_dsdc_num_row[15]), .B2(U_dsdc_n1797), .ZN(U_dsdc_n1782) );
  NOR3_X2 U_dsdc_U1313 ( .A1(U_dsdc_bm_bank_age_2__2_), .A2(U_dsdc_n1859), 
        .A3(U_dsdc_n1856), .ZN(U_dsdc_n1862) );
  OAI21_X2 U_dsdc_U1312 ( .B1(U_dsdc_n1868), .B2(U_dsdc_n1862), .A(U_dsdc_n459), .ZN(U_dsdc_n1863) );
  OAI21_X2 U_dsdc_U1311 ( .B1(U_dsdc_n1864), .B2(U_dsdc_n459), .A(U_dsdc_n1863), .ZN(U_dsdc_n212) );
  AOI21_X2 U_dsdc_U1310 ( .B1(U_dsdc_n1907), .B2(U_dsdc_n1888), .A(
        U_dsdc_n1961), .ZN(U_dsdc_n1891) );
  OAI221_X2 U_dsdc_U1309 ( .B1(U_dsdc_bm_bank_age_3__0_), .B2(U_dsdc_n1900), 
        .C1(U_dsdc_n304), .C2(U_dsdc_n1899), .A(U_dsdc_n1891), .ZN(
        U_dsdc_n1893) );
  OAI21_X2 U_dsdc_U1308 ( .B1(U_dsdc_n302), .B2(U_dsdc_n1893), .A(U_dsdc_n1892), .ZN(U_dsdc_n1894) );
  OAI21_X2 U_dsdc_U1307 ( .B1(U_dsdc_n1899), .B2(U_dsdc_n1896), .A(
        U_dsdc_n1894), .ZN(U_dsdc_n219) );
  AOI21_X2 U_dsdc_U1306 ( .B1(U_dsdc_n1937), .B2(U_dsdc_n1918), .A(
        U_dsdc_n1961), .ZN(U_dsdc_n1921) );
  OAI221_X2 U_dsdc_U1305 ( .B1(U_dsdc_bm_bank_age_1__0_), .B2(U_dsdc_n1930), 
        .C1(U_dsdc_n352), .C2(U_dsdc_n1929), .A(U_dsdc_n1921), .ZN(
        U_dsdc_n1923) );
  OAI21_X2 U_dsdc_U1304 ( .B1(U_dsdc_n335), .B2(U_dsdc_n1923), .A(U_dsdc_n1922), .ZN(U_dsdc_n1924) );
  OAI21_X2 U_dsdc_U1303 ( .B1(U_dsdc_n1929), .B2(U_dsdc_n1926), .A(
        U_dsdc_n1924), .ZN(U_dsdc_n224) );
  NOR2_X2 U_dsdc_U1302 ( .A1(U_dsdc_n994), .A2(U_dsdc_n2071), .ZN(U_dsdc_n704)
         );
  NOR2_X2 U_dsdc_U1301 ( .A1(U_dsdc_n1367), .A2(U_dsdc_n704), .ZN(U_dsdc_n901)
         );
  NOR3_X2 U_dsdc_U1300 ( .A1(U_dsdc_bm_bank_age_1__2_), .A2(U_dsdc_n1929), 
        .A3(U_dsdc_n1926), .ZN(U_dsdc_n1932) );
  OAI21_X2 U_dsdc_U1299 ( .B1(U_dsdc_n1938), .B2(U_dsdc_n1932), .A(U_dsdc_n460), .ZN(U_dsdc_n1933) );
  OAI21_X2 U_dsdc_U1298 ( .B1(U_dsdc_n1934), .B2(U_dsdc_n460), .A(U_dsdc_n1933), .ZN(U_dsdc_n226) );
  OAI21_X2 U_dsdc_U1297 ( .B1(U_dsdc_bm_rc_cnt_2__3_), .B2(U_dsdc_n1202), .A(
        U_dsdc_n310), .ZN(U_dsdc_n1206) );
  OAI22_X2 U_dsdc_U1296 ( .A1(U_dsdc_n1206), .A2(U_dsdc_bm_rc_cnt_2__0_), .B1(
        U_cr_n64), .B2(U_dsdc_n310), .ZN(U_dsdc_N4426) );
  OAI21_X2 U_dsdc_U1295 ( .B1(U_dsdc_bm_rc_cnt_1__3_), .B2(U_dsdc_n1188), .A(
        U_dsdc_n620), .ZN(U_dsdc_n1192) );
  AOI21_X2 U_dsdc_U1294 ( .B1(U_dsdc_bm_rc_cnt_1__0_), .B2(
        U_dsdc_bm_rc_cnt_1__1_), .A(U_dsdc_n1190), .ZN(U_dsdc_n1191) );
  OAI22_X2 U_dsdc_U1293 ( .A1(U_dsdc_n1192), .A2(U_dsdc_n1191), .B1(
        U_dsdc_n620), .B2(U_cr_n106), .ZN(U_dsdc_N4380) );
  AOI21_X2 U_dsdc_U1292 ( .B1(U_dsdc_bm_rc_cnt_2__0_), .B2(
        U_dsdc_bm_rc_cnt_2__1_), .A(U_dsdc_n1204), .ZN(U_dsdc_n1205) );
  OAI22_X2 U_dsdc_U1291 ( .A1(U_dsdc_n1206), .A2(U_dsdc_n1205), .B1(
        U_dsdc_n310), .B2(U_cr_n106), .ZN(U_dsdc_N4427) );
  OAI22_X2 U_dsdc_U1290 ( .A1(U_dsdc_n1192), .A2(U_dsdc_bm_rc_cnt_1__0_), .B1(
        U_cr_n64), .B2(U_dsdc_n620), .ZN(U_dsdc_N4379) );
  NOR4_X2 U_dsdc_U1289 ( .A1(U_dsdc_n1802), .A2(U_dsdc_n968), .A3(U_dsdc_n967), 
        .A4(U_dsdc_n360), .ZN(U_dsdc_n971) );
  AOI22_X2 U_dsdc_U1288 ( .A1(U_dsdc_n969), .A2(U_dsdc_n1038), .B1(U_dsdc_n166), .B2(U_dsdc_n1974), .ZN(U_dsdc_n970) );
  NAND3_X2 U_dsdc_U1287 ( .A1(U_dsdc_n972), .A2(U_dsdc_n971), .A3(U_dsdc_n970), 
        .ZN(U_dsdc_s_dout_valid_nxt) );
  OAI22_X2 U_dsdc_U1286 ( .A1(U_dsdc_n1252), .A2(cr_t_wtr[0]), .B1(
        U_dsdc_wtr_cnt_0_), .B2(U_dsdc_n1251), .ZN(U_dsdc_wtr_cnt_nxt[0]) );
  NAND2_X2 U_dsdc_U1285 ( .A1(n83), .A2(U_dsdc_n1181), .ZN(U_dsdc_n1185) );
  AOI21_X2 U_dsdc_U1284 ( .B1(U_dsdc_bm_ras_cnt_0__0_), .B2(
        U_dsdc_bm_ras_cnt_0__1_), .A(U_dsdc_n1183), .ZN(U_dsdc_n1184) );
  OAI22_X2 U_dsdc_U1282 ( .A1(U_dsdc_n1185), .A2(U_dsdc_n1184), .B1(n83), .B2(
        U_cr_n120), .ZN(U_dsdc_N4320) );
  OAI22_X2 U_dsdc_U1280 ( .A1(U_dsdc_n1185), .A2(U_dsdc_bm_ras_cnt_0__0_), 
        .B1(n83), .B2(n95), .ZN(U_dsdc_N4319) );
  OAI22_X2 U_dsdc_U1279 ( .A1(U_dsdc_n1252), .A2(U_dsdc_n1247), .B1(
        U_dsdc_n1251), .B2(U_dsdc_n1246), .ZN(U_dsdc_wtr_cnt_nxt[1]) );
  NAND2_X2 U_dsdc_U1278 ( .A1(cr_t_wtr[1]), .A2(cr_t_wtr[0]), .ZN(U_dsdc_n1250) );
  AOI21_X2 U_dsdc_U1277 ( .B1(U_dsdc_wtr_cnt_2_), .B2(U_dsdc_n1248), .A(
        U_dsdc_n1284), .ZN(U_dsdc_n1249) );
  OAI22_X2 U_dsdc_U1276 ( .A1(U_dsdc_n1252), .A2(U_dsdc_n1250), .B1(
        U_dsdc_n1251), .B2(U_dsdc_n1249), .ZN(U_dsdc_wtr_cnt_nxt[2]) );
  NAND2_X2 U_dsdc_U1275 ( .A1(U_dsdc_n313), .A2(U_dsdc_n1237), .ZN(
        U_dsdc_n1243) );
  AOI21_X2 U_dsdc_U1274 ( .B1(U_dsdc_bm_ras_cnt_3__0_), .B2(
        U_dsdc_bm_ras_cnt_3__1_), .A(U_dsdc_n1239), .ZN(U_dsdc_n1241) );
  AOI22_X2 U_dsdc_U1273 ( .A1(U_dsdc_num_row[2]), .A2(U_dsdc_n1797), .B1(
        U_dsdc_n325), .B2(U_dsdc_n204), .ZN(U_dsdc_n1777) );
  OAI21_X2 U_dsdc_U1272 ( .B1(U_dsdc_n1778), .B2(U_dsdc_n204), .A(U_dsdc_n1777), .ZN(U_dsdc_n374) );
  NOR3_X2 U_dsdc_U1271 ( .A1(U_dsdc_r_bm_open_bank[0]), .A2(U_dsdc_n1941), 
        .A3(U_dsdc_n384), .ZN(U_dsdc_n1972) );
  NOR3_X2 U_dsdc_U1270 ( .A1(U_dsdc_r_bm_close_bank_0_), .A2(U_dsdc_n384), 
        .A3(U_dsdc_n1942), .ZN(U_dsdc_n2081) );
  INV_X4 U_dsdc_U1269 ( .A(U_dsdc_n2081), .ZN(U_dsdc_n1965) );
  NAND2_X2 U_dsdc_U1268 ( .A1(U_dsdc_n479), .A2(U_dsdc_n478), .ZN(U_dsdc_n480)
         );
  NOR2_X2 U_dsdc_U1267 ( .A1(U_dsdc_n1945), .A2(U_dsdc_n480), .ZN(U_dsdc_n1947) );
  OAI21_X2 U_dsdc_U1263 ( .B1(U_dsdc_n1965), .B2(U_dsdc_n2080), .A(
        U_dsdc_n1956), .ZN(U_dsdc_n2083) );
  AOI221_X2 U_dsdc_U1262 ( .B1(U_dsdc_n2081), .B2(U_dsdc_bm_bank_age_0__0_), 
        .C1(U_dsdc_n1972), .C2(U_dsdc_n201), .A(U_dsdc_n2083), .ZN(
        U_dsdc_n1958) );
  NAND3_X2 U_dsdc_U1261 ( .A1(U_dsdc_n435), .A2(U_dsdc_n201), .A3(U_dsdc_n2080), .ZN(U_dsdc_n1962) );
  OAI221_X2 U_dsdc_U1260 ( .B1(U_dsdc_bm_bank_age_0__1_), .B2(U_dsdc_n1959), 
        .C1(U_dsdc_n435), .C2(U_dsdc_n1958), .A(U_dsdc_n1957), .ZN(U_dsdc_n228) );
  NOR2_X2 U_dsdc_U1259 ( .A1(U_dsdc_n939), .A2(U_dsdc_n1483), .ZN(U_dsdc_n1612) );
  NAND2_X2 U_dsdc_U1258 ( .A1(U_dsdc_n1343), .A2(U_dsdc_n651), .ZN(
        U_dsdc_n1601) );
  NOR3_X2 U_dsdc_U1257 ( .A1(U_dsdc_n1311), .A2(U_dsdc_n1336), .A3(
        U_dsdc_n1495), .ZN(U_dsdc_n1389) );
  NOR3_X2 U_dsdc_U1256 ( .A1(U_dsdc_n1383), .A2(U_dsdc_n659), .A3(U_dsdc_n1592), .ZN(U_dsdc_n1417) );
  NAND2_X2 U_dsdc_U1255 ( .A1(U_dsdc_n310), .A2(U_dsdc_n1209), .ZN(
        U_dsdc_n1213) );
  OAI22_X2 U_dsdc_U1254 ( .A1(U_dsdc_n1213), .A2(U_dsdc_bm_ras_cnt_2__0_), 
        .B1(U_dsdc_n310), .B2(n95), .ZN(U_dsdc_N4413) );
  AOI21_X2 U_dsdc_U1253 ( .B1(U_dsdc_bm_ras_cnt_2__0_), .B2(
        U_dsdc_bm_ras_cnt_2__1_), .A(U_dsdc_n1211), .ZN(U_dsdc_n1212) );
  OAI22_X2 U_dsdc_U1252 ( .A1(U_dsdc_n1213), .A2(U_dsdc_n1212), .B1(
        U_dsdc_n310), .B2(U_cr_n120), .ZN(U_dsdc_N4414) );
  NAND2_X2 U_dsdc_U1251 ( .A1(U_dsdc_n620), .A2(U_dsdc_n1195), .ZN(
        U_dsdc_n1199) );
  OAI22_X2 U_dsdc_U1250 ( .A1(U_dsdc_n1199), .A2(U_dsdc_bm_ras_cnt_1__0_), 
        .B1(U_dsdc_n620), .B2(n95), .ZN(U_dsdc_N4366) );
  AOI21_X2 U_dsdc_U1249 ( .B1(U_dsdc_bm_ras_cnt_1__0_), .B2(
        U_dsdc_bm_ras_cnt_1__1_), .A(U_dsdc_n1197), .ZN(U_dsdc_n1198) );
  OAI22_X2 U_dsdc_U1248 ( .A1(U_dsdc_n1199), .A2(U_dsdc_n1198), .B1(
        U_dsdc_n620), .B2(U_cr_n120), .ZN(U_dsdc_N4367) );
  NOR3_X2 U_dsdc_U1247 ( .A1(U_dsdc_n1534), .A2(U_dsdc_n1533), .A3(
        U_dsdc_n2055), .ZN(U_dsdc_n1541) );
  AOI211_X2 U_dsdc_U1246 ( .C1(U_dsdc_n1431), .C2(U_dsdc_n1621), .A(
        U_dsdc_n1757), .B(U_dsdc_n1538), .ZN(U_dsdc_n1539) );
  NAND2_X2 U_dsdc_U1245 ( .A1(U_dsdc_n1799), .A2(U_dsdc_n590), .ZN(
        U_dsdc_n1792) );
  AOI22_X2 U_dsdc_U1244 ( .A1(U_dsdc_row_cnt_11_), .A2(U_dsdc_n1792), .B1(
        U_dsdc_num_row[11]), .B2(U_dsdc_n1797), .ZN(U_dsdc_n1793) );
  NAND2_X2 U_dsdc_U1243 ( .A1(U_dsdc_n1793), .A2(U_dsdc_n584), .ZN(U_dsdc_n368) );
  NAND2_X2 U_dsdc_U1242 ( .A1(U_dsdc_n1767), .A2(U_dsdc_n583), .ZN(
        U_dsdc_n1763) );
  AOI22_X2 U_dsdc_U1241 ( .A1(U_dsdc_row_cnt_7_), .A2(U_dsdc_n1763), .B1(
        U_dsdc_num_row[7]), .B2(U_dsdc_n1797), .ZN(U_dsdc_n1764) );
  NAND2_X2 U_dsdc_U1240 ( .A1(U_dsdc_n1791), .A2(U_dsdc_n579), .ZN(U_dsdc_n587) );
  NAND2_X2 U_dsdc_U1239 ( .A1(U_dsdc_n1764), .A2(U_dsdc_n587), .ZN(U_dsdc_n379) );
  NAND2_X2 U_dsdc_U1238 ( .A1(U_dsdc_n1790), .A2(U_dsdc_n576), .ZN(
        U_dsdc_n1786) );
  AOI22_X2 U_dsdc_U1237 ( .A1(U_dsdc_row_cnt_13_), .A2(U_dsdc_n1786), .B1(
        U_dsdc_num_row[13]), .B2(U_dsdc_n1797), .ZN(U_dsdc_n1787) );
  NAND2_X2 U_dsdc_U1236 ( .A1(U_dsdc_n1791), .A2(U_dsdc_n585), .ZN(U_dsdc_n588) );
  NAND2_X2 U_dsdc_U1235 ( .A1(U_dsdc_n1787), .A2(U_dsdc_n588), .ZN(U_dsdc_n370) );
  NAND2_X2 U_dsdc_U1234 ( .A1(U_dsdc_n1773), .A2(U_dsdc_n591), .ZN(
        U_dsdc_n1768) );
  AOI22_X2 U_dsdc_U1233 ( .A1(U_dsdc_row_cnt_5_), .A2(U_dsdc_n1768), .B1(
        U_dsdc_num_row[5]), .B2(U_dsdc_n1797), .ZN(U_dsdc_n1769) );
  NAND2_X2 U_dsdc_U1232 ( .A1(U_dsdc_n1791), .A2(U_dsdc_n581), .ZN(U_dsdc_n586) );
  NAND2_X2 U_dsdc_U1231 ( .A1(U_dsdc_n1769), .A2(U_dsdc_n586), .ZN(U_dsdc_n377) );
  NAND2_X2 U_dsdc_U1230 ( .A1(U_dsdc_n1762), .A2(U_dsdc_n592), .ZN(
        U_dsdc_n1759) );
  AOI22_X2 U_dsdc_U1229 ( .A1(U_dsdc_row_cnt_9_), .A2(U_dsdc_n1759), .B1(
        U_dsdc_num_row[9]), .B2(U_dsdc_n1797), .ZN(U_dsdc_n1760) );
  NAND2_X2 U_dsdc_U1228 ( .A1(U_dsdc_n1760), .A2(U_dsdc_n589), .ZN(U_dsdc_n381) );
  INV_X4 U_dsdc_U1227 ( .A(U_dsdc_n1676), .ZN(U_dsdc_n1722) );
  AOI21_X2 U_dsdc_U1226 ( .B1(cr_t_init[2]), .B2(U_dsdc_n1722), .A(
        U_dsdc_n1716), .ZN(U_dsdc_n1717) );
  OAI21_X2 U_dsdc_U1225 ( .B1(U_dsdc_n468), .B2(U_dsdc_n1718), .A(U_dsdc_n1717), .ZN(U_dsdc_n405) );
  AOI21_X2 U_dsdc_U1224 ( .B1(U_dsdc_row_cnt_0_), .B2(U_dsdc_n1791), .A(
        U_dsdc_n1800), .ZN(U_dsdc_n1780) );
  AOI21_X2 U_dsdc_U1223 ( .B1(U_dsdc_n598), .B2(U_dsdc_n1797), .A(U_dsdc_n325), 
        .ZN(U_dsdc_n1779) );
  OAI21_X2 U_dsdc_U1222 ( .B1(U_dsdc_n1780), .B2(U_dsdc_n465), .A(U_dsdc_n1779), .ZN(U_dsdc_n373) );
  OAI211_X2 U_dsdc_U1221 ( .C1(U_dsdc_n1326), .C2(U_dsdc_n1322), .A(cr_t_rp[2]), .B(U_dsdc_n1321), .ZN(U_dsdc_n1324) );
  NAND2_X2 U_dsdc_U1220 ( .A1(U_dsdc_n1324), .A2(U_dsdc_n1323), .ZN(
        U_dsdc_rp_cnt2_nxt[2]) );
  NOR3_X2 U_dsdc_U1219 ( .A1(U_dsdc_bm_bank_age_3__2_), .A2(U_dsdc_n1899), 
        .A3(U_dsdc_n1896), .ZN(U_dsdc_n1902) );
  OAI21_X2 U_dsdc_U1218 ( .B1(U_dsdc_n1908), .B2(U_dsdc_n1902), .A(U_dsdc_n284), .ZN(U_dsdc_n1903) );
  OAI21_X2 U_dsdc_U1217 ( .B1(U_dsdc_n1904), .B2(U_dsdc_n284), .A(U_dsdc_n1903), .ZN(U_dsdc_n221) );
  AOI22_X2 U_dsdc_U1216 ( .A1(U_dsdc_num_row[10]), .A2(U_dsdc_n1797), .B1(
        U_dsdc_n1796), .B2(U_dsdc_n208), .ZN(U_dsdc_n1798) );
  OAI21_X2 U_dsdc_U1215 ( .B1(U_dsdc_n1799), .B2(U_dsdc_n208), .A(U_dsdc_n1798), .ZN(U_dsdc_n367) );
  AOI22_X2 U_dsdc_U1214 ( .A1(U_dsdc_num_row[6]), .A2(U_dsdc_n1797), .B1(
        U_dsdc_n593), .B2(U_dsdc_n206), .ZN(U_dsdc_n1766) );
  OAI21_X2 U_dsdc_U1213 ( .B1(U_dsdc_n1767), .B2(U_dsdc_n206), .A(U_dsdc_n1766), .ZN(U_dsdc_n378) );
  AOI22_X2 U_dsdc_U1212 ( .A1(U_dsdc_num_row[8]), .A2(U_dsdc_n1797), .B1(
        U_dsdc_n595), .B2(U_dsdc_n205), .ZN(U_dsdc_n1761) );
  OAI21_X2 U_dsdc_U1211 ( .B1(U_dsdc_n1762), .B2(U_dsdc_n205), .A(U_dsdc_n1761), .ZN(U_dsdc_n380) );
  AOI22_X2 U_dsdc_U1210 ( .A1(U_dsdc_num_row[4]), .A2(U_dsdc_n1797), .B1(
        U_dsdc_n1771), .B2(U_dsdc_n207), .ZN(U_dsdc_n1772) );
  OAI21_X2 U_dsdc_U1209 ( .B1(U_dsdc_n1773), .B2(U_dsdc_n207), .A(U_dsdc_n1772), .ZN(U_dsdc_n376) );
  AOI22_X2 U_dsdc_U1208 ( .A1(U_dsdc_num_row[14]), .A2(U_dsdc_n1797), .B1(
        U_dsdc_n1783), .B2(U_dsdc_n202), .ZN(U_dsdc_n1784) );
  OAI21_X2 U_dsdc_U1207 ( .B1(U_dsdc_n1785), .B2(U_dsdc_n202), .A(U_dsdc_n1784), .ZN(U_dsdc_n371) );
  AOI22_X2 U_dsdc_U1206 ( .A1(U_dsdc_num_row[12]), .A2(U_dsdc_n1797), .B1(
        U_dsdc_n594), .B2(U_dsdc_n203), .ZN(U_dsdc_n1789) );
  OAI21_X2 U_dsdc_U1205 ( .B1(U_dsdc_n1790), .B2(U_dsdc_n203), .A(U_dsdc_n1789), .ZN(U_dsdc_n369) );
  NAND2_X2 U_dsdc_U1204 ( .A1(U_dsdc_n1159), .A2(U_dsdc_n1152), .ZN(
        U_dsdc_n1160) );
  OAI21_X2 U_dsdc_U1203 ( .B1(U_dsdc_n1160), .B2(U_dsdc_n1158), .A(
        U_dsdc_n1157), .ZN(U_dsdc_N4282) );
  NAND2_X2 U_dsdc_U1202 ( .A1(U_dsdc_n1158), .A2(U_dsdc_bm_ras_cnt_max_2_), 
        .ZN(U_dsdc_n1154) );
  OAI21_X2 U_dsdc_U1201 ( .B1(U_dsdc_n1161), .B2(U_dsdc_n1160), .A(
        U_dsdc_n1155), .ZN(U_dsdc_N4283) );
  OAI221_X2 U_dsdc_U1200 ( .B1(U_dsdc_bm_bank_age_3__2_), .B2(U_dsdc_n1901), 
        .C1(U_dsdc_n303), .C2(U_dsdc_n1898), .A(U_dsdc_n1897), .ZN(U_dsdc_n220) );
  AOI22_X2 U_dsdc_U1199 ( .A1(U_dsdc_init_cnt_4_), .A2(U_dsdc_n1709), .B1(
        cr_t_init[4]), .B2(U_dsdc_n1722), .ZN(U_dsdc_n1710) );
  AOI22_X2 U_dsdc_U1198 ( .A1(U_dsdc_init_cnt_8_), .A2(U_dsdc_n1695), .B1(
        cr_t_init[8]), .B2(U_dsdc_n1722), .ZN(U_dsdc_n1696) );
  AOI22_X2 U_dsdc_U1197 ( .A1(U_dsdc_init_cnt_10_), .A2(U_dsdc_n1688), .B1(
        cr_t_init[10]), .B2(U_dsdc_n1722), .ZN(U_dsdc_n1689) );
  AOI22_X2 U_dsdc_U1196 ( .A1(U_dsdc_init_cnt_6_), .A2(U_dsdc_n1702), .B1(
        cr_t_init[6]), .B2(U_dsdc_n1722), .ZN(U_dsdc_n1703) );
  OAI221_X2 U_dsdc_U1195 ( .B1(U_dsdc_bm_bank_age_2__2_), .B2(U_dsdc_n1861), 
        .C1(U_dsdc_n336), .C2(U_dsdc_n1858), .A(U_dsdc_n1857), .ZN(U_dsdc_n211) );
  OAI221_X2 U_dsdc_U1194 ( .B1(U_dsdc_bm_bank_age_1__2_), .B2(U_dsdc_n1931), 
        .C1(U_dsdc_n337), .C2(U_dsdc_n1928), .A(U_dsdc_n1927), .ZN(U_dsdc_n225) );
  INV_X4 U_dsdc_U1193 ( .A(U_dsdc_n1972), .ZN(U_dsdc_n1966) );
  AOI21_X2 U_dsdc_U1192 ( .B1(U_dsdc_bm_bank_age_0__1_), .B2(
        U_dsdc_bm_bank_age_0__0_), .A(U_dsdc_n1966), .ZN(U_dsdc_n1960) );
  AOI211_X2 U_dsdc_U1191 ( .C1(U_dsdc_n2081), .C2(U_dsdc_n1962), .A(
        U_dsdc_n1961), .B(U_dsdc_n1960), .ZN(U_dsdc_n1964) );
  OAI221_X2 U_dsdc_U1190 ( .B1(U_dsdc_bm_bank_age_0__2_), .B2(U_dsdc_n1966), 
        .C1(U_dsdc_n334), .C2(U_dsdc_n1965), .A(U_dsdc_n1964), .ZN(
        U_dsdc_n1971) );
  NAND3_X2 U_dsdc_U1189 ( .A1(U_dsdc_bm_bank_age_0__1_), .A2(
        U_dsdc_bm_bank_age_0__0_), .A3(U_dsdc_n1972), .ZN(U_dsdc_n1967) );
  NOR2_X2 U_dsdc_U1188 ( .A1(U_dsdc_n334), .A2(U_dsdc_n1967), .ZN(U_dsdc_n1973) );
  NAND3_X2 U_dsdc_U1187 ( .A1(U_dsdc_n1700), .A2(U_dsdc_n1699), .A3(
        U_dsdc_n1698), .ZN(U_dsdc_n410) );
  NAND3_X2 U_dsdc_U1186 ( .A1(U_dsdc_n1693), .A2(U_dsdc_n1692), .A3(
        U_dsdc_n1691), .ZN(U_dsdc_n412) );
  NAND3_X2 U_dsdc_U1185 ( .A1(U_dsdc_n1707), .A2(U_dsdc_n1706), .A3(
        U_dsdc_n1705), .ZN(U_dsdc_n408) );
  OAI211_X2 U_dsdc_U1184 ( .C1(U_dsdc_init_cnt_2_), .C2(U_dsdc_n1711), .A(
        U_dsdc_init_cnt_3_), .B(U_dsdc_n1715), .ZN(U_dsdc_n1713) );
  NAND3_X2 U_dsdc_U1183 ( .A1(U_dsdc_n1714), .A2(U_dsdc_n1713), .A3(
        U_dsdc_n1712), .ZN(U_dsdc_n406) );
  NOR3_X2 U_dsdc_U1182 ( .A1(U_dsdc_bm_bank_age_0__2_), .A2(U_dsdc_n1965), 
        .A3(U_dsdc_n1962), .ZN(U_dsdc_n1968) );
  OAI221_X2 U_dsdc_U1181 ( .B1(U_dsdc_bm_bank_age_0__2_), .B2(U_dsdc_n1967), 
        .C1(U_dsdc_n334), .C2(U_dsdc_n1964), .A(U_dsdc_n1963), .ZN(U_dsdc_n229) );
  OAI221_X2 U_dsdc_U1180 ( .B1(U_dsdc_bm_bank_age_1__0_), .B2(U_dsdc_n1919), 
        .C1(U_dsdc_n352), .C2(U_dsdc_n1921), .A(U_dsdc_n356), .ZN(U_dsdc_n223)
         );
  OAI221_X2 U_dsdc_U1179 ( .B1(U_dsdc_bm_bank_age_3__0_), .B2(U_dsdc_n1889), 
        .C1(U_dsdc_n304), .C2(U_dsdc_n1891), .A(U_dsdc_n185), .ZN(U_dsdc_n218)
         );
  OAI21_X2 U_dsdc_U1178 ( .B1(U_dsdc_n1973), .B2(U_dsdc_n1968), .A(U_dsdc_n458), .ZN(U_dsdc_n1969) );
  OAI21_X2 U_dsdc_U1177 ( .B1(U_dsdc_n1970), .B2(U_dsdc_n458), .A(U_dsdc_n1969), .ZN(U_dsdc_n230) );
  OAI221_X2 U_dsdc_U1176 ( .B1(U_dsdc_bm_bank_age_2__0_), .B2(U_dsdc_n1848), 
        .C1(U_dsdc_n353), .C2(U_dsdc_n1851), .A(U_dsdc_n164), .ZN(U_dsdc_n209)
         );
  OAI221_X2 U_dsdc_U1175 ( .B1(U_dsdc_bm_bank_age_0__0_), .B2(U_dsdc_n2085), 
        .C1(U_dsdc_n201), .C2(U_dsdc_n2084), .A(U_dsdc_n168), .ZN(U_dsdc_n283)
         );
  AOI22_X2 U_dsdc_U1174 ( .A1(U_dsdc_init_cnt_12_), .A2(U_dsdc_n1680), .B1(
        cr_t_init[12]), .B2(U_dsdc_n1722), .ZN(U_dsdc_n1681) );
  INV_X4 U_dsdc_U1173 ( .A(U_dsdc_n765), .ZN(U_dsdc_n287) );
  AOI21_X2 U_dsdc_U1170 ( .B1(U_dsdc_n1270), .B2(hiu_burst_size[0]), .A(
        U_dsdc_n1261), .ZN(U_dsdc_n1339) );
  NAND2_X2 U_dsdc_U1169 ( .A1(U_dsdc_n1339), .A2(U_dsdc_n1281), .ZN(
        U_dsdc_n1282) );
  OAI21_X2 U_dsdc_U1168 ( .B1(U_dsdc_n1266), .B2(U_dsdc_n1263), .A(
        U_dsdc_n1262), .ZN(U_dsdc_n1279) );
  NOR2_X2 U_dsdc_U1167 ( .A1(U_dsdc_n1282), .A2(U_dsdc_n1279), .ZN(
        U_dsdc_n1278) );
  NAND2_X2 U_dsdc_U1166 ( .A1(U_dsdc_n1278), .A2(U_dsdc_n1276), .ZN(
        U_dsdc_n1273) );
  OAI21_X2 U_dsdc_U1165 ( .B1(U_dsdc_n1266), .B2(U_dmc_n16), .A(U_dsdc_n1264), 
        .ZN(U_dsdc_n1274) );
  NOR2_X2 U_dsdc_U1164 ( .A1(U_dsdc_n1273), .A2(U_dsdc_n1274), .ZN(
        U_dsdc_n1272) );
  NOR2_X2 U_dsdc_U1163 ( .A1(U_dsdc_n1271), .A2(U_dsdc_n1340), .ZN(
        U_dsdc_cas_cnt_nxt[5]) );
  AOI21_X2 U_dsdc_U1162 ( .B1(U_dsdc_n1274), .B2(U_dsdc_n1273), .A(
        U_dsdc_n1272), .ZN(U_dsdc_n1275) );
  NOR2_X2 U_dsdc_U1161 ( .A1(U_dsdc_n1275), .A2(U_dsdc_n1340), .ZN(
        U_dsdc_cas_cnt_nxt[4]) );
  OAI22_X2 U_dsdc_U1160 ( .A1(U_dsdc_n1160), .A2(U_dsdc_bm_ras_cnt_max_0_), 
        .B1(U_dsdc_n1159), .B2(n95), .ZN(U_dsdc_N4281) );
  AOI21_X2 U_dsdc_U1159 ( .B1(U_dsdc_init_cnt_1_), .B2(U_dsdc_init_cnt_0_), 
        .A(U_dsdc_n1719), .ZN(U_dsdc_n1721) );
  NAND2_X2 U_dsdc_U1158 ( .A1(cr_t_init[1]), .A2(U_dsdc_n1722), .ZN(
        U_dsdc_n1720) );
  NAND2_X2 U_dsdc_U1157 ( .A1(cr_t_init[0]), .A2(U_dsdc_n1722), .ZN(
        U_dsdc_n1723) );
  AOI211_X2 U_dsdc_U1156 ( .C1(cr_exn_mode_value[10]), .C2(U_dsdc_n1671), .A(
        U_dsdc_n1618), .B(U_dsdc_n1322), .ZN(U_dsdc_n1029) );
  NAND2_X2 U_dsdc_U1155 ( .A1(U_dsdc_n1030), .A2(U_dsdc_n1029), .ZN(
        U_dsdc_N410) );
  NOR3_X2 U_dsdc_U1154 ( .A1(U_dsdc_n1491), .A2(U_dsdc_n1490), .A3(
        U_dsdc_n1521), .ZN(ctl_mode_reg_done) );
  NOR3_X2 U_dsdc_U1153 ( .A1(U_dsdc_n1491), .A2(U_dsdc_n1506), .A3(
        U_dsdc_n1521), .ZN(ctl_ext_mode_reg_done) );
  NOR2_X2 U_dsdc_U1152 ( .A1(U_dsdc_n1277), .A2(U_dsdc_n1340), .ZN(
        U_dsdc_cas_cnt_nxt[3]) );
  AOI21_X2 U_dsdc_U1151 ( .B1(U_dsdc_n1279), .B2(U_dsdc_n1282), .A(
        U_dsdc_n1278), .ZN(U_dsdc_n1280) );
  NOR2_X2 U_dsdc_U1150 ( .A1(U_dsdc_n1280), .A2(U_dsdc_n1340), .ZN(
        U_dsdc_cas_cnt_nxt[2]) );
  AOI21_X2 U_dsdc_U1149 ( .B1(U_dsdc_n1414), .B2(U_dsdc_n1419), .A(
        U_dsdc_n1629), .ZN(U_dsdc_n1630) );
  AOI211_X2 U_dsdc_U1148 ( .C1(U_dsdc_n1632), .C2(U_dsdc_n1420), .A(
        U_dsdc_n1631), .B(U_dsdc_n1630), .ZN(U_dsdc_n1635) );
  NOR3_X2 U_dsdc_U1147 ( .A1(U_dsdc_n1414), .A2(U_dsdc_n1633), .A3(
        U_dsdc_n1632), .ZN(U_dsdc_n1648) );
  OAI21_X2 U_dsdc_U1146 ( .B1(U_dsdc_n1424), .B2(U_dsdc_n1635), .A(
        U_dsdc_n1634), .ZN(U_dsdc_n1639) );
  NAND2_X2 U_dsdc_U1145 ( .A1(U_dsdc_n1414), .A2(U_dsdc_n1872), .ZN(
        U_dsdc_n1636) );
  INV_X4 U_dsdc_U1144 ( .A(U_dsdc_n1636), .ZN(U_dsdc_n1642) );
  NOR2_X2 U_dsdc_U1143 ( .A1(U_dsdc_n1639), .A2(U_dsdc_n1642), .ZN(
        U_dsdc_n1646) );
  AOI22_X2 U_dsdc_U1142 ( .A1(U_dsdc_n1642), .A2(U_dsdc_n1641), .B1(
        U_dsdc_n1640), .B2(U_dsdc_n1639), .ZN(U_dsdc_n1643) );
  OAI21_X2 U_dsdc_U1141 ( .B1(U_dsdc_n1646), .B2(U_dsdc_n200), .A(U_dsdc_n1643), .ZN(U_dsdc_n1647) );
  NOR2_X2 U_dsdc_U1140 ( .A1(U_dsdc_n1876), .A2(U_dsdc_n1359), .ZN(
        U_dsdc_n1379) );
  NOR3_X2 U_dsdc_U1137 ( .A1(U_dsdc_n1444), .A2(U_dsdc_n1640), .A3(
        U_dsdc_n1636), .ZN(U_dsdc_n1649) );
  OAI21_X2 U_dsdc_U1136 ( .B1(U_dsdc_n1419), .B2(U_dsdc_n2069), .A(
        U_dsdc_n1398), .ZN(U_dsdc_n2073) );
  INV_X4 U_dsdc_U1135 ( .A(U_dsdc_n901), .ZN(U_dsdc_n708) );
  NOR2_X2 U_dsdc_U1134 ( .A1(U_dsdc_n708), .A2(U_dsdc_n1416), .ZN(U_dsdc_n1875) );
  NOR2_X2 U_dsdc_U1133 ( .A1(U_dsdc_n461), .A2(U_dsdc_n1881), .ZN(U_dsdc_n1880) );
  AOI21_X2 U_dsdc_U1132 ( .B1(U_dsdc_n1425), .B2(U_dsdc_n1871), .A(
        U_dsdc_n2073), .ZN(U_dsdc_n2072) );
  OAI21_X2 U_dsdc_U1129 ( .B1(U_dsdc_delta_delay_0_), .B2(U_dsdc_n1875), .A(
        U_dsdc_n183), .ZN(U_dsdc_n1879) );
  AOI21_X2 U_dsdc_U1128 ( .B1(U_dsdc_n1874), .B2(U_dsdc_n464), .A(U_dsdc_n1879), .ZN(U_dsdc_n1878) );
  NAND2_X2 U_dsdc_U1127 ( .A1(U_dsdc_delta_delay_1_), .A2(U_dsdc_n1880), .ZN(
        U_dsdc_n1877) );
  AOI22_X2 U_dsdc_U1126 ( .A1(U_dsdc_delta_delay_2_), .A2(U_dsdc_n1878), .B1(
        U_dsdc_n1877), .B2(U_dsdc_n467), .ZN(U_dsdc_n214) );
  AOI211_X2 U_dsdc_U1125 ( .C1(U_dsdc_n1487), .C2(U_dsdc_operation_cs_0_), .A(
        U_dsdc_n1429), .B(U_dsdc_n1486), .ZN(U_dsdc_n1488) );
  AOI21_X2 U_dsdc_U1124 ( .B1(U_dsdc_n1638), .B2(U_dsdc_n1639), .A(
        U_dsdc_n1649), .ZN(U_dsdc_n1645) );
  NOR2_X2 U_dsdc_U1123 ( .A1(U_dsdc_n1359), .A2(U_dsdc_n1414), .ZN(U_dsdc_n770) );
  AOI211_X2 U_dsdc_U1121 ( .C1(U_dsdc_n1427), .C2(U_dsdc_n1975), .A(
        U_dsdc_n1425), .B(U_dsdc_n1974), .ZN(U_dsdc_n1976) );
  NAND3_X2 U_dsdc_U1120 ( .A1(U_dsdc_n869), .A2(U_dsdc_n1397), .A3(
        U_dsdc_n1976), .ZN(U_dsdc_n713) );
  NOR2_X2 U_dsdc_U1119 ( .A1(U_dsdc_n713), .A2(U_dsdc_n1802), .ZN(U_dsdc_n1396) );
  INV_X4 U_dsdc_U1118 ( .A(U_dsdc_n956), .ZN(U_dsdc_n718) );
  NAND2_X2 U_dsdc_U1117 ( .A1(U_dsdc_n1396), .A2(U_dsdc_n718), .ZN(
        U_dsdc_n2067) );
  NOR2_X2 U_dsdc_U1116 ( .A1(U_dsdc_n2067), .A2(U_dsdc_n1411), .ZN(
        U_dsdc_n1395) );
  NAND2_X2 U_dsdc_U1115 ( .A1(U_dsdc_n1347), .A2(U_dsdc_n1346), .ZN(
        U_dsdc_n280) );
  AOI22_X2 U_dsdc_U1114 ( .A1(U_dsdc_N2002), .A2(U_dsdc_n1379), .B1(
        U_dsdc_r_cas_latency_3_), .B2(U_dsdc_n770), .ZN(U_dsdc_n773) );
  NAND2_X2 U_dsdc_U1113 ( .A1(n89), .A2(U_dsdc_N1990), .ZN(U_dsdc_n772) );
  OAI211_X2 U_dsdc_U1112 ( .C1(U_dsdc_n1645), .C2(U_dsdc_n1644), .A(
        U_dsdc_n773), .B(U_dsdc_n772), .ZN(U_dsdc_n774) );
  AOI21_X2 U_dsdc_U1111 ( .B1(U_dsdc_n1647), .B2(U_dsdc_term_cnt_3_), .A(
        U_dsdc_n774), .ZN(U_dsdc_n775) );
  INV_X4 U_dsdc_U1110 ( .A(U_dsdc_n775), .ZN(U_dsdc_term_cnt_nxt[3]) );
  NAND2_X2 U_dsdc_U1109 ( .A1(U_dsdc_n1674), .A2(U_dsdc_n1673), .ZN(
        U_dsdc_n418) );
  NAND2_X2 U_dsdc_U1108 ( .A1(U_dsdc_n879), .A2(U_dsdc_n759), .ZN(U_dsdc_n717)
         );
  AOI22_X2 U_dsdc_U1107 ( .A1(debug_ad_col_addr_2_), .A2(U_dsdc_n2048), .B1(
        U_dsdc_r_col_addr_2_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n1992) );
  OAI21_X2 U_dsdc_U1106 ( .B1(U_dsdc_n1994), .B2(U_dsdc_n1993), .A(
        U_dsdc_n1992), .ZN(U_dsdc_n241) );
  INV_X4 U_dsdc_U1105 ( .A(U_dsdc_n2048), .ZN(U_dsdc_n2010) );
  AOI22_X2 U_dsdc_U1104 ( .A1(U_dsdc_n1405), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_5_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n1999) );
  OAI21_X2 U_dsdc_U1103 ( .B1(U_addrdec_n98), .B2(U_dsdc_n2010), .A(
        U_dsdc_n1999), .ZN(U_dsdc_n244) );
  AOI22_X2 U_dsdc_U1102 ( .A1(debug_ad_col_addr_10_), .A2(U_dsdc_n2048), .B1(
        U_dsdc_r_col_addr_10_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n1983) );
  OAI21_X2 U_dsdc_U1101 ( .B1(U_dsdc_n1994), .B2(U_dsdc_n1984), .A(
        U_dsdc_n1983), .ZN(U_dsdc_n234) );
  AOI22_X2 U_dsdc_U1100 ( .A1(U_dsdc_n1404), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_6_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n2001) );
  OAI21_X2 U_dsdc_U1099 ( .B1(U_addrdec_n99), .B2(U_dsdc_n2010), .A(
        U_dsdc_n2001), .ZN(U_dsdc_n245) );
  AOI22_X2 U_dsdc_U1098 ( .A1(U_dsdc_n1407), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_13_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n1988) );
  OAI21_X2 U_dsdc_U1097 ( .B1(debug_ad_col_addr_13_), .B2(U_dsdc_n2010), .A(
        U_dsdc_n1988), .ZN(U_dsdc_n237) );
  AOI22_X2 U_dsdc_U1096 ( .A1(U_dsdc_n1402), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_9_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n2009) );
  OAI21_X2 U_dsdc_U1095 ( .B1(U_addrdec_n61), .B2(U_dsdc_n2010), .A(
        U_dsdc_n2009), .ZN(U_dsdc_n248) );
  AOI22_X2 U_dsdc_U1094 ( .A1(U_dsdc_n1401), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_8_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n2005) );
  OAI21_X2 U_dsdc_U1093 ( .B1(U_dsdc_n2006), .B2(U_dsdc_n2010), .A(
        U_dsdc_n2005), .ZN(U_dsdc_n247) );
  AOI22_X2 U_dsdc_U1092 ( .A1(U_dsdc_n1399), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_3_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n1995) );
  OAI21_X2 U_dsdc_U1091 ( .B1(U_addrdec_n9), .B2(U_dsdc_n2010), .A(
        U_dsdc_n1995), .ZN(U_dsdc_n242) );
  AOI22_X2 U_dsdc_U1090 ( .A1(U_dsdc_n1400), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_7_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n2003) );
  OAI21_X2 U_dsdc_U1089 ( .B1(U_addrdec_n100), .B2(U_dsdc_n2010), .A(
        U_dsdc_n2003), .ZN(U_dsdc_n246) );
  OAI21_X2 U_dsdc_U1088 ( .B1(U_dsdc_n1994), .B2(U_dsdc_n1986), .A(
        U_dsdc_n1985), .ZN(U_dsdc_n235) );
  AOI22_X2 U_dsdc_U1087 ( .A1(U_dsdc_n1406), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_4_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n1997) );
  OAI21_X2 U_dsdc_U1086 ( .B1(U_addrdec_n97), .B2(U_dsdc_n2010), .A(
        U_dsdc_n1997), .ZN(U_dsdc_n243) );
  AOI22_X2 U_dsdc_U1085 ( .A1(U_dsdc_N1685), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_0_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n1981) );
  OAI21_X2 U_dsdc_U1084 ( .B1(U_dsdc_n1982), .B2(U_dsdc_n2010), .A(
        U_dsdc_n1981), .ZN(U_dsdc_n233) );
  AOI22_X2 U_dsdc_U1083 ( .A1(U_dsdc_n1408), .A2(U_dsdc_n2008), .B1(
        U_dsdc_r_col_addr_12_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n1987) );
  OAI21_X2 U_dsdc_U1082 ( .B1(U_dsdc_n1994), .B2(U_dsdc_n1990), .A(
        U_dsdc_n1989), .ZN(U_dsdc_n238) );
  NOR2_X2 U_dsdc_U1081 ( .A1(U_dsdc_n1341), .A2(U_dsdc_n1340), .ZN(
        U_dsdc_cas_cnt_nxt[0]) );
  NAND3_X2 U_dsdc_U1080 ( .A1(U_dsdc_n717), .A2(U_dsdc_n675), .A3(U_dsdc_n674), 
        .ZN(U_dsdc_n676) );
  AOI22_X2 U_dsdc_U1079 ( .A1(U_dsdc_n1408), .A2(U_dsdc_n1817), .B1(
        U_dsdc_r_col_addr_12_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1547) );
  AOI22_X2 U_dsdc_U1078 ( .A1(U_dsdc_n1407), .A2(U_dsdc_n1817), .B1(
        U_dsdc_r_col_addr_13_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1548) );
  OAI21_X2 U_dsdc_U1077 ( .B1(debug_ad_col_addr_13_), .B2(U_dsdc_n1819), .A(
        U_dsdc_n1548), .ZN(U_dsdc_i_col_addr_nxt[13]) );
  AOI22_X2 U_dsdc_U1076 ( .A1(U_dsdc_xsr_cnt_4_), .A2(U_dsdc_n1741), .B1(
        cr_t_xsr[4]), .B2(U_dsdc_n1754), .ZN(U_dsdc_n1742) );
  OAI21_X2 U_dsdc_U1075 ( .B1(U_dsdc_xsr_cnt_4_), .B2(U_dsdc_n1744), .A(
        U_dsdc_n1742), .ZN(U_dsdc_n390) );
  AOI22_X2 U_dsdc_U1074 ( .A1(debug_ad_col_addr_5_), .A2(U_dsdc_n1815), .B1(
        U_dsdc_n1405), .B2(U_dsdc_n1817), .ZN(U_dsdc_n1553) );
  NAND2_X2 U_dsdc_U1073 ( .A1(U_dsdc_n1553), .A2(U_dsdc_n1552), .ZN(
        U_dsdc_i_col_addr_nxt[5]) );
  AOI22_X2 U_dsdc_U1072 ( .A1(debug_ad_col_addr_4_), .A2(U_dsdc_n1815), .B1(
        U_dsdc_n1406), .B2(U_dsdc_n1817), .ZN(U_dsdc_n1551) );
  NAND2_X2 U_dsdc_U1071 ( .A1(U_dsdc_n1551), .A2(U_dsdc_n1550), .ZN(
        U_dsdc_i_col_addr_nxt[4]) );
  AOI22_X2 U_dsdc_U1070 ( .A1(debug_ad_col_addr_1_), .A2(U_dsdc_n1815), .B1(
        U_dsdc_n354), .B2(U_dsdc_n1817), .ZN(U_dsdc_n1813) );
  NAND2_X2 U_dsdc_U1069 ( .A1(U_dsdc_n1813), .A2(U_dsdc_n1812), .ZN(
        U_dsdc_n319) );
  AOI22_X2 U_dsdc_U1068 ( .A1(debug_ad_col_addr_6_), .A2(U_dsdc_n1815), .B1(
        U_dsdc_n1404), .B2(U_dsdc_n1817), .ZN(U_dsdc_n1555) );
  NAND2_X2 U_dsdc_U1067 ( .A1(U_dsdc_n1555), .A2(U_dsdc_n1554), .ZN(
        U_dsdc_i_col_addr_nxt[6]) );
  NOR2_X2 U_dsdc_U1066 ( .A1(U_dsdc_n719), .A2(U_dsdc_n881), .ZN(U_dsdc_n2018)
         );
  OAI22_X2 U_dsdc_U1065 ( .A1(U_dsdc_n2020), .A2(U_dsdc_n2015), .B1(
        U_dsdc_n2018), .B2(U_dsdc_n469), .ZN(U_dsdc_n249) );
  OAI22_X2 U_dsdc_U1064 ( .A1(U_dsdc_n2020), .A2(U_dsdc_n2017), .B1(
        U_dsdc_n2018), .B2(U_dsdc_n471), .ZN(U_dsdc_n251) );
  OAI22_X2 U_dsdc_U1063 ( .A1(U_dsdc_n2020), .A2(U_dsdc_n2016), .B1(
        U_dsdc_n2018), .B2(U_dsdc_n470), .ZN(U_dsdc_n250) );
  OAI22_X2 U_dsdc_U1062 ( .A1(U_dsdc_n2020), .A2(U_dsdc_n2019), .B1(
        U_dsdc_n2018), .B2(U_dsdc_n472), .ZN(U_dsdc_n252) );
  NOR2_X2 U_dsdc_U1061 ( .A1(U_dsdc_xsr_cnt_0_), .A2(U_dsdc_xsr_cnt_1_), .ZN(
        U_dsdc_n1747) );
  NAND2_X2 U_dsdc_U1060 ( .A1(U_dsdc_n1747), .A2(U_dsdc_n1750), .ZN(
        U_dsdc_n1751) );
  NOR2_X2 U_dsdc_U1059 ( .A1(U_dsdc_n1747), .A2(U_dsdc_n1756), .ZN(
        U_dsdc_n1748) );
  AOI22_X2 U_dsdc_U1058 ( .A1(U_dsdc_xsr_cnt_2_), .A2(U_dsdc_n1748), .B1(
        cr_t_xsr[2]), .B2(U_dsdc_n1754), .ZN(U_dsdc_n1749) );
  OAI21_X2 U_dsdc_U1057 ( .B1(U_dsdc_xsr_cnt_2_), .B2(U_dsdc_n1751), .A(
        U_dsdc_n1749), .ZN(U_dsdc_n388) );
  AOI22_X2 U_dsdc_U1056 ( .A1(U_dsdc_n1401), .A2(U_dsdc_n1817), .B1(
        U_dsdc_r_col_addr_8_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1807) );
  OAI21_X2 U_dsdc_U1055 ( .B1(U_dsdc_n1819), .B2(U_dsdc_n2006), .A(
        U_dsdc_n1807), .ZN(U_dsdc_n323) );
  AOI22_X2 U_dsdc_U1054 ( .A1(U_dsdc_N1685), .A2(U_dsdc_n1817), .B1(
        U_dsdc_r_col_addr_0_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1818) );
  OAI21_X2 U_dsdc_U1053 ( .B1(U_dsdc_n1819), .B2(U_dsdc_n1982), .A(
        U_dsdc_n1818), .ZN(U_dsdc_n315) );
  AOI22_X2 U_dsdc_U1052 ( .A1(U_dsdc_n1402), .A2(U_dsdc_n1817), .B1(
        U_dsdc_r_col_addr_9_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1806) );
  OAI21_X2 U_dsdc_U1051 ( .B1(U_dsdc_n1819), .B2(U_addrdec_n61), .A(
        U_dsdc_n1806), .ZN(U_dsdc_n324) );
  AOI22_X2 U_dsdc_U1050 ( .A1(U_dsdc_n1399), .A2(U_dsdc_n1817), .B1(
        U_dsdc_r_col_addr_3_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1809) );
  OAI21_X2 U_dsdc_U1049 ( .B1(U_dsdc_n1819), .B2(U_addrdec_n9), .A(
        U_dsdc_n1809), .ZN(U_dsdc_n321) );
  AOI22_X2 U_dsdc_U1048 ( .A1(U_dsdc_n1400), .A2(U_dsdc_n1817), .B1(
        U_dsdc_r_col_addr_7_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1808) );
  OAI21_X2 U_dsdc_U1047 ( .B1(U_dsdc_n1819), .B2(U_addrdec_n100), .A(
        U_dsdc_n1808), .ZN(U_dsdc_n322) );
  AOI22_X2 U_dsdc_U1046 ( .A1(debug_ad_row_addr[11]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_11_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2025) );
  INV_X4 U_dsdc_U1045 ( .A(U_dsdc_n2025), .ZN(U_dsdc_n257) );
  AOI22_X2 U_dsdc_U1044 ( .A1(debug_ad_row_addr[10]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_10_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2024) );
  INV_X4 U_dsdc_U1043 ( .A(U_dsdc_n2024), .ZN(U_dsdc_n256) );
  AOI22_X2 U_dsdc_U1042 ( .A1(debug_ad_row_addr[0]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_0_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2023) );
  INV_X4 U_dsdc_U1041 ( .A(U_dsdc_n2023), .ZN(U_dsdc_n255) );
  AOI22_X2 U_dsdc_U1040 ( .A1(debug_ad_row_addr[15]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_15_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2029) );
  INV_X4 U_dsdc_U1039 ( .A(U_dsdc_n2029), .ZN(U_dsdc_n261) );
  AOI22_X2 U_dsdc_U1038 ( .A1(debug_ad_row_addr[1]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_1_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2030) );
  INV_X4 U_dsdc_U1037 ( .A(U_dsdc_n2030), .ZN(U_dsdc_n262) );
  AOI22_X2 U_dsdc_U1036 ( .A1(debug_ad_row_addr[2]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_2_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2031) );
  INV_X4 U_dsdc_U1035 ( .A(U_dsdc_n2031), .ZN(U_dsdc_n263) );
  AOI22_X2 U_dsdc_U1034 ( .A1(debug_ad_row_addr[3]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_3_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2032) );
  INV_X4 U_dsdc_U1033 ( .A(U_dsdc_n2032), .ZN(U_dsdc_n264) );
  AOI22_X2 U_dsdc_U1032 ( .A1(debug_ad_row_addr[4]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_4_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2033) );
  INV_X4 U_dsdc_U1031 ( .A(U_dsdc_n2033), .ZN(U_dsdc_n265) );
  AOI22_X2 U_dsdc_U1030 ( .A1(debug_ad_row_addr[14]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_14_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2028) );
  INV_X4 U_dsdc_U1029 ( .A(U_dsdc_n2028), .ZN(U_dsdc_n260) );
  AOI22_X2 U_dsdc_U1028 ( .A1(debug_ad_row_addr[6]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_6_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2035) );
  INV_X4 U_dsdc_U1027 ( .A(U_dsdc_n2035), .ZN(U_dsdc_n267) );
  AOI22_X2 U_dsdc_U1026 ( .A1(debug_ad_row_addr[8]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_8_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2037) );
  INV_X4 U_dsdc_U1025 ( .A(U_dsdc_n2037), .ZN(U_dsdc_n269) );
  AOI22_X2 U_dsdc_U1024 ( .A1(debug_ad_row_addr[9]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_9_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2040) );
  INV_X4 U_dsdc_U1023 ( .A(U_dsdc_n2040), .ZN(U_dsdc_n270) );
  AOI22_X2 U_dsdc_U1022 ( .A1(debug_ad_row_addr[12]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_12_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2026) );
  INV_X4 U_dsdc_U1021 ( .A(U_dsdc_n2026), .ZN(U_dsdc_n258) );
  AOI22_X2 U_dsdc_U1020 ( .A1(debug_ad_row_addr[5]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_5_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2034) );
  INV_X4 U_dsdc_U1019 ( .A(U_dsdc_n2034), .ZN(U_dsdc_n266) );
  AOI22_X2 U_dsdc_U1018 ( .A1(debug_ad_row_addr[13]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_13_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2027) );
  INV_X4 U_dsdc_U1017 ( .A(U_dsdc_n2027), .ZN(U_dsdc_n259) );
  AOI22_X2 U_dsdc_U1016 ( .A1(debug_ad_row_addr[7]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_row_addr_7_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2036) );
  INV_X4 U_dsdc_U1015 ( .A(U_dsdc_n2036), .ZN(U_dsdc_n268) );
  AOI22_X2 U_dsdc_U1014 ( .A1(U_dsdc_delta_delay_0_), .A2(U_dsdc_n183), .B1(
        U_dsdc_n1881), .B2(U_dsdc_n461), .ZN(U_dsdc_n216) );
  NOR3_X2 U_dsdc_U1013 ( .A1(U_dsdc_n1416), .A2(U_dsdc_n1412), .A3(
        U_dsdc_n2070), .ZN(U_dsdc_n2075) );
  NAND2_X2 U_dsdc_U1012 ( .A1(U_dsdc_n2041), .A2(U_dsdc_n1396), .ZN(
        U_dsdc_n2049) );
  NOR4_X2 U_dsdc_U1011 ( .A1(U_dsdc_mrd_cnt_0_), .A2(U_dsdc_n1430), .A3(
        U_dsdc_n1671), .A4(U_dsdc_n1670), .ZN(U_dsdc_N4174) );
  AOI211_X2 U_dsdc_U1010 ( .C1(U_dsdc_mrd_cnt_1_), .C2(U_dsdc_mrd_cnt_0_), .A(
        U_dsdc_n1671), .B(U_dsdc_n1670), .ZN(U_dsdc_n1672) );
  INV_X4 U_dsdc_U1009 ( .A(U_dsdc_n1672), .ZN(U_dsdc_n423) );
  AOI22_X2 U_dsdc_U1008 ( .A1(U_dsdc_n1395), .A2(U_dsdc_n1438), .B1(
        U_dsdc_n166), .B2(U_dsdc_n2068), .ZN(U_dsdc_n279) );
  NAND3_X2 U_dsdc_U1007 ( .A1(U_dsdc_n1746), .A2(U_dsdc_n1745), .A3(
        U_dsdc_n1744), .ZN(U_dsdc_n389) );
  NAND2_X2 U_dsdc_U1006 ( .A1(U_dsdc_n1739), .A2(U_dsdc_n1738), .ZN(
        U_dsdc_n391) );
  OAI21_X2 U_dsdc_U1005 ( .B1(U_dsdc_n2079), .B2(U_dsdc_n2078), .A(
        U_dsdc_n2077), .ZN(U_dsdc_n282) );
  NAND3_X2 U_dsdc_U1004 ( .A1(U_dsdc_n1753), .A2(U_dsdc_n1752), .A3(
        U_dsdc_n1751), .ZN(U_dsdc_n387) );
  NAND2_X2 U_dsdc_U1003 ( .A1(U_dsdc_n1729), .A2(U_dsdc_n1750), .ZN(
        U_dsdc_n1734) );
  NAND2_X2 U_dsdc_U1002 ( .A1(U_dsdc_n1735), .A2(U_dsdc_n1734), .ZN(
        U_dsdc_n392) );
  NOR2_X2 U_dsdc_U1001 ( .A1(U_dsdc_n1592), .A2(U_dsdc_n1591), .ZN(
        U_dsdc_n1597) );
  INV_X4 U_dsdc_U1000 ( .A(U_dsdc_n1597), .ZN(U_dsdc_n1609) );
  NAND2_X2 U_dsdc_U999 ( .A1(U_dsdc_rcar_cnt2_3_), .A2(U_dsdc_n1609), .ZN(
        U_dsdc_n1615) );
  NAND2_X2 U_dsdc_U998 ( .A1(U_cr_n127), .A2(U_cr_n151), .ZN(U_dsdc_n1603) );
  NAND2_X2 U_dsdc_U997 ( .A1(U_cr_n151), .A2(U_cr_n104), .ZN(U_dsdc_n1593) );
  OAI21_X2 U_dsdc_U996 ( .B1(cr_t_rcar[3]), .B2(U_dsdc_n1593), .A(U_dsdc_n1612), .ZN(U_dsdc_n1596) );
  INV_X4 U_dsdc_U995 ( .A(U_dsdc_n1596), .ZN(U_dsdc_n1602) );
  AOI21_X2 U_dsdc_U994 ( .B1(U_dsdc_n1603), .B2(U_dsdc_n1602), .A(U_dsdc_n1601), .ZN(U_dsdc_n1610) );
  AOI21_X2 U_dsdc_U993 ( .B1(U_dsdc_n1612), .B2(cr_t_rcar[2]), .A(U_dsdc_n1611), .ZN(U_dsdc_n1614) );
  OAI22_X2 U_dsdc_U992 ( .A1(U_dsdc_n1616), .A2(U_dsdc_n1615), .B1(
        U_dsdc_n1614), .B2(U_cr_n72), .ZN(U_dsdc_rcar_cnt2_nxt[3]) );
  NAND2_X2 U_dsdc_U991 ( .A1(U_dsdc_n1568), .A2(U_dsdc_n1580), .ZN(
        U_dsdc_n1573) );
  NOR3_X2 U_dsdc_U990 ( .A1(U_dsdc_num_init_ref_cnt_0_), .A2(
        U_dsdc_num_init_ref_cnt_1_), .A3(U_dsdc_n2063), .ZN(U_dsdc_n1666) );
  AOI22_X2 U_dsdc_U989 ( .A1(U_dsdc_num_init_ref_cnt_2_), .A2(U_dsdc_n1571), 
        .B1(U_dsdc_n1667), .B2(cr_num_init_ref[2]), .ZN(U_dsdc_n1572) );
  OAI21_X2 U_dsdc_U988 ( .B1(U_dsdc_num_init_ref_cnt_2_), .B2(U_dsdc_n1573), 
        .A(U_dsdc_n1572), .ZN(U_dsdc_num_init_ref_cnt_nxt[2]) );
  NOR2_X2 U_dsdc_U987 ( .A1(U_dsdc_rcar_cnt2_1_), .A2(U_dsdc_rcar_cnt2_0_), 
        .ZN(U_dsdc_n1604) );
  OAI221_X2 U_dsdc_U986 ( .B1(cr_t_rcar[2]), .B2(U_dsdc_n1608), .C1(U_cr_n104), 
        .C2(U_dsdc_n1610), .A(U_dsdc_n1606), .ZN(U_dsdc_rcar_cnt2_nxt[2]) );
  AOI21_X2 U_dsdc_U985 ( .B1(U_dsdc_n1666), .B2(U_dsdc_n473), .A(U_dsdc_n2051), 
        .ZN(U_dsdc_n1668) );
  AOI22_X2 U_dsdc_U984 ( .A1(U_dsdc_num_init_ref_cnt_3_), .A2(U_dsdc_n1668), 
        .B1(U_dsdc_n1667), .B2(cr_num_init_ref[3]), .ZN(U_dsdc_n1669) );
  INV_X4 U_dsdc_U983 ( .A(U_dsdc_n1669), .ZN(U_dsdc_n431) );
  AOI22_X2 U_dsdc_U982 ( .A1(cr_t_rcar[0]), .A2(U_dsdc_n1601), .B1(
        U_dsdc_n1602), .B2(U_cr_n127), .ZN(U_dsdc_n1594) );
  OAI221_X2 U_dsdc_U981 ( .B1(U_dsdc_n1604), .B2(U_dsdc_rcar_cnt2_0_), .C1(
        U_dsdc_n1604), .C2(U_dsdc_rcar_cnt2_1_), .A(U_dsdc_n1609), .ZN(
        U_dsdc_n1598) );
  OAI211_X2 U_dsdc_U980 ( .C1(U_dsdc_n1600), .C2(U_cr_n151), .A(U_dsdc_n1608), 
        .B(U_dsdc_n1598), .ZN(U_dsdc_rcar_cnt2_nxt[1]) );
  OAI21_X2 U_dsdc_U979 ( .B1(U_dsdc_num_init_ref_cnt_0_), .B2(U_dsdc_n1567), 
        .A(U_dsdc_n1566), .ZN(U_dsdc_num_init_ref_cnt_nxt[0]) );
  NAND2_X2 U_dsdc_U978 ( .A1(U_dsdc_n1726), .A2(U_dsdc_n1725), .ZN(U_dsdc_n394) );
  NAND3_X2 U_dsdc_U977 ( .A1(U_dsdc_n1570), .A2(U_dsdc_n1573), .A3(
        U_dsdc_n1569), .ZN(U_dsdc_num_init_ref_cnt_nxt[1]) );
  INV_X4 U_dsdc_U976 ( .A(U_dsdc_n1618), .ZN(U_dsdc_n1622) );
  NOR2_X2 U_dsdc_U975 ( .A1(U_dsdc_rp_cnt1_1_), .A2(U_dsdc_rp_cnt1_0_), .ZN(
        U_dsdc_n1624) );
  AOI21_X2 U_dsdc_U974 ( .B1(U_dsdc_rp_cnt1_0_), .B2(U_dsdc_rp_cnt1_1_), .A(
        U_dsdc_n1624), .ZN(U_dsdc_n1620) );
  OAI22_X2 U_dsdc_U973 ( .A1(U_dsdc_n1622), .A2(U_cr_n147), .B1(U_dsdc_n1620), 
        .B2(U_dsdc_n1619), .ZN(U_dsdc_rp_cnt1_nxt[1]) );
  NAND2_X2 U_dsdc_U972 ( .A1(U_dsdc_rp_cnt1_2_), .A2(U_dsdc_n1621), .ZN(
        U_dsdc_n1623) );
  OAI22_X2 U_dsdc_U971 ( .A1(U_dsdc_n1624), .A2(U_dsdc_n1623), .B1(
        U_dsdc_n1622), .B2(U_cr_n148), .ZN(U_dsdc_rp_cnt1_nxt[2]) );
  OAI22_X2 U_dsdc_U970 ( .A1(U_dsdc_rp_cnt1_0_), .A2(U_dsdc_n1619), .B1(
        U_dsdc_n1622), .B2(U_cr_n45), .ZN(U_dsdc_rp_cnt1_nxt[0]) );
  NOR2_X2 U_dsdc_U969 ( .A1(U_dsdc_access_cs_3_), .A2(U_dsdc_access_cs_1_), 
        .ZN(U_dsdc_n1445) );
  NOR2_X4 U_dsdc_U968 ( .A1(debug_ad_bank_addr[1]), .A2(debug_ad_bank_addr[0]), 
        .ZN(U_dsdc_n998) );
  OAI21_X2 U_dsdc_U967 ( .B1(U_dsdc_n1428), .B2(debug_ref_req), .A(
        U_dsdc_n2056), .ZN(U_dsdc_n1473) );
  AOI222_X2 U_dsdc_U965 ( .A1(U_dsdc_n1917), .A2(U_dsdc_n349), .B1(
        U_dsdc_n1917), .B2(U_dsdc_n1954), .C1(U_dsdc_n349), .C2(U_dsdc_n1954), 
        .ZN(U_dsdc_n1920) );
  NAND2_X2 U_dsdc_U964 ( .A1(U_dsdc_n903), .A2(U_dsdc_n1411), .ZN(U_dsdc_n1315) );
  NOR2_X1 U_dsdc_U963 ( .A1(U_dsdc_n1557), .A2(hiu_rw), .ZN(U_dsdc_n883) );
  INV_X1 U_dsdc_U962 ( .A(U_dsdc_n884), .ZN(U_dsdc_n885) );
  AOI211_X2 U_dsdc_U961 ( .C1(ad_sdram_chip_select_0_), .C2(U_dsdc_n850), .A(
        U_dsdc_n849), .B(U_dsdc_n899), .ZN(U_dsdc_n851) );
  OAI211_X1 U_dsdc_U960 ( .C1(U_dsdc_n1043), .C2(U_dsdc_n914), .A(U_dsdc_n913), 
        .B(U_dsdc_n912), .ZN(U_dsdc_n925) );
  NAND3_X1 U_dsdc_U959 ( .A1(U_dsdc_n1166), .A2(U_dsdc_bm_num_open_bank_0_), 
        .A3(U_dsdc_n180), .ZN(U_dsdc_n1008) );
  OAI22_X2 U_dsdc_U958 ( .A1(debug_ref_req), .A2(U_dsdc_n1537), .B1(
        U_dsdc_n1492), .B2(U_dsdc_n2063), .ZN(U_dsdc_n1493) );
  OAI21_X2 U_dsdc_U957 ( .B1(U_dsdc_n1508), .B2(U_dsdc_n432), .A(U_dsdc_n1507), 
        .ZN(U_dsdc_n1527) );
  INV_X1 U_dsdc_U956 ( .A(U_dsdc_n1320), .ZN(U_dsdc_n1125) );
  INV_X1 U_dsdc_U955 ( .A(U_dsdc_n1286), .ZN(U_dsdc_n1373) );
  NOR4_X2 U_dsdc_U954 ( .A1(U_dsdc_init_cnt_0_), .A2(U_dsdc_init_cnt_1_), .A3(
        U_dsdc_init_cnt_2_), .A4(U_dsdc_n1724), .ZN(U_dsdc_n1716) );
  INV_X1 U_dsdc_U953 ( .A(U_dsdc_n1679), .ZN(U_dsdc_n1686) );
  AOI22_X2 U_dsdc_U952 ( .A1(U_dsdc_n1268), .A2(U_dsdc_cas_cnt_4_), .B1(
        U_dsdc_r_burst_size_4_), .B2(U_dsdc_n1269), .ZN(U_dsdc_n1264) );
  AOI22_X1 U_dsdc_U950 ( .A1(debug_ad_bank_addr[0]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_bank_addr_0_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2021) );
  NAND2_X2 U_dsdc_U949 ( .A1(U_dsdc_n891), .A2(U_dsdc_n1412), .ZN(U_dsdc_n974)
         );
  OAI222_X2 U_dsdc_U929 ( .A1(U_dsdc_n182), .A2(U_dsdc_n1258), .B1(U_dsdc_n347), .B2(U_dsdc_n601), .C1(U_dsdc_n1546), .C2(U_dsdc_n1253), .ZN(
        U_dsdc_DP_OP_1642_126_2028_I5_0_) );
  INV_X1 U_dsdc_U928 ( .A(U_dsdc_n998), .ZN(U_dsdc_n572) );
  INV_X1 U_dsdc_U926 ( .A(U_dsdc_n981), .ZN(U_dsdc_n820) );
  OAI21_X1 U_dsdc_U925 ( .B1(U_dsdc_n914), .B2(U_dsdc_n932), .A(U_dsdc_n824), 
        .ZN(U_dsdc_n849) );
  AOI21_X1 U_dsdc_U924 ( .B1(U_dsdc_n910), .B2(U_dsdc_n976), .A(U_dsdc_n836), 
        .ZN(U_dsdc_n848) );
  INV_X1 U_dsdc_U923 ( .A(U_dsdc_n1776), .ZN(U_dsdc_n574) );
  INV_X1 U_dsdc_U922 ( .A(debug_ad_bank_addr[1]), .ZN(U_dsdc_n1130) );
  INV_X1 U_dsdc_U921 ( .A(U_dsdc_n1794), .ZN(U_dsdc_n580) );
  INV_X1 U_dsdc_U920 ( .A(U_dsdc_n1765), .ZN(U_dsdc_n579) );
  INV_X1 U_dsdc_U919 ( .A(U_dsdc_n1770), .ZN(U_dsdc_n581) );
  INV_X1 U_dsdc_U918 ( .A(U_dsdc_n1795), .ZN(U_dsdc_n575) );
  NOR2_X2 U_dsdc_U917 ( .A1(U_dsdc_n716), .A2(U_dsdc_n676), .ZN(U_dsdc_n2041)
         );
  AOI22_X1 U_dsdc_U916 ( .A1(debug_ad_bank_addr[1]), .A2(U_dsdc_n2039), .B1(
        U_dsdc_r_bank_addr_1_), .B2(U_dsdc_n2038), .ZN(U_dsdc_n2022) );
  NAND2_X1 U_dsdc_U915 ( .A1(U_dsdc_n167), .A2(U_dsdc_n1445), .ZN(U_dsdc_n666)
         );
  NAND2_X2 U_dsdc_U914 ( .A1(U_dsdc_n1422), .A2(U_dsdc_n1384), .ZN(
        U_dsdc_n1136) );
  INV_X4 U_dsdc_U913 ( .A(U_dsdc_n184), .ZN(U_dsdc_n619) );
  AOI21_X2 U_dsdc_U912 ( .B1(U_dsdc_n1260), .B2(U_dsdc_n1068), .A(U_dsdc_n354), 
        .ZN(U_dsdc_n1138) );
  OAI21_X2 U_dsdc_U911 ( .B1(U_dsdc_n643), .B2(U_dsdc_n1509), .A(U_dsdc_n1513), 
        .ZN(U_dsdc_n1671) );
  NOR4_X2 U_dsdc_U910 ( .A1(U_dsdc_n1411), .A2(U_dsdc_n1427), .A3(U_dsdc_n1418), .A4(U_dsdc_n1802), .ZN(U_dsdc_n1804) );
  INV_X1 U_dsdc_U909 ( .A(debug_ad_col_addr_8_), .ZN(U_dsdc_n2006) );
  NOR4_X1 U_dsdc_U908 ( .A1(cr_row_addr_width[1]), .A2(cr_row_addr_width[0]), 
        .A3(cr_row_addr_width[2]), .A4(cr_row_addr_width[3]), .ZN(U_dsdc_N4239) );
  OAI22_X1 U_dsdc_U907 ( .A1(U_dsdc_n1391), .A2(U_dsdc_n987), .B1(U_dsdc_n999), 
        .B2(U_dsdc_n1390), .ZN(U_dsdc_bm_close_bank_3_) );
  OAI22_X1 U_dsdc_U906 ( .A1(U_dsdc_n1391), .A2(U_dsdc_n599), .B1(
        U_dsdc_oldest_bank_0_), .B2(U_dsdc_n1390), .ZN(U_dsdc_bm_close_bank_2_) );
  AOI21_X1 U_dsdc_U905 ( .B1(U_dsdc_n1791), .B2(U_dsdc_n1795), .A(U_dsdc_n1800), .ZN(U_dsdc_n1799) );
  AOI21_X1 U_dsdc_U904 ( .B1(U_dsdc_n1791), .B2(U_dsdc_n1770), .A(U_dsdc_n1800), .ZN(U_dsdc_n1767) );
  AOI21_X1 U_dsdc_U903 ( .B1(U_dsdc_n1791), .B2(U_dsdc_n1794), .A(U_dsdc_n1800), .ZN(U_dsdc_n1790) );
  AOI21_X1 U_dsdc_U902 ( .B1(U_dsdc_n1791), .B2(U_dsdc_n1776), .A(U_dsdc_n1800), .ZN(U_dsdc_n1773) );
  AOI21_X1 U_dsdc_U901 ( .B1(U_dsdc_n1791), .B2(U_dsdc_n1765), .A(U_dsdc_n1800), .ZN(U_dsdc_n1762) );
  INV_X4 U_dsdc_U900 ( .A(U_dsdc_n1724), .ZN(U_dsdc_n1715) );
  AOI21_X2 U_dsdc_U899 ( .B1(U_dsdc_n2014), .B2(U_dsdc_n2013), .A(U_dsdc_n2067), .ZN(U_dsdc_n2039) );
  OAI21_X2 U_dsdc_U898 ( .B1(U_dsdc_n891), .B2(U_dsdc_n1309), .A(U_dsdc_n720), 
        .ZN(U_dsdc_n2038) );
  OAI221_X2 U_dsdc_U897 ( .B1(U_dsdc_n1616), .B2(U_dsdc_rcar_cnt2_2_), .C1(
        U_dsdc_n1616), .C2(U_dsdc_n1605), .A(U_dsdc_n1609), .ZN(U_dsdc_n1606)
         );
  INV_X1 U_dsdc_U896 ( .A(U_dsdc_n1625), .ZN(U_dsdc_n1626) );
  NOR2_X2 U_dsdc_U895 ( .A1(U_dsdc_n667), .A2(U_dsdc_n666), .ZN(U_dsdc_n1412)
         );
  NAND2_X2 U_dsdc_U894 ( .A1(U_dsdc_n998), .A2(U_dsdc_bm_row_addr_0__6_), .ZN(
        U_dsdc_n501) );
  NOR2_X2 U_dsdc_U893 ( .A1(U_dsdc_n903), .A2(U_dsdc_n759), .ZN(U_dsdc_n891)
         );
  NOR2_X1 U_dsdc_U892 ( .A1(U_dsdc_n741), .A2(U_dsdc_access_cs_0_), .ZN(
        U_dsdc_n1416) );
  NAND4_X2 U_dsdc_U891 ( .A1(U_dsdc_n167), .A2(U_dsdc_access_cs_2_), .A3(
        U_dsdc_access_cs_0_), .A4(U_dsdc_n1445), .ZN(U_dsdc_n1633) );
  NAND3_X1 U_dsdc_U890 ( .A1(cr_do_self_ref_rp), .A2(U_dsdc_n1478), .A3(
        U_dsdc_n1577), .ZN(U_dsdc_n2062) );
  AOI22_X2 U_dsdc_U889 ( .A1(U_dsdc_bm_bank_status_0_), .A2(U_dsdc_n2082), 
        .B1(U_dsdc_n2081), .B2(U_dsdc_n2080), .ZN(U_dsdc_n2085) );
  AOI21_X2 U_dsdc_U888 ( .B1(U_dsdc_n720), .B2(U_dsdc_n1413), .A(U_dsdc_n1395), 
        .ZN(U_dsdc_n719) );
  AOI22_X2 U_dsdc_U887 ( .A1(U_dsdc_n1736), .A2(U_dsdc_n1750), .B1(cr_t_xsr[5]), .B2(U_dsdc_n1754), .ZN(U_dsdc_n1739) );
  NAND2_X1 U_dsdc_U886 ( .A1(U_dsdc_n964), .A2(U_dsdc_n167), .ZN(U_dsdc_n2014)
         );
  AOI21_X2 U_dsdc_U884 ( .B1(U_dsdc_n976), .B2(U_dsdc_n988), .A(U_dsdc_n1546), 
        .ZN(U_dsdc_n977) );
  NAND2_X1 U_dsdc_U883 ( .A1(U_dsdc_n196), .A2(U_dsdc_n432), .ZN(U_dsdc_n641)
         );
  AOI21_X1 U_dsdc_U882 ( .B1(U_dsdc_n1318), .B2(U_dsdc_access_cs_3_), .A(
        U_dsdc_n1317), .ZN(U_dsdc_n1319) );
  NAND2_X2 U_dsdc_U881 ( .A1(U_dsdc_n1676), .A2(U_dsdc_n1675), .ZN(
        U_dsdc_n1724) );
  AOI22_X2 U_dsdc_U880 ( .A1(U_dsdc_bm_bank_status_3_), .A2(U_dsdc_n2082), 
        .B1(U_dsdc_n1907), .B2(U_dsdc_n1890), .ZN(U_dsdc_n1889) );
  AOI21_X2 U_dsdc_U879 ( .B1(U_dsdc_n1977), .B2(U_dsdc_n2014), .A(U_dsdc_n2012), .ZN(U_dsdc_n2048) );
  AOI21_X2 U_dsdc_U878 ( .B1(U_dsdc_n1410), .B2(U_dsdc_n1413), .A(U_dsdc_n2039), .ZN(U_dsdc_n2020) );
  NOR2_X2 U_dsdc_U877 ( .A1(U_dsdc_n692), .A2(U_dsdc_n711), .ZN(U_dsdc_n1411)
         );
  AOI211_X2 U_dsdc_U876 ( .C1(U_dsdc_n984), .C2(U_dsdc_n986), .A(U_dsdc_n911), 
        .B(U_dsdc_n910), .ZN(U_dsdc_n912) );
  OAI21_X2 U_dsdc_U875 ( .B1(U_dsdc_n1391), .B2(U_dsdc_n1127), .A(U_dsdc_n1123), .ZN(U_dsdc_close_bank_addr_0_) );
  NAND2_X2 U_dsdc_U874 ( .A1(U_dsdc_n1708), .A2(U_dsdc_n1715), .ZN(
        U_dsdc_n1712) );
  NAND2_X2 U_dsdc_U873 ( .A1(U_dsdc_n1701), .A2(U_dsdc_n1715), .ZN(
        U_dsdc_n1705) );
  AOI22_X2 U_dsdc_U872 ( .A1(debug_ad_col_addr_11_), .A2(U_dsdc_n2048), .B1(
        U_dsdc_r_col_addr_11_), .B2(U_dsdc_n2007), .ZN(U_dsdc_n1985) );
  NOR2_X1 U_dsdc_U871 ( .A1(U_dsdc_n712), .A2(U_dsdc_n170), .ZN(U_dsdc_n871)
         );
  NAND2_X1 U_dsdc_U870 ( .A1(U_dsdc_n871), .A2(U_dsdc_n355), .ZN(U_dsdc_n1650)
         );
  NAND2_X2 U_dsdc_U869 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__11_), 
        .ZN(U_dsdc_n789) );
  NAND2_X2 U_dsdc_U868 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__15_), 
        .ZN(U_dsdc_n782) );
  NOR2_X1 U_dsdc_U867 ( .A1(U_dsdc_n936), .A2(U_dsdc_n935), .ZN(U_dsdc_n1059)
         );
  NAND3_X1 U_dsdc_U866 ( .A1(U_dsdc_n173), .A2(U_dsdc_n167), .A3(
        U_dsdc_access_cs_1_), .ZN(U_dsdc_n660) );
  NAND2_X2 U_dsdc_U865 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__5_), .ZN(
        U_dsdc_n792) );
  NAND2_X2 U_dsdc_U864 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__6_), .ZN(
        U_dsdc_n500) );
  AOI22_X2 U_dsdc_U863 ( .A1(U_dsdc_bm_bank_status_1_), .A2(U_dsdc_n2082), 
        .B1(U_dsdc_n1937), .B2(U_dsdc_n1920), .ZN(U_dsdc_n1919) );
  AOI222_X4 U_dsdc_U862 ( .A1(U_dsdc_DP_OP_1642_126_2028_n85), .A2(
        U_dsdc_data_cnt_1_), .B1(U_dsdc_n751), .B2(U_dsdc_r_burst_size_1_), 
        .C1(U_dsdc_n983), .C2(hiu_burst_size[1]), .ZN(U_dsdc_n752) );
  NAND2_X4 U_dsdc_U861 ( .A1(U_dsdc_n670), .A2(U_dsdc_n1038), .ZN(U_dsdc_n1546) );
  INV_X8 U_dsdc_U860 ( .A(U_dsdc_RSOP_1683_C2_CONTROL1), .ZN(U_dsdc_n601) );
  AOI22_X1 U_dsdc_U859 ( .A1(U_dsdc_RSOP_1683_C2_CONTROL1), .A2(
        U_dsdc_data_cnt_4_), .B1(U_dsdc_n751), .B2(U_dsdc_r_burst_size_4_), 
        .ZN(U_dsdc_n748) );
  NAND2_X4 U_dsdc_U858 ( .A1(U_dsdc_n1391), .A2(U_dsdc_n1004), .ZN(
        U_dsdc_n1326) );
  NAND2_X4 U_dsdc_U857 ( .A1(U_dsdc_n981), .A2(U_dsdc_n980), .ZN(U_dsdc_n1391)
         );
  NAND2_X1 U_dsdc_U855 ( .A1(U_dsdc_n992), .A2(U_dsdc_n991), .ZN(U_dsdc_n1386)
         );
  OAI211_X1 U_dsdc_U854 ( .C1(U_dsdc_n991), .C2(U_dsdc_n860), .A(U_dsdc_n944), 
        .B(U_dsdc_n859), .ZN(U_dsdc_n877) );
  NAND3_X1 U_dsdc_U853 ( .A1(U_dsdc_n1978), .A2(U_dsdc_n991), .A3(U_dsdc_n974), 
        .ZN(U_dsdc_dqs_mask_end_nxt) );
  NAND2_X2 U_dsdc_U852 ( .A1(U_dsdc_n936), .A2(U_dsdc_n1312), .ZN(U_dsdc_n738)
         );
  NAND2_X1 U_dsdc_U851 ( .A1(U_dsdc_n1558), .A2(U_dsdc_n181), .ZN(U_dsdc_n933)
         );
  NAND2_X1 U_dsdc_U850 ( .A1(U_dsdc_n1410), .A2(U_dsdc_n1558), .ZN(
        U_dsdc_n1651) );
  NOR3_X1 U_dsdc_U849 ( .A1(U_dsdc_n1558), .A2(U_dsdc_n1557), .A3(U_dsdc_n1556), .ZN(U_dsdc_n1563) );
  AOI211_X1 U_dsdc_U848 ( .C1(U_dsdc_n1558), .C2(U_dsdc_n724), .A(U_dsdc_n723), 
        .B(U_dsdc_n722), .ZN(U_dsdc_n727) );
  NOR2_X1 U_dsdc_U847 ( .A1(U_dsdc_n1558), .A2(U_dsdc_n165), .ZN(U_dsdc_n1413)
         );
  AOI22_X4 U_dsdc_U846 ( .A1(U_dsdc_DP_OP_1642_126_2028_n5), .A2(
        U_dsdc_DP_OP_1642_126_2028_n14), .B1(U_dsdc_DP_OP_1642_126_2028_n60), 
        .B2(U_dsdc_DP_OP_1642_126_2028_n19), .ZN(U_dsdc_DP_OP_1642_126_2028_n4) );
  AOI22_X4 U_dsdc_U845 ( .A1(U_dsdc_DP_OP_1642_126_2028_n7), .A2(
        U_dsdc_DP_OP_1642_126_2028_n15), .B1(U_dsdc_DP_OP_1642_126_2028_n59), 
        .B2(U_dsdc_DP_OP_1642_126_2028_n20), .ZN(U_dsdc_DP_OP_1642_126_2028_n6) );
  AOI22_X2 U_dsdc_U844 ( .A1(U_dsdc_DP_OP_1642_126_2028_n13), .A2(
        U_dsdc_DP_OP_1642_126_2028_n3), .B1(U_dsdc_DP_OP_1642_126_2028_n61), 
        .B2(U_dsdc_DP_OP_1642_126_2028_n85), .ZN(U_dsdc_DP_OP_1642_126_2028_n2) );
  XNOR2_X2 U_dsdc_U843 ( .A(U_dsdc_DP_OP_1642_126_2028_n86), .B(
        U_dsdc_DP_OP_1642_126_2028_n85), .ZN(U_dsdc_n162) );
  XNOR2_X2 U_dsdc_U842 ( .A(U_dsdc_n162), .B(U_dsdc_DP_OP_1642_126_2028_n85), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n11) );
  INV_X2 U_dsdc_U841 ( .A(s_rd_ready), .ZN(U_dsdc_n1484) );
  NAND2_X1 U_dsdc_U840 ( .A1(U_dsdc_bm_ras_cnt_max_0_), .A2(
        U_dsdc_bm_ras_cnt_max_1_), .ZN(U_dsdc_n1156) );
  NOR3_X2 U_dsdc_U839 ( .A1(U_dsdc_operation_cs_3_), .A2(
        U_dsdc_operation_cs_2_), .A3(U_dsdc_n432), .ZN(U_dsdc_n1512) );
  NAND2_X1 U_dsdc_U837 ( .A1(U_dsdc_n354), .A2(cr_delayed_precharge), .ZN(
        U_dsdc_n855) );
  NAND3_X2 U_dsdc_U836 ( .A1(U_dsdc_n298), .A2(U_dsdc_n167), .A3(
        U_dsdc_access_cs_3_), .ZN(U_dsdc_n692) );
  NOR2_X2 U_dsdc_U834 ( .A1(U_dsdc_n355), .A2(U_dsdc_n170), .ZN(U_dsdc_n1458)
         );
  NOR2_X1 U_dsdc_U833 ( .A1(U_dsdc_num_init_ref_cnt_0_), .A2(
        U_dsdc_num_init_ref_cnt_1_), .ZN(U_dsdc_n1568) );
  NAND2_X1 U_dsdc_U832 ( .A1(U_dsdc_n306), .A2(U_dsdc_data_flag), .ZN(
        U_dsdc_n739) );
  OR2_X1 U_dsdc_U831 ( .A1(U_dsdc_term_cnt_3_), .A2(U_dsdc_term_cnt_2_), .ZN(
        U_dsdc_n1644) );
  OR4_X2 U_dsdc_U830 ( .A1(U_dsdc_cas_cnt_5_), .A2(U_dsdc_cas_cnt_3_), .A3(
        U_dsdc_cas_cnt_4_), .A4(U_dsdc_cas_cnt_1_), .ZN(U_dsdc_n1446) );
  NAND3_X2 U_dsdc_U829 ( .A1(U_dsdc_n167), .A2(U_dsdc_access_cs_3_), .A3(
        U_dsdc_access_cs_1_), .ZN(U_dsdc_n712) );
  OR4_X2 U_dsdc_U828 ( .A1(U_dsdc_r_bm_close_bank_2_), .A2(
        U_dsdc_r_bm_close_bank_0_), .A3(U_dsdc_r_bm_close_bank_1_), .A4(
        U_dsdc_r_bm_close_bank_3_), .ZN(U_dsdc_n1846) );
  NAND2_X2 U_dsdc_U825 ( .A1(U_dsdc_n170), .A2(U_dsdc_access_cs_2_), .ZN(
        U_dsdc_n667) );
  NOR3_X2 U_dsdc_U824 ( .A1(U_dsdc_rcar_cnt2_2_), .A2(U_dsdc_rcar_cnt2_1_), 
        .A3(U_dsdc_rcar_cnt2_0_), .ZN(U_dsdc_n1616) );
  NAND2_X2 U_dsdc_U820 ( .A1(U_dsdc_n355), .A2(U_dsdc_n170), .ZN(U_dsdc_n711)
         );
  NAND2_X2 U_dsdc_U819 ( .A1(U_dsdc_operation_cs_1_), .A2(
        U_dsdc_operation_cs_0_), .ZN(U_dsdc_n1522) );
  OR4_X2 U_dsdc_U818 ( .A1(U_dsdc_row_cnt_0_), .A2(U_dsdc_row_cnt_1_), .A3(
        U_dsdc_row_cnt_2_), .A4(U_dsdc_row_cnt_3_), .ZN(U_dsdc_n1776) );
  NAND3_X2 U_dsdc_U815 ( .A1(U_dsdc_operation_cs_3_), .A2(
        U_dsdc_operation_cs_2_), .A3(U_dsdc_n432), .ZN(U_dsdc_n1485) );
  NAND2_X2 U_dsdc_U814 ( .A1(U_dsdc_n343), .A2(U_dsdc_n344), .ZN(U_dsdc_n1490)
         );
  NOR2_X2 U_dsdc_U813 ( .A1(U_dsdc_operation_cs_1_), .A2(U_dsdc_n344), .ZN(
        U_dsdc_n1435) );
  NAND2_X2 U_dsdc_U812 ( .A1(U_dsdc_operation_cs_1_), .A2(U_dsdc_n344), .ZN(
        U_dsdc_n1455) );
  NAND3_X2 U_dsdc_U811 ( .A1(U_dsdc_operation_cs_3_), .A2(U_dsdc_n432), .A3(
        U_dsdc_n341), .ZN(U_dsdc_n1451) );
  XNOR2_X1 U_dsdc_U810 ( .A(U_dsdc_n195), .B(U_dsdc_wr_cnt_0_), .ZN(
        U_dsdc_n1305) );
  AND2_X2 U_dsdc_U808 ( .A1(U_dsdc_n1842), .A2(U_dsdc_bm_bank_age_0__2_), .ZN(
        U_dsdc_n308) );
  INV_X1 U_dsdc_U807 ( .A(U_dsdc_n1583), .ZN(U_dsdc_n1585) );
  INV_X1 U_dsdc_U806 ( .A(U_dsdc_n1189), .ZN(U_dsdc_n1190) );
  OAI21_X1 U_dsdc_U805 ( .B1(U_dsdc_n171), .B2(U_dsdc_n309), .A(U_dsdc_n1329), 
        .ZN(U_dsdc_n1330) );
  INV_X2 U_dsdc_U804 ( .A(U_dsdc_n1509), .ZN(U_dsdc_n1431) );
  OAI21_X1 U_dsdc_U803 ( .B1(U_dsdc_i_col_addr_1_), .B2(U_dsdc_i_col_addr_2_), 
        .A(U_dsdc_n1810), .ZN(U_dsdc_n1993) );
  INV_X1 U_dsdc_U802 ( .A(U_dsdc_n1153), .ZN(U_dsdc_n1158) );
  INV_X1 U_dsdc_U801 ( .A(U_dsdc_n1196), .ZN(U_dsdc_n1197) );
  INV_X2 U_dsdc_U800 ( .A(U_dsdc_n1522), .ZN(U_dsdc_n642) );
  INV_X1 U_dsdc_U799 ( .A(U_dsdc_n1747), .ZN(U_dsdc_n1743) );
  INV_X2 U_dsdc_U798 ( .A(U_dsdc_n1841), .ZN(U_dsdc_n476) );
  NAND2_X1 U_dsdc_U797 ( .A1(n90), .A2(s_cas_latency[1]), .ZN(U_dsdc_n1460) );
  OR4_X2 U_dsdc_U796 ( .A1(cr_row_addr_width[2]), .A2(cr_row_addr_width[0]), 
        .A3(U_cr_n42), .A4(U_cr_n70), .ZN(U_dsdc_n357) );
  INV_X1 U_dsdc_U795 ( .A(U_dsdc_n692), .ZN(U_dsdc_n657) );
  NAND3_X1 U_dsdc_U794 ( .A1(U_dsdc_n687), .A2(U_dsdc_n172), .A3(U_dsdc_n301), 
        .ZN(U_dsdc_n688) );
  INV_X2 U_dsdc_U793 ( .A(U_dsdc_n1455), .ZN(U_dsdc_n661) );
  INV_X1 U_dsdc_U792 ( .A(U_dsdc_n1719), .ZN(U_dsdc_n1711) );
  INV_X1 U_dsdc_U791 ( .A(U_dsdc_n1210), .ZN(U_dsdc_n1211) );
  INV_X1 U_dsdc_U790 ( .A(U_dsdc_n1490), .ZN(U_dsdc_n645) );
  NOR2_X2 U_dsdc_U789 ( .A1(U_dsdc_n649), .A2(U_dsdc_access_cs_1_), .ZN(
        U_dsdc_n1427) );
  INV_X1 U_dsdc_U788 ( .A(U_dsdc_n1082), .ZN(U_dsdc_n1087) );
  NAND2_X1 U_dsdc_U787 ( .A1(U_dsdc_n1638), .A2(U_dsdc_n1637), .ZN(
        U_dsdc_n1641) );
  INV_X1 U_dsdc_U786 ( .A(U_dsdc_n1203), .ZN(U_dsdc_n1204) );
  INV_X2 U_dsdc_U785 ( .A(U_dsdc_n1419), .ZN(U_dsdc_n1632) );
  INV_X1 U_dsdc_U784 ( .A(U_dsdc_n712), .ZN(U_dsdc_n915) );
  INV_X1 U_dsdc_U783 ( .A(U_dsdc_n711), .ZN(U_dsdc_n652) );
  INV_X2 U_dsdc_U782 ( .A(U_dsdc_n1458), .ZN(U_dsdc_n658) );
  INV_X1 U_dsdc_U781 ( .A(U_dsdc_n660), .ZN(U_dsdc_n654) );
  INV_X2 U_dsdc_U780 ( .A(U_dsdc_n1436), .ZN(U_dsdc_n1465) );
  INV_X1 U_dsdc_U779 ( .A(U_dsdc_n1175), .ZN(U_dsdc_n1176) );
  INV_X1 U_dsdc_U778 ( .A(U_dsdc_n1228), .ZN(U_dsdc_n1229) );
  INV_X2 U_dsdc_U777 ( .A(U_dsdc_n1604), .ZN(U_dsdc_n1605) );
  NAND2_X1 U_dsdc_U776 ( .A1(cr_row_addr_width[1]), .A2(U_cr_n21), .ZN(
        U_dsdc_n1658) );
  OR3_X2 U_dsdc_U775 ( .A1(U_dsdc_row_cnt_5_), .A2(U_dsdc_row_cnt_4_), .A3(
        U_dsdc_n1776), .ZN(U_dsdc_n1770) );
  INV_X1 U_dsdc_U774 ( .A(U_dsdc_n1485), .ZN(U_dsdc_n1487) );
  INV_X2 U_dsdc_U773 ( .A(U_dsdc_n1662), .ZN(U_dsdc_n1652) );
  OR4_X2 U_dsdc_U772 ( .A1(cr_row_addr_width[1]), .A2(cr_row_addr_width[0]), 
        .A3(cr_row_addr_width[2]), .A4(U_cr_n70), .ZN(U_dsdc_n358) );
  INV_X1 U_dsdc_U771 ( .A(U_dsdc_n1238), .ZN(U_dsdc_n1239) );
  NOR2_X1 U_dsdc_U770 ( .A1(U_dsdc_n1040), .A2(n84), .ZN(U_dsdc_n714) );
  NAND2_X1 U_dsdc_U769 ( .A1(cr_row_addr_width[0]), .A2(U_cr_n42), .ZN(
        U_dsdc_n1659) );
  INV_X1 U_dsdc_U768 ( .A(U_dsdc_n1182), .ZN(U_dsdc_n1183) );
  OAI22_X1 U_dsdc_U767 ( .A1(U_dsdc_n1163), .A2(U_dsdc_n1165), .B1(U_dsdc_n326), .B2(U_dsdc_n174), .ZN(U_dsdc_n1162) );
  INV_X1 U_dsdc_U766 ( .A(U_dsdc_n871), .ZN(U_dsdc_n872) );
  NOR2_X1 U_dsdc_U765 ( .A1(U_dsdc_n1244), .A2(U_dsdc_n382), .ZN(U_dsdc_n1245)
         );
  NOR2_X1 U_dsdc_U764 ( .A1(U_dsdc_n1186), .A2(U_dsdc_n363), .ZN(U_dsdc_n1187)
         );
  NAND3_X1 U_dsdc_U763 ( .A1(U_dsdc_n1434), .A2(U_dsdc_n343), .A3(U_dsdc_n1491), .ZN(U_dsdc_n926) );
  INV_X1 U_dsdc_U762 ( .A(U_dsdc_n1434), .ZN(U_dsdc_n949) );
  INV_X1 U_dsdc_U761 ( .A(U_dsdc_n1425), .ZN(U_dsdc_n857) );
  OAI21_X1 U_dsdc_U760 ( .B1(U_dsdc_n1841), .B2(U_dsdc_n304), .A(U_dsdc_n1831), 
        .ZN(U_dsdc_n1832) );
  OAI21_X1 U_dsdc_U759 ( .B1(U_dsdc_n1841), .B2(U_dsdc_n302), .A(U_dsdc_n1829), 
        .ZN(U_dsdc_n1830) );
  AOI21_X1 U_dsdc_U758 ( .B1(U_dsdc_operation_cs_2_), .B2(U_dsdc_n1506), .A(
        U_dsdc_operation_cs_3_), .ZN(U_dsdc_n1508) );
  INV_X1 U_dsdc_U757 ( .A(U_dsdc_n1454), .ZN(U_dsdc_n662) );
  INV_X1 U_dsdc_U756 ( .A(U_dsdc_n1961), .ZN(U_dsdc_n1956) );
  INV_X1 U_dsdc_U755 ( .A(U_dsdc_n1284), .ZN(U_dsdc_n1037) );
  NOR2_X1 U_dsdc_U754 ( .A1(U_dsdc_n1163), .A2(U_dsdc_rcd_cnt_0_), .ZN(
        U_dsdc_n1164) );
  XNOR2_X1 U_dsdc_U753 ( .A(U_dsdc_n1460), .B(s_cas_latency[2]), .ZN(
        U_dsdc_n1088) );
  INV_X2 U_dsdc_U752 ( .A(U_dsdc_n1464), .ZN(U_dsdc_n1461) );
  NAND2_X1 U_dsdc_U751 ( .A1(U_dsdc_n1460), .A2(s_cas_latency[2]), .ZN(
        U_dsdc_n1081) );
  INV_X2 U_dsdc_U750 ( .A(U_dsdc_n1536), .ZN(U_dsdc_n1452) );
  NAND2_X2 U_dsdc_U749 ( .A1(U_dsdc_n663), .A2(U_dsdc_n327), .ZN(U_dsdc_n1558)
         );
  AOI21_X1 U_dsdc_U748 ( .B1(U_dsdc_n699), .B2(U_dsdc_i_col_addr_4_), .A(
        U_dsdc_i_col_addr_5_), .ZN(U_dsdc_n680) );
  INV_X1 U_dsdc_U747 ( .A(U_dsdc_n1633), .ZN(U_dsdc_n1420) );
  NAND2_X2 U_dsdc_U746 ( .A1(U_dsdc_n1427), .A2(U_dsdc_access_cs_0_), .ZN(
        U_dsdc_n966) );
  NOR2_X1 U_dsdc_U745 ( .A1(U_dsdc_N4240), .A2(U_dsdc_N4239), .ZN(U_dsdc_n612)
         );
  NOR2_X1 U_dsdc_U744 ( .A1(U_dsdc_n1214), .A2(U_dsdc_n365), .ZN(U_dsdc_n1215)
         );
  AOI21_X1 U_dsdc_U743 ( .B1(U_dsdc_rcar_cnt1_2_), .B2(U_dsdc_n1585), .A(
        U_dsdc_n1584), .ZN(U_dsdc_n1586) );
  NOR2_X1 U_dsdc_U742 ( .A1(U_dsdc_n1200), .A2(U_dsdc_n364), .ZN(U_dsdc_n1201)
         );
  NAND2_X1 U_dsdc_U741 ( .A1(U_dsdc_rcar_cnt1_3_), .A2(U_dsdc_n1587), .ZN(
        U_dsdc_n1589) );
  OR3_X2 U_dsdc_U740 ( .A1(U_dsdc_row_cnt_7_), .A2(U_dsdc_row_cnt_6_), .A3(
        U_dsdc_n1770), .ZN(U_dsdc_n1765) );
  INV_X1 U_dsdc_U739 ( .A(U_dsdc_n1427), .ZN(U_dsdc_n1348) );
  INV_X1 U_dsdc_U738 ( .A(U_dsdc_n1426), .ZN(U_dsdc_n1360) );
  NAND2_X1 U_dsdc_U737 ( .A1(U_dsdc_n1425), .A2(U_dsdc_r_rw), .ZN(U_dsdc_n1628) );
  INV_X2 U_dsdc_U736 ( .A(U_dsdc_n1418), .ZN(U_dsdc_n710) );
  NAND2_X1 U_dsdc_U735 ( .A1(U_dsdc_n1434), .A2(U_dsdc_n343), .ZN(U_dsdc_n1531) );
  INV_X2 U_dsdc_U734 ( .A(U_dsdc_n1312), .ZN(U_dsdc_n1300) );
  OAI21_X1 U_dsdc_U733 ( .B1(U_dsdc_n692), .B2(U_dsdc_n667), .A(U_dsdc_n653), 
        .ZN(U_dsdc_n1357) );
  INV_X2 U_dsdc_U732 ( .A(U_dsdc_n1437), .ZN(U_dsdc_n1152) );
  NAND2_X1 U_dsdc_U731 ( .A1(U_dsdc_n904), .A2(U_dsdc_n1415), .ZN(U_dsdc_n937)
         );
  INV_X2 U_dsdc_U730 ( .A(U_dsdc_n681), .ZN(U_dsdc_n696) );
  NAND2_X1 U_dsdc_U729 ( .A1(U_dsdc_n988), .A2(U_dsdc_n940), .ZN(U_dsdc_n828)
         );
  NAND2_X1 U_dsdc_U728 ( .A1(U_dsdc_n904), .A2(U_dsdc_n1412), .ZN(U_dsdc_n674)
         );
  NOR2_X1 U_dsdc_U727 ( .A1(U_dsdc_n1362), .A2(U_dsdc_n1803), .ZN(U_dsdc_n1365) );
  OR3_X2 U_dsdc_U726 ( .A1(U_dsdc_row_cnt_9_), .A2(U_dsdc_row_cnt_8_), .A3(
        U_dsdc_n1765), .ZN(U_dsdc_n1795) );
  INV_X2 U_dsdc_U725 ( .A(U_dsdc_n904), .ZN(U_dsdc_n668) );
  NAND2_X1 U_dsdc_U724 ( .A1(U_dsdc_n867), .A2(U_dsdc_n866), .ZN(U_dsdc_n868)
         );
  INV_X1 U_dsdc_U723 ( .A(U_dsdc_n1292), .ZN(U_dsdc_n659) );
  NAND2_X1 U_dsdc_U722 ( .A1(U_dsdc_n1362), .A2(U_dsdc_n1384), .ZN(U_dsdc_n852) );
  NAND2_X1 U_dsdc_U721 ( .A1(U_dsdc_n1564), .A2(U_dsdc_n1577), .ZN(U_dsdc_n648) );
  INV_X2 U_dsdc_U720 ( .A(U_dsdc_n1432), .ZN(U_dsdc_n643) );
  OAI21_X2 U_dsdc_U719 ( .B1(U_dsdc_n1532), .B2(cr_do_self_ref_rp), .A(
        U_dsdc_n1497), .ZN(U_dsdc_n1754) );
  INV_X2 U_dsdc_U718 ( .A(U_dsdc_n1424), .ZN(U_dsdc_n684) );
  INV_X2 U_dsdc_U717 ( .A(hiu_rw), .ZN(U_dsdc_n1438) );
  INV_X2 U_dsdc_U716 ( .A(U_dsdc_n741), .ZN(U_dsdc_n736) );
  INV_X2 U_dsdc_U715 ( .A(U_dsdc_n1510), .ZN(U_dsdc_n1524) );
  INV_X2 U_dsdc_U714 ( .A(U_dsdc_n1414), .ZN(U_dsdc_n1079) );
  INV_X1 U_dsdc_U713 ( .A(U_dsdc_n1479), .ZN(U_dsdc_n1471) );
  NAND2_X1 U_dsdc_U712 ( .A1(U_dsdc_n1428), .A2(U_dsdc_n1436), .ZN(
        U_dsdc_n1469) );
  INV_X4 U_dsdc_U711 ( .A(U_dsdc_n1558), .ZN(U_dsdc_n703) );
  NAND2_X1 U_dsdc_U710 ( .A1(U_dsdc_n1414), .A2(U_cr_n58), .ZN(U_dsdc_n735) );
  INV_X2 U_dsdc_U709 ( .A(U_dsdc_n1628), .ZN(U_dsdc_n1631) );
  INV_X2 U_dsdc_U708 ( .A(U_dsdc_n1499), .ZN(U_dsdc_n1470) );
  NOR2_X1 U_dsdc_U707 ( .A1(U_dsdc_n904), .A2(U_dsdc_n165), .ZN(U_dsdc_n905)
         );
  INV_X2 U_dsdc_U706 ( .A(U_dsdc_n2053), .ZN(U_dsdc_n927) );
  INV_X2 U_dsdc_U705 ( .A(U_dsdc_n1505), .ZN(U_dsdc_n950) );
  INV_X2 U_dsdc_U704 ( .A(U_dsdc_n1195), .ZN(U_dsdc_n837) );
  INV_X2 U_dsdc_U703 ( .A(U_dsdc_n1181), .ZN(U_dsdc_n838) );
  INV_X2 U_dsdc_U702 ( .A(U_dsdc_n1237), .ZN(U_dsdc_n841) );
  INV_X2 U_dsdc_U701 ( .A(U_dsdc_n1209), .ZN(U_dsdc_n842) );
  NAND3_X1 U_dsdc_U700 ( .A1(U_dsdc_bm_bank_age_3__1_), .A2(
        U_dsdc_bm_bank_age_3__0_), .A3(U_dsdc_n1906), .ZN(U_dsdc_n1901) );
  OAI21_X1 U_dsdc_U699 ( .B1(U_dsdc_n966), .B2(U_dsdc_n466), .A(U_dsdc_n1309), 
        .ZN(U_dsdc_n968) );
  XNOR2_X1 U_dsdc_U698 ( .A(U_dsdc_n1088), .B(s_read_pipe[0]), .ZN(
        U_dsdc_add_x_2600_1_n8) );
  INV_X2 U_dsdc_U697 ( .A(U_dsdc_n1258), .ZN(U_dsdc_n751) );
  NAND2_X1 U_dsdc_U696 ( .A1(debug_ref_req), .A2(U_dsdc_n1437), .ZN(
        U_dsdc_n1447) );
  NAND2_X1 U_dsdc_U695 ( .A1(U_dsdc_bm_bank_age_0__0_), .A2(U_dsdc_n1972), 
        .ZN(U_dsdc_n1959) );
  INV_X2 U_dsdc_U694 ( .A(U_dsdc_n926), .ZN(U_dsdc_n897) );
  INV_X2 U_dsdc_U693 ( .A(U_dsdc_n903), .ZN(U_dsdc_n1061) );
  NAND2_X1 U_dsdc_U692 ( .A1(U_dsdc_n1437), .A2(U_cr_n58), .ZN(U_dsdc_n856) );
  NOR2_X1 U_dsdc_U691 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n450), .ZN(U_dsdc_n1115)
         );
  NAND2_X1 U_dsdc_U690 ( .A1(U_dsdc_n1871), .A2(U_dsdc_r_rw), .ZN(U_dsdc_n858)
         );
  INV_X2 U_dsdc_U689 ( .A(U_dsdc_n1136), .ZN(U_dsdc_n1109) );
  NAND4_X1 U_dsdc_U688 ( .A1(U_dsdc_n1574), .A2(U_dsdc_n926), .A3(U_dsdc_n1501), .A4(U_dsdc_n1510), .ZN(U_dsdc_n928) );
  NOR2_X1 U_dsdc_U687 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n454), .ZN(U_dsdc_n1132)
         );
  NOR2_X1 U_dsdc_U686 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n455), .ZN(U_dsdc_n1134)
         );
  NOR2_X1 U_dsdc_U685 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n456), .ZN(U_dsdc_n1137)
         );
  NAND2_X1 U_dsdc_U684 ( .A1(U_dsdc_n856), .A2(U_dsdc_n855), .ZN(U_dsdc_n860)
         );
  NAND2_X1 U_dsdc_U683 ( .A1(U_dsdc_n1410), .A2(U_dsdc_n1413), .ZN(
        U_dsdc_n1044) );
  NOR2_X1 U_dsdc_U682 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n451), .ZN(U_dsdc_n1116)
         );
  XNOR2_X1 U_dsdc_U681 ( .A(U_dsdc_n1092), .B(s_read_pipe[2]), .ZN(
        U_dsdc_n1091) );
  INV_X1 U_dsdc_U680 ( .A(hiu_burst_size[2]), .ZN(U_dsdc_n1263) );
  NAND2_X1 U_dsdc_U678 ( .A1(U_dsdc_n477), .A2(U_dsdc_n334), .ZN(U_dsdc_n478)
         );
  AOI21_X1 U_dsdc_U677 ( .B1(U_dsdc_n1944), .B2(U_dsdc_bm_bank_age_0__1_), .A(
        U_dsdc_bm_bank_age_0__0_), .ZN(U_dsdc_n1946) );
  NOR2_X1 U_dsdc_U676 ( .A1(U_dsdc_bm_bank_age_1__3_), .A2(U_dsdc_n1953), .ZN(
        U_dsdc_n1913) );
  NOR2_X1 U_dsdc_U674 ( .A1(U_dsdc_n1438), .A2(U_dsdc_n1284), .ZN(U_dsdc_n822)
         );
  NOR2_X1 U_dsdc_U673 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n452), .ZN(U_dsdc_n1117)
         );
  NOR2_X1 U_dsdc_U672 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n453), .ZN(U_dsdc_n1122)
         );
  OAI21_X1 U_dsdc_U671 ( .B1(U_dsdc_n304), .B2(U_dsdc_n1900), .A(U_dsdc_n302), 
        .ZN(U_dsdc_n1892) );
  NOR2_X1 U_dsdc_U670 ( .A1(U_dsdc_bm_bank_age_3__3_), .A2(U_dsdc_n1953), .ZN(
        U_dsdc_n1883) );
  OAI21_X1 U_dsdc_U669 ( .B1(U_dsdc_n1860), .B2(U_dsdc_n353), .A(U_dsdc_n178), 
        .ZN(U_dsdc_n1852) );
  INV_X1 U_dsdc_U668 ( .A(U_dsdc_n1727), .ZN(U_dsdc_n1729) );
  NAND2_X1 U_dsdc_U667 ( .A1(cr_t_xsr[8]), .A2(U_dsdc_n1754), .ZN(U_dsdc_n1726) );
  NOR2_X1 U_dsdc_U666 ( .A1(n84), .A2(U_dsdc_n1537), .ZN(U_dsdc_n1538) );
  OAI21_X1 U_dsdc_U665 ( .B1(U_dsdc_n1825), .B2(U_dsdc_n436), .A(U_dsdc_n1823), 
        .ZN(U_dsdc_n1824) );
  NAND2_X1 U_dsdc_U664 ( .A1(U_dsdc_n1496), .A2(U_dsdc_n865), .ZN(U_dsdc_n1385) );
  INV_X2 U_dsdc_U663 ( .A(U_dsdc_n1416), .ZN(U_dsdc_n2069) );
  OR4_X2 U_dsdc_U661 ( .A1(hiu_burst_size[5]), .A2(hiu_burst_size[3]), .A3(
        hiu_burst_size[2]), .A4(hiu_burst_size[1]), .ZN(U_dsdc_n1448) );
  INV_X2 U_dsdc_U660 ( .A(U_dsdc_n2058), .ZN(U_dsdc_n1511) );
  NAND3_X1 U_dsdc_U659 ( .A1(U_dsdc_n881), .A2(U_dsdc_n880), .A3(U_dsdc_n181), 
        .ZN(U_dsdc_n1065) );
  INV_X2 U_dsdc_U658 ( .A(U_dsdc_n1805), .ZN(U_dsdc_n721) );
  NAND2_X1 U_dsdc_U657 ( .A1(U_dsdc_n736), .A2(U_dsdc_n1419), .ZN(U_dsdc_n737)
         );
  AND2_X2 U_dsdc_U656 ( .A1(U_dsdc_n648), .A2(U_dsdc_n1433), .ZN(U_dsdc_n362)
         );
  INV_X1 U_dsdc_U655 ( .A(U_dsdc_n1876), .ZN(U_dsdc_n761) );
  INV_X1 U_dsdc_U654 ( .A(hiu_burst_size[0]), .ZN(U_dsdc_n1253) );
  NOR2_X1 U_dsdc_U653 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n447), .ZN(U_dsdc_n1069)
         );
  INV_X2 U_dsdc_U652 ( .A(U_dsdc_n648), .ZN(U_dsdc_n644) );
  INV_X2 U_dsdc_U651 ( .A(U_dsdc_n1315), .ZN(U_dsdc_n723) );
  INV_X2 U_dsdc_U650 ( .A(U_dsdc_n1648), .ZN(U_dsdc_n1634) );
  AOI21_X1 U_dsdc_U649 ( .B1(U_dsdc_n697), .B2(U_dsdc_i_col_addr_8_), .A(
        U_dsdc_i_col_addr_9_), .ZN(U_dsdc_n694) );
  NOR2_X1 U_dsdc_U648 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n448), .ZN(U_dsdc_n1073)
         );
  AOI21_X1 U_dsdc_U647 ( .B1(U_dsdc_n696), .B2(U_dsdc_i_col_addr_6_), .A(
        U_dsdc_i_col_addr_7_), .ZN(U_dsdc_n698) );
  INV_X2 U_dsdc_U646 ( .A(U_dsdc_n881), .ZN(U_dsdc_n675) );
  NAND2_X1 U_dsdc_U645 ( .A1(U_dsdc_n1496), .A2(U_dsdc_n1483), .ZN(
        U_dsdc_n1353) );
  INV_X2 U_dsdc_U644 ( .A(U_dsdc_n879), .ZN(U_dsdc_n682) );
  INV_X1 U_dsdc_U643 ( .A(U_dsdc_n1357), .ZN(U_dsdc_n1361) );
  NOR2_X1 U_dsdc_U642 ( .A1(U_dsdc_n1136), .A2(U_dsdc_n449), .ZN(U_dsdc_n1095)
         );
  OR3_X2 U_dsdc_U641 ( .A1(U_dsdc_row_cnt_11_), .A2(U_dsdc_row_cnt_10_), .A3(
        U_dsdc_n1795), .ZN(U_dsdc_n1794) );
  INV_X1 U_dsdc_U640 ( .A(U_dsdc_n1269), .ZN(U_dsdc_n1259) );
  NOR2_X1 U_dsdc_U639 ( .A1(U_dsdc_n934), .A2(U_dsdc_n933), .ZN(U_dsdc_n935)
         );
  INV_X2 U_dsdc_U638 ( .A(U_dsdc_n852), .ZN(U_dsdc_n1592) );
  NAND2_X1 U_dsdc_U637 ( .A1(cr_t_xsr[3]), .A2(U_dsdc_n1754), .ZN(U_dsdc_n1746) );
  INV_X2 U_dsdc_U636 ( .A(U_dsdc_n1860), .ZN(U_dsdc_n1866) );
  NAND2_X1 U_dsdc_U635 ( .A1(cr_t_xsr[0]), .A2(U_dsdc_n1754), .ZN(U_dsdc_n1755) );
  INV_X2 U_dsdc_U634 ( .A(U_dsdc_n1656), .ZN(U_dsdc_n1654) );
  NAND2_X1 U_dsdc_U633 ( .A1(cr_t_xsr[1]), .A2(U_dsdc_n1754), .ZN(U_dsdc_n1753) );
  AOI21_X1 U_dsdc_U631 ( .B1(U_dsdc_n1805), .B2(U_dsdc_n440), .A(
        U_dsdc_early_term_flag), .ZN(U_dsdc_n733) );
  AOI22_X1 U_dsdc_U630 ( .A1(U_dsdc_n1565), .A2(U_dsdc_num_init_ref_cnt_0_), 
        .B1(U_dsdc_n1667), .B2(cr_num_init_ref[0]), .ZN(U_dsdc_n1566) );
  NAND2_X1 U_dsdc_U629 ( .A1(U_dsdc_n2051), .A2(U_dsdc_n1574), .ZN(
        U_dsdc_n1575) );
  OAI211_X1 U_dsdc_U628 ( .C1(U_dsdc_num_init_ref_cnt_0_), .C2(U_dsdc_n2063), 
        .A(U_dsdc_n1433), .B(U_dsdc_num_init_ref_cnt_1_), .ZN(U_dsdc_n1569) );
  NAND2_X1 U_dsdc_U627 ( .A1(U_dsdc_n1667), .A2(cr_num_init_ref[1]), .ZN(
        U_dsdc_n1570) );
  NAND3_X1 U_dsdc_U626 ( .A1(U_dsdc_n1292), .A2(U_dsdc_n2014), .A3(
        U_dsdc_n1650), .ZN(U_dsdc_n1295) );
  NOR2_X1 U_dsdc_U625 ( .A1(U_dsdc_n988), .A2(U_dsdc_n989), .ZN(U_dsdc_n911)
         );
  NAND2_X1 U_dsdc_U624 ( .A1(U_dsdc_bm_bank_age_2__2_), .A2(U_dsdc_n1911), 
        .ZN(U_dsdc_n1837) );
  NOR2_X1 U_dsdc_U623 ( .A1(U_dsdc_n2014), .A2(U_dsdc_n1483), .ZN(U_dsdc_n1474) );
  OAI21_X1 U_dsdc_U622 ( .B1(U_dsdc_n1496), .B2(U_dsdc_n1650), .A(U_dsdc_n1342), .ZN(U_dsdc_n993) );
  NAND2_X1 U_dsdc_U621 ( .A1(U_dsdc_n1430), .A2(U_dsdc_n1728), .ZN(
        U_dsdc_n1476) );
  INV_X2 U_dsdc_U620 ( .A(U_dsdc_n1065), .ZN(U_dsdc_n1066) );
  NOR2_X1 U_dsdc_U619 ( .A1(U_dsdc_n988), .A2(U_dsdc_n1353), .ZN(U_dsdc_n836)
         );
  NAND3_X1 U_dsdc_U618 ( .A1(U_dsdc_n989), .A2(U_dsdc_r_chip_slct_0_), .A3(
        ad_sdram_type_0_), .ZN(U_dsdc_n824) );
  NAND2_X1 U_dsdc_U617 ( .A1(U_dsdc_n165), .A2(U_dsdc_n1397), .ZN(U_dsdc_n2078) );
  NAND2_X1 U_dsdc_U616 ( .A1(U_dsdc_n1423), .A2(U_dsdc_n1425), .ZN(U_dsdc_n651) );
  INV_X2 U_dsdc_U615 ( .A(U_dsdc_n702), .ZN(U_dsdc_n695) );
  NOR2_X2 U_dsdc_U614 ( .A1(U_dsdc_n1794), .A2(U_dsdc_n597), .ZN(U_dsdc_n1478)
         );
  NAND3_X1 U_dsdc_U613 ( .A1(U_dsdc_n1385), .A2(U_dsdc_n869), .A3(U_dsdc_n868), 
        .ZN(U_dsdc_n1350) );
  INV_X1 U_dsdc_U612 ( .A(U_dsdc_n989), .ZN(U_dsdc_n853) );
  INV_X2 U_dsdc_U611 ( .A(U_dsdc_n860), .ZN(U_dsdc_n916) );
  NAND2_X1 U_dsdc_U610 ( .A1(U_dsdc_n879), .A2(U_dsdc_n1060), .ZN(U_dsdc_n1313) );
  NAND3_X1 U_dsdc_U609 ( .A1(U_dsdc_n1629), .A2(U_dsdc_n1358), .A3(
        U_dsdc_n1633), .ZN(U_dsdc_n870) );
  NOR3_X1 U_dsdc_U608 ( .A1(cr_delayed_precharge), .A2(U_dsdc_n1651), .A3(
        U_dsdc_n181), .ZN(U_dsdc_wrapped_pop_flag_nxt) );
  NOR2_X1 U_dsdc_U607 ( .A1(U_dsdc_n1729), .A2(U_dsdc_n1754), .ZN(U_dsdc_n1730) );
  OAI21_X1 U_dsdc_U606 ( .B1(U_dsdc_n359), .B2(U_dsdc_n1736), .A(U_dsdc_n1733), 
        .ZN(U_dsdc_n1732) );
  NAND2_X1 U_dsdc_U605 ( .A1(U_dsdc_bm_bank_age_1__2_), .A2(U_dsdc_n1911), 
        .ZN(U_dsdc_n1915) );
  INV_X2 U_dsdc_U604 ( .A(U_dsdc_n1911), .ZN(U_dsdc_n1951) );
  INV_X2 U_dsdc_U603 ( .A(U_dsdc_n1946), .ZN(U_dsdc_n479) );
  NAND2_X1 U_dsdc_U602 ( .A1(cr_t_init[15]), .A2(U_dsdc_n1722), .ZN(
        U_dsdc_n1674) );
  INV_X2 U_dsdc_U601 ( .A(U_dsdc_n1943), .ZN(U_dsdc_n1948) );
  NAND3_X1 U_dsdc_U600 ( .A1(U_dsdc_n349), .A2(U_dsdc_n1938), .A3(
        U_dsdc_bm_bank_age_1__3_), .ZN(U_dsdc_n1939) );
  NAND2_X1 U_dsdc_U599 ( .A1(cr_t_init[9]), .A2(U_dsdc_n1722), .ZN(
        U_dsdc_n1693) );
  INV_X1 U_dsdc_U598 ( .A(U_dsdc_n1580), .ZN(U_dsdc_n1567) );
  NAND2_X1 U_dsdc_U597 ( .A1(cr_t_init[7]), .A2(U_dsdc_n1722), .ZN(
        U_dsdc_n1700) );
  NAND2_X1 U_dsdc_U596 ( .A1(cr_t_init[5]), .A2(U_dsdc_n1722), .ZN(
        U_dsdc_n1707) );
  NAND2_X1 U_dsdc_U595 ( .A1(cr_t_init[3]), .A2(U_dsdc_n1722), .ZN(
        U_dsdc_n1714) );
  OR3_X2 U_dsdc_U594 ( .A1(U_dsdc_row_cnt_13_), .A2(U_dsdc_row_cnt_12_), .A3(
        U_dsdc_n1794), .ZN(U_dsdc_n1788) );
  NOR2_X1 U_dsdc_U593 ( .A1(U_dsdc_n1666), .A2(U_dsdc_n2051), .ZN(U_dsdc_n1571) );
  INV_X2 U_dsdc_U592 ( .A(U_dsdc_n1535), .ZN(U_dsdc_n1621) );
  OAI211_X1 U_dsdc_U591 ( .C1(U_cr_n39), .C2(U_dsdc_n1532), .A(U_dsdc_n1535), 
        .B(U_dsdc_n1531), .ZN(U_dsdc_n2055) );
  OAI211_X1 U_dsdc_U590 ( .C1(U_dsdc_xsr_cnt_7_), .C2(U_dsdc_n1727), .A(
        U_dsdc_xsr_cnt_8_), .B(U_dsdc_n1733), .ZN(U_dsdc_n1725) );
  NAND2_X1 U_dsdc_U589 ( .A1(U_dsdc_bm_bank_age_3__2_), .A2(U_dsdc_n1911), 
        .ZN(U_dsdc_n1885) );
  INV_X2 U_dsdc_U585 ( .A(U_dsdc_n1788), .ZN(U_dsdc_n585) );
  INV_X1 U_dsdc_U582 ( .A(debug_ad_col_addr_0_), .ZN(U_dsdc_n1982) );
  INV_X4 U_dsdc_U581 ( .A(U_dsdc_n991), .ZN(U_dsdc_n1344) );
  OAI211_X1 U_dsdc_U580 ( .C1(U_dsdc_xsr_cnt_2_), .C2(U_dsdc_n1743), .A(
        U_dsdc_xsr_cnt_3_), .B(U_dsdc_n1750), .ZN(U_dsdc_n1745) );
  INV_X2 U_dsdc_U579 ( .A(U_dsdc_n1617), .ZN(U_dsdc_n1619) );
  NAND3_X1 U_dsdc_U578 ( .A1(U_dsdc_n1651), .A2(U_dsdc_n1313), .A3(
        U_dsdc_n1065), .ZN(U_dsdc_n895) );
  INV_X2 U_dsdc_U577 ( .A(U_dsdc_n1500), .ZN(U_dsdc_n1502) );
  AOI22_X1 U_dsdc_U576 ( .A1(U_dsdc_xsr_cnt_7_), .A2(U_dsdc_n1730), .B1(
        cr_t_xsr[7]), .B2(U_dsdc_n1754), .ZN(U_dsdc_n1731) );
  NAND3_X1 U_dsdc_U575 ( .A1(U_dsdc_n1059), .A2(U_dsdc_n1064), .A3(U_dsdc_n937), .ZN(U_dsdc_n942) );
  OAI21_X1 U_dsdc_U574 ( .B1(cr_t_xsr[6]), .B2(U_dsdc_n1733), .A(U_dsdc_n1732), 
        .ZN(U_dsdc_n1735) );
  OAI211_X1 U_dsdc_U573 ( .C1(U_dsdc_xsr_cnt_4_), .C2(U_dsdc_n1737), .A(
        U_dsdc_xsr_cnt_5_), .B(U_dsdc_n1750), .ZN(U_dsdc_n1738) );
  INV_X2 U_dsdc_U572 ( .A(U_dsdc_n1750), .ZN(U_dsdc_n1756) );
  NAND3_X1 U_dsdc_U571 ( .A1(U_dsdc_xsr_cnt_0_), .A2(U_dsdc_xsr_cnt_1_), .A3(
        U_dsdc_n1750), .ZN(U_dsdc_n1752) );
  NAND3_X1 U_dsdc_U570 ( .A1(U_dsdc_n1335), .A2(U_dsdc_rp_cnt2_2_), .A3(
        U_dsdc_n1329), .ZN(U_dsdc_n1323) );
  INV_X2 U_dsdc_U568 ( .A(U_dsdc_n760), .ZN(U_dsdc_n669) );
  INV_X2 U_dsdc_U567 ( .A(U_dsdc_n1059), .ZN(U_dsdc_n1062) );
  NOR2_X1 U_dsdc_U565 ( .A1(U_dsdc_n1350), .A2(U_dsdc_n1349), .ZN(U_dsdc_n1351) );
  OAI21_X1 U_dsdc_U564 ( .B1(U_dsdc_n873), .B2(U_dsdc_n1974), .A(
        U_dsdc_r_chip_slct_0_), .ZN(U_dsdc_n874) );
  OAI211_X1 U_dsdc_U562 ( .C1(U_dsdc_n1627), .C2(U_dsdc_n165), .A(U_dsdc_n1343), .B(U_dsdc_n1342), .ZN(U_dsdc_n1363) );
  NAND2_X1 U_dsdc_U559 ( .A1(U_dsdc_n1038), .A2(debug_ref_req), .ZN(
        U_dsdc_n939) );
  OAI21_X1 U_dsdc_U558 ( .B1(U_dsdc_n1822), .B2(U_dsdc_n437), .A(U_dsdc_n1820), 
        .ZN(U_dsdc_n1821) );
  INV_X2 U_dsdc_U557 ( .A(U_dsdc_n891), .ZN(U_dsdc_n1031) );
  INV_X1 U_dsdc_U556 ( .A(U_dsdc_n1429), .ZN(U_dsdc_n1543) );
  INV_X2 U_dsdc_U555 ( .A(U_dsdc_n2075), .ZN(U_dsdc_n2076) );
  INV_X2 U_dsdc_U554 ( .A(U_dsdc_n1758), .ZN(U_dsdc_n1579) );
  NAND2_X1 U_dsdc_U553 ( .A1(U_dsdc_n1031), .A2(U_dsdc_n181), .ZN(U_dsdc_n864)
         );
  OAI21_X1 U_dsdc_U552 ( .B1(U_dsdc_xsr_cnt_7_), .B2(U_dsdc_n1734), .A(
        U_dsdc_n1731), .ZN(U_dsdc_n393) );
  NOR2_X1 U_dsdc_U551 ( .A1(U_dsdc_n1740), .A2(U_dsdc_n1756), .ZN(U_dsdc_n1741) );
  NOR3_X1 U_dsdc_U550 ( .A1(U_dsdc_n1344), .A2(U_dsdc_n1802), .A3(U_dsdc_n1349), .ZN(U_dsdc_n938) );
  NAND3_X1 U_dsdc_U549 ( .A1(U_dsdc_bm_bank_age_2__3_), .A2(U_dsdc_n1868), 
        .A3(U_dsdc_n350), .ZN(U_dsdc_n1869) );
  AOI21_X1 U_dsdc_U548 ( .B1(U_dsdc_n902), .B2(U_dsdc_n933), .A(
        U_dsdc_i_col_addr_1_), .ZN(U_dsdc_n863) );
  INV_X2 U_dsdc_U547 ( .A(U_dsdc_n700), .ZN(U_dsdc_n677) );
  NAND2_X1 U_dsdc_U546 ( .A1(U_dsdc_n1429), .A2(cr_mode_reg_update), .ZN(
        U_dsdc_n646) );
  INV_X2 U_dsdc_U545 ( .A(U_dsdc_n2008), .ZN(U_dsdc_n1994) );
  OR3_X2 U_dsdc_U544 ( .A1(U_dsdc_n1336), .A2(cr_t_rp[1]), .A3(cr_t_rp[0]), 
        .ZN(U_dsdc_n1321) );
  AOI22_X1 U_dsdc_U543 ( .A1(U_dsdc_n1062), .A2(U_dsdc_n1061), .B1(
        U_dsdc_n1410), .B2(U_dsdc_n1060), .ZN(U_dsdc_n1063) );
  INV_X2 U_dsdc_U542 ( .A(debug_ad_row_addr[15]), .ZN(U_dsdc_n806) );
  OAI211_X1 U_dsdc_U541 ( .C1(U_dsdc_n1316), .C2(U_dsdc_n1315), .A(
        U_dsdc_n1314), .B(U_dsdc_n1313), .ZN(U_dsdc_n1317) );
  NOR2_X2 U_dsdc_U540 ( .A1(U_dsdc_n573), .A2(U_dsdc_n2063), .ZN(U_dsdc_n1791)
         );
  NAND2_X2 U_dsdc_U539 ( .A1(U_dsdc_n1403), .A2(U_dsdc_n1063), .ZN(
        U_dsdc_n1268) );
  AND2_X2 U_dsdc_U537 ( .A1(U_dsdc_n861), .A2(U_dsdc_r_chip_slct_0_), .ZN(
        U_dsdc_n862) );
  OAI211_X1 U_dsdc_U536 ( .C1(U_dsdc_n1361), .C2(U_dsdc_n1360), .A(
        U_dsdc_n1359), .B(U_dsdc_n1358), .ZN(U_dsdc_n1366) );
  AND2_X2 U_dsdc_U535 ( .A1(U_dsdc_n2013), .A2(U_dsdc_n1409), .ZN(U_dsdc_n1977) );
  INV_X1 U_dsdc_U534 ( .A(debug_ad_col_addr_14_), .ZN(U_dsdc_n1141) );
  OAI21_X1 U_dsdc_U533 ( .B1(U_dsdc_n2079), .B2(U_dsdc_n2076), .A(
        U_dsdc_early_term_flag), .ZN(U_dsdc_n2077) );
  INV_X2 U_dsdc_U532 ( .A(U_dsdc_n1409), .ZN(U_dsdc_n1056) );
  OAI21_X1 U_dsdc_U531 ( .B1(U_dsdc_n1372), .B2(debug_ref_req), .A(
        U_dsdc_n1038), .ZN(U_dsdc_n957) );
  INV_X2 U_dsdc_U530 ( .A(U_dsdc_n1812), .ZN(U_dsdc_n1118) );
  NAND2_X1 U_dsdc_U529 ( .A1(U_dsdc_n864), .A2(U_dsdc_n1412), .ZN(U_dsdc_n992)
         );
  OAI21_X1 U_dsdc_U527 ( .B1(U_dsdc_n940), .B2(U_dsdc_n939), .A(U_dsdc_n938), 
        .ZN(U_dsdc_n941) );
  OR2_X2 U_dsdc_U526 ( .A1(U_dsdc_n1612), .A2(U_dsdc_n1601), .ZN(U_dsdc_n1495)
         );
  NAND2_X1 U_dsdc_U525 ( .A1(U_dsdc_n1791), .A2(U_dsdc_row_cnt_12_), .ZN(
        U_dsdc_n576) );
  NOR3_X1 U_dsdc_U524 ( .A1(U_dsdc_n1507), .A2(U_dsdc_access_cs_4_), .A3(
        U_dsdc_n1348), .ZN(U_dsdc_n1356) );
  NAND2_X1 U_dsdc_U523 ( .A1(U_dsdc_n1791), .A2(U_dsdc_row_cnt_6_), .ZN(
        U_dsdc_n583) );
  NAND2_X1 U_dsdc_U522 ( .A1(U_dsdc_n1671), .A2(cr_exn_mode_value[8]), .ZN(
        U_dsdc_n1074) );
  AOI21_X1 U_dsdc_U521 ( .B1(U_dsdc_n354), .B2(U_dsdc_n942), .A(U_dsdc_n941), 
        .ZN(U_dsdc_n943) );
  NAND2_X1 U_dsdc_U520 ( .A1(U_dsdc_n1791), .A2(U_dsdc_row_cnt_10_), .ZN(
        U_dsdc_n590) );
  INV_X2 U_dsdc_U519 ( .A(ad_data_mask[0]), .ZN(U_dsdc_n2015) );
  INV_X1 U_dsdc_U518 ( .A(U_dsdc_n1875), .ZN(U_dsdc_n1874) );
  NAND2_X1 U_dsdc_U517 ( .A1(U_dsdc_n1791), .A2(U_dsdc_row_cnt_4_), .ZN(
        U_dsdc_n591) );
  AOI22_X1 U_dsdc_U516 ( .A1(U_dsdc_n1268), .A2(U_dsdc_cas_cnt_2_), .B1(
        U_dsdc_n1269), .B2(U_dsdc_r_burst_size_2_), .ZN(U_dsdc_n1262) );
  INV_X2 U_dsdc_U515 ( .A(U_dsdc_n932), .ZN(U_dsdc_n948) );
  NAND2_X1 U_dsdc_U514 ( .A1(U_dsdc_n1791), .A2(U_dsdc_row_cnt_14_), .ZN(
        U_dsdc_n578) );
  INV_X2 U_dsdc_U512 ( .A(U_dsdc_n1670), .ZN(U_dsdc_n1108) );
  NAND2_X1 U_dsdc_U511 ( .A1(U_dsdc_n1791), .A2(U_dsdc_row_cnt_2_), .ZN(
        U_dsdc_n577) );
  NAND2_X1 U_dsdc_U510 ( .A1(U_dsdc_n1671), .A2(cr_exn_mode_value[4]), .ZN(
        U_dsdc_n1107) );
  OR2_X2 U_dsdc_U509 ( .A1(U_dsdc_n1581), .A2(U_dsdc_n1495), .ZN(U_dsdc_N430)
         );
  INV_X2 U_dsdc_U508 ( .A(U_dsdc_n992), .ZN(U_dsdc_n767) );
  NOR2_X1 U_dsdc_U507 ( .A1(U_dsdc_n1679), .A2(U_dsdc_n1722), .ZN(U_dsdc_n1680) );
  NAND2_X1 U_dsdc_U506 ( .A1(U_dsdc_n1627), .A2(U_dsdc_n1626), .ZN(
        U_dsdc_s_rd_end_nxt) );
  AOI22_X1 U_dsdc_U505 ( .A1(U_dsdc_n1671), .A2(cr_exn_mode_value[11]), .B1(
        U_dsdc_r_col_addr_10_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1070) );
  OR2_X2 U_dsdc_U503 ( .A1(U_dsdc_n1603), .A2(U_dsdc_n1596), .ZN(U_dsdc_n1608)
         );
  NAND2_X1 U_dsdc_U502 ( .A1(U_dsdc_n1791), .A2(U_dsdc_row_cnt_8_), .ZN(
        U_dsdc_n592) );
  NAND2_X1 U_dsdc_U501 ( .A1(U_dsdc_n1671), .A2(cr_exn_mode_value[5]), .ZN(
        U_dsdc_n1101) );
  NAND2_X1 U_dsdc_U500 ( .A1(U_dsdc_n1671), .A2(cr_exn_mode_value[6]), .ZN(
        U_dsdc_n1096) );
  INV_X2 U_dsdc_U498 ( .A(U_dsdc_n588), .ZN(U_dsdc_n1783) );
  INV_X1 U_dsdc_U497 ( .A(debug_ad_row_addr[6]), .ZN(U_dsdc_n1098) );
  INV_X2 U_dsdc_U496 ( .A(U_dsdc_n584), .ZN(U_dsdc_n594) );
  NAND2_X1 U_dsdc_U495 ( .A1(U_dsdc_n1417), .A2(U_dsdc_n1650), .ZN(
        U_dsdc_n1318) );
  INV_X2 U_dsdc_U494 ( .A(ad_data_mask[2]), .ZN(U_dsdc_n2017) );
  INV_X1 U_dsdc_U493 ( .A(debug_ad_row_addr[4]), .ZN(U_dsdc_n1111) );
  INV_X2 U_dsdc_U492 ( .A(ad_data_mask[1]), .ZN(U_dsdc_n2016) );
  INV_X2 U_dsdc_U491 ( .A(U_dsdc_n587), .ZN(U_dsdc_n595) );
  NAND4_X1 U_dsdc_U490 ( .A1(U_dsdc_n1436), .A2(U_dsdc_n1428), .A3(
        U_dsdc_n1038), .A4(U_dsdc_n1449), .ZN(U_dsdc_n921) );
  OAI22_X1 U_dsdc_U489 ( .A1(U_dsdc_n1260), .A2(U_dsdc_n327), .B1(U_dsdc_n1259), .B2(U_dsdc_n182), .ZN(U_dsdc_n1261) );
  INV_X2 U_dsdc_U488 ( .A(debug_ad_row_addr[13]), .ZN(U_dsdc_n800) );
  NAND4_X1 U_dsdc_U487 ( .A1(U_dsdc_n1978), .A2(U_dsdc_n944), .A3(U_dsdc_n943), 
        .A4(U_dsdc_n992), .ZN(U_dsdc_n947) );
  OAI211_X1 U_dsdc_U486 ( .C1(U_dsdc_init_cnt_12_), .C2(U_dsdc_n1686), .A(
        U_dsdc_init_cnt_13_), .B(U_dsdc_n1676), .ZN(U_dsdc_n1678) );
  INV_X2 U_dsdc_U485 ( .A(U_dsdc_n582), .ZN(U_dsdc_n1771) );
  AOI21_X1 U_dsdc_U484 ( .B1(cr_t_rcar[0]), .B2(U_dsdc_n1602), .A(U_dsdc_n1601), .ZN(U_dsdc_n1600) );
  OR3_X2 U_dsdc_U483 ( .A1(U_dsdc_init_cnt_15_), .A2(U_dsdc_init_cnt_14_), 
        .A3(U_dsdc_n482), .ZN(U_dsdc_n1675) );
  INV_X1 U_dsdc_U482 ( .A(debug_ad_row_addr[10]), .ZN(U_dsdc_n1028) );
  OAI211_X1 U_dsdc_U481 ( .C1(U_dsdc_n875), .C2(U_dsdc_n934), .A(U_dsdc_n922), 
        .B(U_dsdc_n874), .ZN(U_dsdc_n876) );
  INV_X2 U_dsdc_U480 ( .A(U_dsdc_n586), .ZN(U_dsdc_n593) );
  INV_X1 U_dsdc_U479 ( .A(debug_ad_row_addr[8]), .ZN(U_dsdc_n1076) );
  OAI22_X1 U_dsdc_U478 ( .A1(U_dsdc_n1590), .A2(U_cr_n72), .B1(U_dsdc_n1589), 
        .B2(U_dsdc_n1588), .ZN(U_dsdc_rcar_cnt1_nxt[3]) );
  INV_X2 U_dsdc_U477 ( .A(U_dsdc_n1610), .ZN(U_dsdc_n1611) );
  INV_X4 U_dsdc_U476 ( .A(debug_ad_bank_addr[0]), .ZN(U_dsdc_n1127) );
  OAI22_X1 U_dsdc_U475 ( .A1(U_dsdc_n1590), .A2(U_cr_n104), .B1(U_dsdc_n1586), 
        .B2(U_dsdc_n1588), .ZN(U_dsdc_rcar_cnt1_nxt[2]) );
  NAND4_X1 U_dsdc_U474 ( .A1(U_dsdc_n922), .A2(U_dsdc_n921), .A3(U_dsdc_n920), 
        .A4(U_dsdc_n958), .ZN(U_dsdc_n923) );
  INV_X2 U_dsdc_U473 ( .A(U_dsdc_oldest_bank_1_), .ZN(U_dsdc_n1000) );
  XNOR2_X1 U_dsdc_U472 ( .A(U_dsdc_n618), .B(U_dsdc_n358), .ZN(
        U_dsdc_num_row[9]) );
  INV_X1 U_dsdc_U471 ( .A(U_dsdc_n1849), .ZN(U_dsdc_n1847) );
  OAI21_X1 U_dsdc_U470 ( .B1(U_dsdc_rcar_cnt2_0_), .B2(U_dsdc_n1597), .A(
        U_dsdc_n1594), .ZN(U_dsdc_rcar_cnt2_nxt[0]) );
  INV_X1 U_dsdc_U469 ( .A(U_dsdc_n1890), .ZN(U_dsdc_n1888) );
  OAI22_X1 U_dsdc_U468 ( .A1(U_dsdc_n1590), .A2(U_cr_n151), .B1(U_dsdc_n1582), 
        .B2(U_dsdc_n1588), .ZN(U_dsdc_rcar_cnt1_nxt[1]) );
  INV_X2 U_dsdc_U467 ( .A(U_dsdc_n1542), .ZN(U_dsdc_n1545) );
  INV_X2 U_dsdc_U466 ( .A(ad_data_mask[3]), .ZN(U_dsdc_n2019) );
  INV_X1 U_dsdc_U465 ( .A(U_dsdc_n1920), .ZN(U_dsdc_n1918) );
  AOI21_X1 U_dsdc_U464 ( .B1(U_dsdc_n1867), .B2(U_dsdc_n1849), .A(U_dsdc_n1850), .ZN(U_dsdc_n1848) );
  INV_X2 U_dsdc_U463 ( .A(U_dsdc_n1138), .ZN(U_dsdc_n605) );
  AOI22_X1 U_dsdc_U462 ( .A1(U_dsdc_n1138), .A2(U_dsdc_n1408), .B1(
        U_dsdc_r_col_addr_12_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1133) );
  INV_X2 U_dsdc_U461 ( .A(U_dsdc_n1990), .ZN(U_dsdc_n1139) );
  AOI22_X1 U_dsdc_U460 ( .A1(U_dsdc_n1138), .A2(U_dsdc_n1407), .B1(
        U_dsdc_r_col_addr_13_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1135) );
  OAI21_X1 U_dsdc_U459 ( .B1(U_dsdc_n1546), .B2(U_dsdc_n1263), .A(U_dsdc_n750), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_I5_2_) );
  NAND3_X1 U_dsdc_U458 ( .A1(U_dsdc_n853), .A2(U_dsdc_n1038), .A3(U_dsdc_n1473), .ZN(U_dsdc_n854) );
  OAI21_X1 U_dsdc_U457 ( .B1(U_dsdc_n1546), .B2(U_dmc_n16), .A(U_dsdc_n748), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_I5_4_) );
  NOR2_X1 U_dsdc_U456 ( .A1(U_dsdc_n1694), .A2(U_dsdc_n1724), .ZN(U_dsdc_n1695) );
  NAND4_X1 U_dsdc_U455 ( .A1(U_dsdc_n605), .A2(U_dsdc_n184), .A3(U_dsdc_n1409), 
        .A4(U_dsdc_n1136), .ZN(U_dsdc_n1128) );
  NOR2_X1 U_dsdc_U454 ( .A1(U_dsdc_n1701), .A2(U_dsdc_n1724), .ZN(U_dsdc_n1702) );
  NOR2_X1 U_dsdc_U453 ( .A1(U_dsdc_n1708), .A2(U_dsdc_n1724), .ZN(U_dsdc_n1709) );
  NOR2_X1 U_dsdc_U452 ( .A1(U_dsdc_n1687), .A2(U_dsdc_n1724), .ZN(U_dsdc_n1688) );
  OAI211_X2 U_dsdc_U451 ( .C1(U_dsdc_n1545), .C2(U_dsdc_n432), .A(U_dsdc_n1544), .B(U_dsdc_n1543), .ZN(U_dsdc_n2093) );
  OAI211_X1 U_dsdc_U450 ( .C1(U_dsdc_n1724), .C2(U_dsdc_n482), .A(U_dsdc_n1678), .B(U_dsdc_n1677), .ZN(U_dsdc_n416) );
  OAI21_X1 U_dsdc_U449 ( .B1(U_dsdc_n1721), .B2(U_dsdc_n1724), .A(U_dsdc_n1720), .ZN(U_dsdc_n404) );
  OAI21_X1 U_dsdc_U448 ( .B1(U_dsdc_init_cnt_0_), .B2(U_dsdc_n1724), .A(
        U_dsdc_n1723), .ZN(U_dsdc_n403) );
  AOI22_X1 U_dsdc_U446 ( .A1(debug_ad_col_addr_11_), .A2(U_dsdc_n1815), .B1(
        U_dsdc_r_col_addr_11_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1814) );
  AOI22_X1 U_dsdc_U445 ( .A1(debug_ad_col_addr_10_), .A2(U_dsdc_n1815), .B1(
        U_dsdc_r_col_addr_10_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1816) );
  INV_X2 U_dsdc_U444 ( .A(U_dsdc_n1902), .ZN(U_dsdc_n1897) );
  INV_X2 U_dsdc_U443 ( .A(U_dsdc_n1396), .ZN(U_dsdc_n2012) );
  INV_X2 U_dsdc_U442 ( .A(U_dsdc_n753), .ZN(U_dsdc_n754) );
  OAI21_X1 U_dsdc_U441 ( .B1(U_dsdc_init_cnt_0_), .B2(U_dsdc_init_cnt_1_), .A(
        U_dsdc_n1715), .ZN(U_dsdc_n1718) );
  INV_X2 U_dsdc_U440 ( .A(U_dsdc_n2083), .ZN(U_dsdc_n2084) );
  OAI211_X1 U_dsdc_U439 ( .C1(U_dsdc_init_cnt_4_), .C2(U_dsdc_n1704), .A(
        U_dsdc_init_cnt_5_), .B(U_dsdc_n1715), .ZN(U_dsdc_n1706) );
  XNOR2_X1 U_dsdc_U438 ( .A(U_dsdc_n607), .B(U_dsdc_n357), .ZN(
        U_dsdc_num_row[11]) );
  INV_X2 U_dsdc_U437 ( .A(U_dsdc_n1862), .ZN(U_dsdc_n1857) );
  OAI211_X1 U_dsdc_U436 ( .C1(U_dsdc_init_cnt_6_), .C2(U_dsdc_n1697), .A(
        U_dsdc_init_cnt_7_), .B(U_dsdc_n1715), .ZN(U_dsdc_n1699) );
  OR2_X2 U_dsdc_U435 ( .A1(U_dsdc_n1965), .A2(U_dsdc_n1962), .ZN(U_dsdc_n1957)
         );
  NAND2_X1 U_dsdc_U434 ( .A1(U_dsdc_n1687), .A2(U_dsdc_n1715), .ZN(
        U_dsdc_n1691) );
  OAI211_X1 U_dsdc_U432 ( .C1(U_dsdc_init_cnt_8_), .C2(U_dsdc_n1690), .A(
        U_dsdc_init_cnt_9_), .B(U_dsdc_n1715), .ZN(U_dsdc_n1692) );
  AOI22_X1 U_dsdc_U431 ( .A1(debug_ad_col_addr_14_), .A2(U_dsdc_n1815), .B1(
        U_dsdc_r_col_addr_14_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1549) );
  OAI211_X1 U_dsdc_U430 ( .C1(U_dsdc_init_cnt_10_), .C2(U_dsdc_n1683), .A(
        U_dsdc_init_cnt_11_), .B(U_dsdc_n1715), .ZN(U_dsdc_n1685) );
  INV_X2 U_dsdc_U429 ( .A(U_dsdc_n1932), .ZN(U_dsdc_n1927) );
  NAND2_X1 U_dsdc_U428 ( .A1(U_dsdc_n1679), .A2(U_dsdc_n1715), .ZN(
        U_dsdc_n1682) );
  AOI22_X1 U_dsdc_U427 ( .A1(debug_ad_col_addr_2_), .A2(U_dsdc_n1815), .B1(
        U_dsdc_r_col_addr_2_), .B2(U_dsdc_n619), .ZN(U_dsdc_n1811) );
  INV_X2 U_dsdc_U426 ( .A(U_dsdc_n749), .ZN(U_dsdc_DP_OP_1642_126_2028_I5_3_)
         );
  INV_X2 U_dsdc_U425 ( .A(U_dsdc_n1865), .ZN(U_dsdc_n1864) );
  INV_X2 U_dsdc_U424 ( .A(U_dsdc_n1968), .ZN(U_dsdc_n1963) );
  NOR3_X1 U_dsdc_U423 ( .A1(hiu_terminate), .A2(U_dsdc_dqs_mask_end), .A3(
        U_dsdc_n475), .ZN(U_dsdc_n973) );
  INV_X2 U_dsdc_U422 ( .A(U_dsdc_n747), .ZN(U_dsdc_DP_OP_1642_126_2028_I5_5_)
         );
  OAI21_X1 U_dsdc_U421 ( .B1(U_dsdc_n2041), .B2(U_dsdc_n1990), .A(U_dsdc_n1549), .ZN(U_dsdc_i_col_addr_nxt[14]) );
  INV_X2 U_dsdc_U420 ( .A(U_dsdc_n1905), .ZN(U_dsdc_n1904) );
  OAI21_X1 U_dsdc_U419 ( .B1(U_dsdc_n2041), .B2(U_dsdc_n1993), .A(U_dsdc_n1811), .ZN(U_dsdc_n320) );
  OAI21_X1 U_dsdc_U418 ( .B1(U_dsdc_n2041), .B2(U_dsdc_n1986), .A(U_dsdc_n1814), .ZN(U_dsdc_n317) );
  OAI21_X1 U_dsdc_U417 ( .B1(U_dsdc_n2041), .B2(U_dsdc_n1984), .A(U_dsdc_n1816), .ZN(U_dsdc_n316) );
  INV_X2 U_dsdc_U416 ( .A(U_dsdc_n1935), .ZN(U_dsdc_n1934) );
  OAI21_X1 U_dsdc_U415 ( .B1(U_dsdc_init_cnt_12_), .B2(U_dsdc_n1682), .A(
        U_dsdc_n1681), .ZN(U_dsdc_n415) );
  OAI211_X1 U_dsdc_U414 ( .C1(U_dsdc_n1430), .C2(U_dsdc_n1505), .A(
        U_dsdc_n2060), .B(U_dsdc_n1504), .ZN(U_dsdc_n1516) );
  OAI21_X1 U_dsdc_U413 ( .B1(U_dsdc_init_cnt_6_), .B2(U_dsdc_n1705), .A(
        U_dsdc_n1703), .ZN(U_dsdc_n409) );
  OAI211_X1 U_dsdc_U412 ( .C1(U_dsdc_n1724), .C2(U_dsdc_n1686), .A(
        U_dsdc_n1685), .B(U_dsdc_n1684), .ZN(U_dsdc_n414) );
  INV_X2 U_dsdc_U411 ( .A(U_dsdc_n2067), .ZN(U_dsdc_n720) );
  OAI21_X1 U_dsdc_U410 ( .B1(U_dsdc_init_cnt_10_), .B2(U_dsdc_n1691), .A(
        U_dsdc_n1689), .ZN(U_dsdc_n413) );
  OAI21_X1 U_dsdc_U409 ( .B1(U_dsdc_init_cnt_8_), .B2(U_dsdc_n1698), .A(
        U_dsdc_n1696), .ZN(U_dsdc_n411) );
  OR2_X2 U_dsdc_U408 ( .A1(U_dsdc_n973), .A2(s_rd_start), .ZN(U_dsdc_n217) );
  AOI22_X1 U_dsdc_U407 ( .A1(U_dsdc_n2049), .A2(U_dsdc_r_burst_size_5_), .B1(
        hiu_burst_size[5]), .B2(U_dsdc_n2048), .ZN(U_dsdc_n2047) );
  AOI22_X1 U_dsdc_U406 ( .A1(U_dsdc_n2049), .A2(U_dsdc_r_burst_size_1_), .B1(
        hiu_burst_size[1]), .B2(U_dsdc_n2048), .ZN(U_dsdc_n2043) );
  AOI22_X1 U_dsdc_U405 ( .A1(U_dsdc_n2049), .A2(U_dsdc_r_burst_size_3_), .B1(
        hiu_burst_size[3]), .B2(U_dsdc_n2048), .ZN(U_dsdc_n2045) );
  AOI22_X1 U_dsdc_U404 ( .A1(U_dsdc_n2049), .A2(U_dsdc_r_burst_size_0_), .B1(
        hiu_burst_size[0]), .B2(U_dsdc_n2048), .ZN(U_dsdc_n2042) );
  AOI22_X1 U_dsdc_U403 ( .A1(U_dsdc_n2049), .A2(U_dsdc_r_burst_size_4_), .B1(
        hiu_burst_size[4]), .B2(U_dsdc_n2048), .ZN(U_dsdc_n2046) );
  INV_X4 U_dsdc_U402 ( .A(U_dsdc_n987), .ZN(U_dsdc_n978) );
  AOI22_X1 U_dsdc_U401 ( .A1(U_dsdc_n2049), .A2(U_dsdc_r_wrapped_burst), .B1(
        hiu_wrapped_burst), .B2(U_dsdc_n2048), .ZN(U_dsdc_n2050) );
  INV_X2 U_dsdc_U400 ( .A(U_dsdc_n1971), .ZN(U_dsdc_n1970) );
  AOI22_X1 U_dsdc_U399 ( .A1(U_dsdc_n2049), .A2(U_dsdc_r_burst_size_2_), .B1(
        hiu_burst_size[2]), .B2(U_dsdc_n2048), .ZN(U_dsdc_n2044) );
  AND2_X2 U_dsdc_U397 ( .A1(U_dsdc_bm_row_addr_1__10_), .A2(U_dsdc_n604), .ZN(
        U_dsdc_n176) );
  INV_X2 U_dsdc_U396 ( .A(U_dsdc_n1270), .ZN(U_dsdc_n1266) );
  OAI211_X1 U_dsdc_U395 ( .C1(U_dsdc_n1354), .C2(U_dsdc_n1353), .A(
        U_dsdc_n1352), .B(U_dsdc_n1351), .ZN(U_dsdc_n1355) );
  INV_X2 U_dsdc_U394 ( .A(U_dsdc_n1395), .ZN(U_dsdc_n2068) );
  OAI211_X1 U_dsdc_U393 ( .C1(U_dsdc_n989), .C2(U_dsdc_n1354), .A(U_dsdc_n919), 
        .B(U_dsdc_n918), .ZN(U_dsdc_n924) );
  INV_X2 U_dsdc_U392 ( .A(U_dsdc_n1339), .ZN(U_dsdc_n1341) );
  NAND2_X1 U_dsdc_U391 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__7_), .ZN(
        U_dsdc_n797) );
  OAI211_X1 U_dsdc_U390 ( .C1(U_dsdc_n1541), .C2(U_dsdc_n341), .A(U_dsdc_n1540), .B(U_dsdc_n1539), .ZN(U_dsdc_n2095) );
  INV_X2 U_dsdc_U389 ( .A(U_dsdc_n2046), .ZN(U_dsdc_n275) );
  INV_X2 U_dsdc_U388 ( .A(U_dsdc_n2047), .ZN(U_dsdc_n276) );
  INV_X2 U_dsdc_U387 ( .A(U_dsdc_n2050), .ZN(U_dsdc_n277) );
  NAND2_X1 U_dsdc_U386 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__13_), 
        .ZN(U_dsdc_n778) );
  OAI21_X1 U_dsdc_U385 ( .B1(U_dsdc_bm_rc_cnt_3__2_), .B2(
        U_dsdc_bm_rc_cnt_3__3_), .A(U_dsdc_n978), .ZN(U_dsdc_n831) );
  INV_X2 U_dsdc_U384 ( .A(U_dsdc_n2045), .ZN(U_dsdc_n274) );
  INV_X2 U_dsdc_U383 ( .A(U_dsdc_n2044), .ZN(U_dsdc_n273) );
  AOI22_X1 U_dsdc_U382 ( .A1(U_dsdc_n2007), .A2(U_dsdc_r_col_addr_1_), .B1(
        debug_ad_col_addr_1_), .B2(U_dsdc_n2048), .ZN(U_dsdc_n1991) );
  INV_X2 U_dsdc_U381 ( .A(U_dsdc_n2043), .ZN(U_dsdc_n272) );
  OAI21_X1 U_dsdc_U379 ( .B1(U_dsdc_n2068), .B2(U_dsdc_n1483), .A(
        U_dsdc_r_chip_slct_0_), .ZN(U_dsdc_n1346) );
  INV_X2 U_dsdc_U378 ( .A(U_dsdc_n2042), .ZN(U_dsdc_n271) );
  AOI22_X1 U_dsdc_U377 ( .A1(U_dsdc_r_col_addr_14_), .A2(U_dsdc_n2007), .B1(
        debug_ad_col_addr_14_), .B2(U_dsdc_n2048), .ZN(U_dsdc_n1989) );
  INV_X2 U_dsdc_U376 ( .A(U_dsdc_n2022), .ZN(U_dsdc_n254) );
  INV_X2 U_dsdc_U375 ( .A(U_dsdc_n2021), .ZN(U_dsdc_n253) );
  INV_X2 U_dsdc_U374 ( .A(U_dsdc_n1991), .ZN(U_dsdc_n240) );
  INV_X1 U_dsdc_U373 ( .A(U_dsdc_n1283), .ZN(U_dsdc_n1288) );
  OAI21_X1 U_dsdc_U372 ( .B1(debug_ad_col_addr_12_), .B2(U_dsdc_n2010), .A(
        U_dsdc_n1987), .ZN(U_dsdc_n236) );
  AND4_X2 U_dsdc_U371 ( .A1(U_dsdc_n832), .A2(U_dsdc_n831), .A3(U_dsdc_n830), 
        .A4(U_dsdc_n829), .ZN(U_dsdc_n835) );
  INV_X2 U_dsdc_U370 ( .A(U_dsdc_n808), .ZN(U_dsdc_n809) );
  AND2_X2 U_dsdc_U369 ( .A1(U_dsdc_n785), .A2(U_dsdc_n800), .ZN(U_dsdc_n333)
         );
  OR3_X2 U_dsdc_U368 ( .A1(U_dsdc_n602), .A2(U_dsdc_n816), .A3(
        U_dsdc_bm_row_addr_0__7_), .ZN(U_dsdc_n332) );
  AND2_X2 U_dsdc_U367 ( .A1(U_dsdc_n813), .A2(debug_ad_row_addr[1]), .ZN(
        U_dsdc_n318) );
  NAND2_X1 U_dsdc_U366 ( .A1(U_dsdc_n1394), .A2(U_dsdc_bm_bank_status_1_), 
        .ZN(U_dsdc_n997) );
  NAND2_X1 U_dsdc_U365 ( .A1(U_dsdc_n1394), .A2(U_dsdc_bm_bank_status_3_), 
        .ZN(U_dsdc_n996) );
  NAND2_X1 U_dsdc_U364 ( .A1(U_dsdc_n1394), .A2(U_dsdc_bm_bank_status_0_), 
        .ZN(U_dsdc_n1002) );
  NAND2_X1 U_dsdc_U363 ( .A1(U_dsdc_n1394), .A2(U_dsdc_bm_bank_status_2_), 
        .ZN(U_dsdc_n1392) );
  INV_X2 U_dsdc_U362 ( .A(U_dsdc_n1394), .ZN(U_dsdc_n1322) );
  AND2_X2 U_dsdc_U361 ( .A1(U_dsdc_n533), .A2(U_dsdc_n425), .ZN(U_dsdc_n177)
         );
  INV_X2 U_dsdc_U360 ( .A(U_dsdc_n818), .ZN(U_dsdc_n817) );
  NAND3_X1 U_dsdc_U359 ( .A1(U_dsdc_n986), .A2(U_dsdc_n984), .A3(U_dsdc_n982), 
        .ZN(U_dsdc_n847) );
  NAND3_X1 U_dsdc_U358 ( .A1(U_dsdc_n984), .A2(U_dsdc_n983), .A3(U_dsdc_n982), 
        .ZN(U_dsdc_n985) );
  NAND2_X1 U_dsdc_U357 ( .A1(U_dsdc_n975), .A2(U_dsdc_n828), .ZN(U_dsdc_n910)
         );
  NAND3_X1 U_dsdc_U356 ( .A1(U_dsdc_n1003), .A2(U_dsdc_n1000), .A3(U_dsdc_n999), .ZN(U_dsdc_n1001) );
  NAND2_X2 U_dsdc_U355 ( .A1(U_dsdc_n1345), .A2(U_dsdc_n977), .ZN(U_dsdc_n1112) );
  NAND2_X2 U_dsdc_U354 ( .A1(U_dsdc_n1112), .A2(U_dsdc_n1136), .ZN(
        U_dsdc_n1166) );
  INV_X1 U_dsdc_U353 ( .A(U_dsdc_n1146), .ZN(U_dsdc_n1030) );
  INV_X2 U_dsdc_U352 ( .A(U_dsdc_n1166), .ZN(U_dsdc_n1159) );
  INV_X2 U_dsdc_U351 ( .A(U_dsdc_n1020), .ZN(U_dsdc_n1012) );
  NOR3_X1 U_dsdc_U350 ( .A1(U_dsdc_n1020), .A2(U_dsdc_n179), .A3(U_dsdc_n338), 
        .ZN(U_dsdc_n1021) );
  OAI21_X1 U_dsdc_U349 ( .B1(U_dsdc_bm_close_bank_2_), .B2(U_dsdc_n1392), .A(
        U_dsdc_n310), .ZN(U_dsdc_N4449) );
  OAI21_X1 U_dsdc_U347 ( .B1(U_dsdc_bm_close_bank_3_), .B2(U_dsdc_n996), .A(
        U_dsdc_n313), .ZN(U_dsdc_N4496) );
  INV_X2 U_dsdc_U346 ( .A(U_dsdc_n960), .ZN(U_dsdc_n894) );
  INV_X2 U_dsdc_U345 ( .A(U_dsdc_n1017), .ZN(U_dsdc_n1013) );
  INV_X2 U_dsdc_U344 ( .A(U_dsdc_n972), .ZN(U_dsdc_n946) );
  INV_X1 U_dsdc_U343 ( .A(U_dsdc_n1328), .ZN(U_dsdc_n1327) );
  INV_X2 U_dsdc_U342 ( .A(U_dsdc_n963), .ZN(U_dsdc_n961) );
  NAND2_X2 U_dsdc_U341 ( .A1(U_dsdc_n1320), .A2(U_dsdc_n1057), .ZN(
        U_dsdc_n1121) );
  NAND3_X1 U_dsdc_U340 ( .A1(U_dsdc_n1389), .A2(U_dsdc_n1320), .A3(
        U_dsdc_n1319), .ZN(U_dsdc_n[2089]) );
  INV_X1 U_dsdc_U339 ( .A(U_dsdc_n1039), .ZN(U_dsdc_n962) );
  OR3_X2 U_dsdc_U338 ( .A1(hiu_terminate), .A2(U_dsdc_n1374), .A3(U_dsdc_n963), 
        .ZN(U_dsdc_N429) );
  INV_X1 U_dsdc_U337 ( .A(U_dsdc_n1374), .ZN(U_dsdc_n1376) );
  INV_X2 U_dsdc_U336 ( .A(U_dsdc_n1051), .ZN(U_dsdc_n1052) );
  OR2_X2 U_dsdc_U335 ( .A1(U_dsdc_bm_num_open_bank_4_), .A2(U_dsdc_n1026), 
        .ZN(U_dsdc_n603) );
  OAI21_X1 U_dsdc_U334 ( .B1(U_dsdc_n1131), .B2(U_dsdc_n1127), .A(U_dsdc_n1126), .ZN(U_dsdc_N422) );
  NAND2_X2 U_dsdc_U331 ( .A1(U_dsdc_n173), .A2(U_dsdc_n355), .ZN(U_dsdc_n649)
         );
  NOR2_X1 U_dsdc_U330 ( .A1(U_dsdc_init_cnt_0_), .A2(U_dsdc_init_cnt_1_), .ZN(
        U_dsdc_n1719) );
  XNOR2_X1 U_dsdc_U328 ( .A(U_dsdc_n194), .B(U_dsdc_wtr_cnt_0_), .ZN(
        U_dsdc_n1246) );
  NOR2_X1 U_dsdc_U327 ( .A1(U_dsdc_rcar_cnt1_1_), .A2(U_dsdc_rcar_cnt1_0_), 
        .ZN(U_dsdc_n1583) );
  NAND2_X2 U_dsdc_U326 ( .A1(U_dsdc_n355), .A2(U_dsdc_access_cs_0_), .ZN(
        U_dsdc_n690) );
  INV_X2 U_dsdc_U325 ( .A(U_dsdc_N4239), .ZN(U_dsdc_n598) );
  INV_X2 U_dsdc_U324 ( .A(U_dsdc_n1708), .ZN(U_dsdc_n1704) );
  NOR2_X1 U_dsdc_U323 ( .A1(U_dsdc_n1536), .A2(U_dsdc_n1581), .ZN(U_dsdc_n2053) );
  INV_X2 U_dsdc_U322 ( .A(U_dsdc_n1234), .ZN(U_dsdc_n1227) );
  INV_X2 U_dsdc_U321 ( .A(U_dsdc_n1193), .ZN(U_dsdc_n1188) );
  INV_X2 U_dsdc_U320 ( .A(U_dsdc_n1207), .ZN(U_dsdc_n1202) );
  INV_X2 U_dsdc_U319 ( .A(U_dsdc_n1179), .ZN(U_dsdc_n1174) );
  NAND2_X1 U_dsdc_U318 ( .A1(U_dsdc_n1458), .A2(U_dsdc_n657), .ZN(U_dsdc_n1292) );
  NAND2_X1 U_dsdc_U317 ( .A1(U_dsdc_n1434), .A2(U_dsdc_n1435), .ZN(
        U_dsdc_n1505) );
  INV_X2 U_dsdc_U316 ( .A(U_dsdc_n1650), .ZN(U_dsdc_n865) );
  NAND2_X1 U_dsdc_U315 ( .A1(U_dsdc_n360), .A2(U_dsdc_n1426), .ZN(U_dsdc_n1343) );
  NOR2_X1 U_dsdc_U314 ( .A1(U_dsdc_n1422), .A2(U_dsdc_n1803), .ZN(U_dsdc_n1591) );
  INV_X2 U_dsdc_U313 ( .A(U_dsdc_n1701), .ZN(U_dsdc_n1697) );
  INV_X2 U_dsdc_U312 ( .A(U_dsdc_n1526), .ZN(U_dsdc_n2065) );
  OAI21_X1 U_dsdc_U311 ( .B1(U_dsdc_n352), .B2(U_dsdc_n1930), .A(U_dsdc_n335), 
        .ZN(U_dsdc_n1922) );
  INV_X2 U_dsdc_U310 ( .A(U_dsdc_n933), .ZN(U_dsdc_n1060) );
  INV_X2 U_dsdc_U309 ( .A(U_dsdc_n945), .ZN(U_dsdc_n869) );
  INV_X2 U_dsdc_U308 ( .A(U_dsdc_n1754), .ZN(U_dsdc_n1733) );
  INV_X2 U_dsdc_U307 ( .A(U_dsdc_add_x_2600_1_n8), .ZN(U_dsdc_n1089) );
  INV_X2 U_dsdc_U306 ( .A(U_dsdc_n856), .ZN(U_dsdc_n994) );
  NAND3_X1 U_dsdc_U305 ( .A1(U_dsdc_n1866), .A2(U_dsdc_bm_bank_age_2__1_), 
        .A3(U_dsdc_bm_bank_age_2__0_), .ZN(U_dsdc_n1861) );
  NAND2_X1 U_dsdc_U304 ( .A1(cr_t_init[11]), .A2(U_dsdc_n1722), .ZN(
        U_dsdc_n1684) );
  NAND2_X1 U_dsdc_U303 ( .A1(cr_t_init[13]), .A2(U_dsdc_n1722), .ZN(
        U_dsdc_n1677) );
  NAND2_X1 U_dsdc_U302 ( .A1(U_dsdc_n1556), .A2(U_dsdc_n758), .ZN(U_dsdc_n672)
         );
  INV_X2 U_dsdc_U301 ( .A(U_dsdc_n982), .ZN(U_dsdc_n826) );
  NAND2_X1 U_dsdc_U300 ( .A1(U_dsdc_bm_bank_age_3__3_), .A2(U_dsdc_n1908), 
        .ZN(U_dsdc_n1909) );
  INV_X4 U_dsdc_U299 ( .A(U_dsdc_n1629), .ZN(U_dsdc_n685) );
  INV_X2 U_dsdc_U298 ( .A(U_dsdc_n1694), .ZN(U_dsdc_n1690) );
  NAND2_X1 U_dsdc_U297 ( .A1(U_dsdc_n1740), .A2(U_dsdc_n1750), .ZN(
        U_dsdc_n1744) );
  INV_X2 U_dsdc_U296 ( .A(U_dsdc_n1456), .ZN(U_dsdc_n1457) );
  INV_X2 U_dsdc_U295 ( .A(U_dsdc_n1687), .ZN(U_dsdc_n1683) );
  INV_X2 U_dsdc_U294 ( .A(U_dsdc_DP_OP_1642_126_2028_I4), .ZN(U_dsdc_n755) );
  NAND4_X1 U_dsdc_U293 ( .A1(U_dsdc_n902), .A2(U_dsdc_n903), .A3(U_dsdc_n904), 
        .A4(U_dsdc_n181), .ZN(U_dsdc_n861) );
  OAI21_X1 U_dsdc_U292 ( .B1(U_dsdc_n933), .B2(U_dsdc_n903), .A(U_dsdc_n902), 
        .ZN(U_dsdc_n906) );
  OAI21_X1 U_dsdc_U291 ( .B1(U_dsdc_xsr_cnt_0_), .B2(U_dsdc_n1756), .A(
        U_dsdc_n1755), .ZN(U_dsdc_n386) );
  OAI211_X1 U_dsdc_U290 ( .C1(U_dsdc_n1492), .C2(U_dsdc_n2063), .A(
        U_dsdc_n1540), .B(U_dsdc_n1488), .ZN(U_dsdc_auto_ref_en_nxt) );
  INV_X1 U_dsdc_U289 ( .A(U_dsdc_n1525), .ZN(U_dsdc_n1529) );
  OAI21_X1 U_dsdc_U288 ( .B1(U_dsdc_n906), .B2(U_dsdc_n905), .A(U_dsdc_n1412), 
        .ZN(U_dsdc_n920) );
  NOR2_X1 U_dsdc_U286 ( .A1(debug_ref_req), .A2(sdram_req_i), .ZN(U_dsdc_n1449) );
  INV_X4 U_dsdc_U285 ( .A(U_dsdc_n764), .ZN(U_dsdc_n1382) );
  NAND2_X1 U_dsdc_U283 ( .A1(U_dsdc_n1791), .A2(U_dsdc_n575), .ZN(U_dsdc_n589)
         );
  NAND2_X1 U_dsdc_U282 ( .A1(U_dsdc_n1791), .A2(U_dsdc_n580), .ZN(U_dsdc_n584)
         );
  INV_X1 U_dsdc_U280 ( .A(U_dsdc_n589), .ZN(U_dsdc_n1796) );
  AND2_X2 U_dsdc_U279 ( .A1(U_dsdc_n921), .A2(U_dsdc_n852), .ZN(U_dsdc_n1352)
         );
  NAND2_X1 U_dsdc_U278 ( .A1(U_dsdc_n1694), .A2(U_dsdc_n1715), .ZN(
        U_dsdc_n1698) );
  OAI21_X1 U_dsdc_U277 ( .B1(debug_ad_col_addr_12_), .B2(U_dsdc_n1819), .A(
        U_dsdc_n1547), .ZN(U_dsdc_i_col_addr_nxt[12]) );
  OAI21_X1 U_dsdc_U276 ( .B1(U_dsdc_init_cnt_4_), .B2(U_dsdc_n1712), .A(
        U_dsdc_n1710), .ZN(U_dsdc_n407) );
  NAND2_X1 U_dsdc_U275 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__13_), 
        .ZN(U_dsdc_n776) );
  NAND2_X1 U_dsdc_U273 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__7_), .ZN(
        U_dsdc_n795) );
  NAND2_X1 U_dsdc_U272 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__9_), .ZN(
        U_dsdc_n786) );
  INV_X4 U_dsdc_U271 ( .A(U_dsdc_n599), .ZN(U_dsdc_n159) );
  NAND2_X1 U_dsdc_U270 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__12_), 
        .ZN(U_dsdc_n516) );
  OAI21_X1 U_dsdc_U269 ( .B1(U_dsdc_bm_rc_cnt_2__2_), .B2(
        U_dsdc_bm_rc_cnt_2__3_), .A(U_dsdc_n159), .ZN(U_dsdc_n832) );
  NAND2_X1 U_dsdc_U268 ( .A1(U_dsdc_n159), .A2(U_dsdc_bm_row_addr_2__13_), 
        .ZN(U_dsdc_n777) );
  NAND2_X1 U_dsdc_U267 ( .A1(U_dsdc_n978), .A2(U_dsdc_bm_row_addr_3__9_), .ZN(
        U_dsdc_n788) );
  NAND2_X1 U_dsdc_U266 ( .A1(U_dsdc_n159), .A2(U_dsdc_bm_row_addr_2__7_), .ZN(
        U_dsdc_n796) );
  OAI21_X1 U_dsdc_U264 ( .B1(U_dsdc_bm_rc_cnt_1__2_), .B2(
        U_dsdc_bm_rc_cnt_1__3_), .A(U_dsdc_n604), .ZN(U_dsdc_n830) );
  INV_X2 U_dsdc_U263 ( .A(U_dsdc_n1782), .ZN(U_dsdc_n372) );
  NAND2_X4 U_dsdc_U261 ( .A1(U_dsdc_n1166), .A2(U_dsdc_n978), .ZN(U_dsdc_n313)
         );
  NOR3_X1 U_dsdc_U260 ( .A1(U_dsdc_n1020), .A2(U_dsdc_bm_num_open_bank_3_), 
        .A3(U_dsdc_n338), .ZN(U_dsdc_n1018) );
  OAI22_X1 U_dsdc_U259 ( .A1(U_dsdc_n1243), .A2(U_dsdc_n1241), .B1(U_dsdc_n313), .B2(U_cr_n120), .ZN(U_dsdc_N4461) );
  OAI22_X1 U_dsdc_U258 ( .A1(U_dsdc_n1243), .A2(U_dsdc_bm_ras_cnt_3__0_), .B1(
        U_dsdc_n313), .B2(n95), .ZN(U_dsdc_N4460) );
  NOR2_X2 U_dsdc_U257 ( .A1(U_dsdc_n887), .A2(U_dsdc_n817), .ZN(U_dsdc_n981)
         );
  NOR3_X1 U_dsdc_U256 ( .A1(U_dsdc_n1310), .A2(cr_delayed_precharge), .A3(
        U_dsdc_n1309), .ZN(U_dsdc_n1311) );
  NOR2_X1 U_dsdc_U255 ( .A1(U_dsdc_n1310), .A2(U_cr_n58), .ZN(U_dsdc_n1035) );
  OAI21_X1 U_dsdc_U254 ( .B1(U_dsdc_bm_close_bank_0_), .B2(U_dsdc_n1002), .A(
        n83), .ZN(U_dsdc_N4355) );
  NOR3_X1 U_dsdc_U253 ( .A1(U_dsdc_n1286), .A2(U_dsdc_n1285), .A3(U_dsdc_n1557), .ZN(U_dsdc_n1287) );
  OAI21_X1 U_dsdc_U252 ( .B1(U_dsdc_bm_close_bank_1_), .B2(U_dsdc_n997), .A(
        U_dsdc_n620), .ZN(U_dsdc_N4402) );
  OAI21_X2 U_dsdc_U251 ( .B1(U_dsdc_n1006), .B2(U_dsdc_n340), .A(U_dsdc_n1005), 
        .ZN(U_dsdc_n293) );
  NAND2_X4 U_dsdc_U250 ( .A1(U_dsdc_n1166), .A2(U_dsdc_n159), .ZN(U_dsdc_n310)
         );
  AOI22_X1 U_dsdc_U249 ( .A1(U_dsdc_n1092), .A2(s_read_pipe[2]), .B1(
        U_dsdc_n1093), .B2(U_dsdc_n158), .ZN(U_dsdc_n554) );
  INV_X1 U_dsdc_U248 ( .A(U_dsdc_n1091), .ZN(U_dsdc_n158) );
  XOR2_X1 U_dsdc_U247 ( .A(U_dsdc_n1085), .B(U_dsdc_n1084), .Z(
        U_dsdc_cas_latency_1_) );
  NAND2_X1 U_dsdc_U246 ( .A1(U_dsdc_n1393), .A2(U_dsdc_n157), .ZN(
        U_dsdc_n[2091]) );
  AOI211_X1 U_dsdc_U245 ( .C1(U_dsdc_access_cs_1_), .C2(U_dsdc_n154), .A(
        U_dsdc_n1388), .B(U_dsdc_n156), .ZN(U_dsdc_n157) );
  OAI211_X1 U_dsdc_U244 ( .C1(cr_delayed_precharge), .C2(U_dsdc_n155), .A(
        U_dsdc_n1387), .B(U_dsdc_n1389), .ZN(U_dsdc_n156) );
  INV_X1 U_dsdc_U243 ( .A(U_dsdc_n1386), .ZN(U_dsdc_n155) );
  NAND3_X1 U_dsdc_U242 ( .A1(U_dsdc_n2069), .A2(U_dsdc_n1385), .A3(U_dsdc_n153), .ZN(U_dsdc_n154) );
  NOR2_X1 U_dsdc_U241 ( .A1(U_dsdc_n1384), .A2(U_dsdc_n1383), .ZN(U_dsdc_n153)
         );
  OAI21_X1 U_dsdc_U240 ( .B1(U_dsdc_n462), .B2(U_dsdc_n151), .A(U_dsdc_n152), 
        .ZN(U_dsdc_n366) );
  AOI21_X1 U_dsdc_U239 ( .B1(U_dsdc_n1791), .B2(U_dsdc_n462), .A(U_dsdc_n1797), 
        .ZN(U_dsdc_n152) );
  INV_X1 U_dsdc_U238 ( .A(U_dsdc_n1800), .ZN(U_dsdc_n151) );
  OAI211_X1 U_dsdc_U237 ( .C1(U_dsdc_init_cnt_14_), .C2(U_dsdc_n148), .A(
        U_dsdc_n149), .B(U_dsdc_n150), .ZN(U_dsdc_n417) );
  NAND2_X1 U_dsdc_U236 ( .A1(U_dsdc_n1722), .A2(cr_t_init[14]), .ZN(
        U_dsdc_n150) );
  NAND3_X1 U_dsdc_U235 ( .A1(U_dsdc_n1676), .A2(U_dsdc_init_cnt_14_), .A3(
        U_dsdc_n482), .ZN(U_dsdc_n149) );
  NAND2_X1 U_dsdc_U234 ( .A1(U_dsdc_n1715), .A2(U_dsdc_n147), .ZN(U_dsdc_n148)
         );
  INV_X1 U_dsdc_U233 ( .A(U_dsdc_n482), .ZN(U_dsdc_n147) );
  AOI22_X1 U_dsdc_U232 ( .A1(U_dsdc_n313), .A2(U_dsdc_n145), .B1(U_cr_n128), 
        .B2(U_dsdc_n144), .ZN(U_dsdc_N4462) );
  AOI22_X1 U_dsdc_U230 ( .A1(U_dsdc_bm_ras_cnt_3__2_), .A2(U_dsdc_n1238), .B1(
        U_dsdc_bm_ras_cnt_3__3_), .B2(U_dsdc_n1244), .ZN(U_dsdc_n145) );
  AOI22_X1 U_dsdc_U229 ( .A1(U_dsdc_n313), .A2(U_dsdc_n143), .B1(n96), .B2(
        U_dsdc_n144), .ZN(U_dsdc_N4475) );
  INV_X1 U_dsdc_U228 ( .A(U_dsdc_n313), .ZN(U_dsdc_n144) );
  AOI22_X1 U_dsdc_U227 ( .A1(U_dsdc_bm_rc_cnt_3__2_), .A2(U_dsdc_n1228), .B1(
        U_dsdc_bm_rc_cnt_3__3_), .B2(U_dsdc_n1234), .ZN(U_dsdc_n143) );
  OAI211_X1 U_dsdc_U226 ( .C1(U_dsdc_n1382), .C2(U_dsdc_n139), .A(U_dsdc_n140), 
        .B(U_dsdc_n142), .ZN(U_dsdc_n288) );
  OAI211_X1 U_dsdc_U225 ( .C1(U_dsdc_DP_OP_1642_126_2028_n15), .C2(
        U_dsdc_DP_OP_1642_126_2028_n7), .A(U_dsdc_n1380), .B(U_dsdc_n141), 
        .ZN(U_dsdc_n142) );
  NAND2_X1 U_dsdc_U224 ( .A1(U_dsdc_DP_OP_1642_126_2028_n15), .A2(
        U_dsdc_DP_OP_1642_126_2028_n7), .ZN(U_dsdc_n141) );
  NAND2_X1 U_dsdc_U223 ( .A1(U_dsdc_n1381), .A2(U_dsdc_N1764), .ZN(U_dsdc_n140) );
  AOI21_X1 U_dsdc_U222 ( .B1(U_dsdc_n1823), .B2(U_dsdc_data_cnt_2_), .A(
        U_dsdc_n1822), .ZN(U_dsdc_n139) );
  OAI21_X1 U_dsdc_U221 ( .B1(U_dsdc_n1473), .B2(debug_ref_req), .A(
        U_dsdc_n1038), .ZN(U_dsdc_n1354) );
  NOR4_X1 U_dsdc_U219 ( .A1(U_dsdc_n1581), .A2(U_dsdc_n1667), .A3(U_dsdc_n1580), .A4(U_dsdc_n137), .ZN(U_dsdc_n1590) );
  NAND3_X1 U_dsdc_U218 ( .A1(U_dsdc_n1579), .A2(U_dsdc_n1578), .A3(U_dsdc_n92), 
        .ZN(U_dsdc_n137) );
  OR3_X1 U_dsdc_U216 ( .A1(U_dsdc_N4241), .A2(U_dsdc_N4240), .A3(U_dsdc_N4239), 
        .ZN(U_dsdc_n613) );
  OAI21_X1 U_dsdc_U214 ( .B1(U_dsdc_n701), .B2(U_dsdc_i_col_addr_11_), .A(
        U_dsdc_n700), .ZN(U_dsdc_n1986) );
  OAI21_X1 U_dsdc_U213 ( .B1(cr_num_open_banks[4]), .B2(U_dsdc_n385), .A(
        U_dsdc_n134), .ZN(U_dsdc_n982) );
  OAI221_X1 U_dsdc_U212 ( .B1(U_dsdc_n131), .B2(U_dsdc_bm_num_open_bank_3_), 
        .C1(U_dsdc_n131), .C2(n92), .A(U_dsdc_n133), .ZN(U_dsdc_n134) );
  AOI22_X1 U_dsdc_U211 ( .A1(cr_num_open_banks[4]), .A2(U_dsdc_n385), .B1(
        cr_num_open_banks[3]), .B2(U_dsdc_n179), .ZN(U_dsdc_n133) );
  AOI21_X1 U_dsdc_U209 ( .B1(U_dsdc_n338), .B2(cr_num_open_banks[2]), .A(
        U_dsdc_n130), .ZN(U_dsdc_n131) );
  NOR2_X1 U_dsdc_U208 ( .A1(U_dsdc_n128), .A2(U_dsdc_n129), .ZN(U_dsdc_n130)
         );
  AOI22_X1 U_dsdc_U207 ( .A1(cr_num_open_banks[1]), .A2(U_dsdc_n180), .B1(
        U_dsdc_n340), .B2(cr_num_open_banks[0]), .ZN(U_dsdc_n129) );
  OAI22_X1 U_dsdc_U206 ( .A1(cr_num_open_banks[2]), .A2(U_dsdc_n338), .B1(
        cr_num_open_banks[1]), .B2(U_dsdc_n180), .ZN(U_dsdc_n128) );
  NAND3_X1 U_dsdc_U204 ( .A1(U_dsdc_n125), .A2(U_dsdc_n493), .A3(U_dsdc_n126), 
        .ZN(U_dsdc_n496) );
  AOI22_X1 U_dsdc_U203 ( .A1(U_dsdc_n816), .A2(U_dsdc_bm_row_addr_0__7_), .B1(
        U_dsdc_n801), .B2(U_dsdc_bm_row_addr_0__3_), .ZN(U_dsdc_n126) );
  AOI21_X1 U_dsdc_U202 ( .B1(U_dsdc_bm_row_addr_0__9_), .B2(U_dsdc_n803), .A(
        U_dsdc_n572), .ZN(U_dsdc_n125) );
  OAI211_X1 U_dsdc_U201 ( .C1(U_dsdc_n1382), .C2(U_dsdc_n120), .A(U_dsdc_n121), 
        .B(U_dsdc_n124), .ZN(U_dsdc_n286) );
  OAI221_X1 U_dsdc_U200 ( .B1(U_dsdc_DP_OP_1642_126_2028_n28), .B2(U_dsdc_n25), 
        .C1(U_dsdc_n123), .C2(U_dsdc_DP_OP_1642_126_2028_n11), .A(U_dsdc_n1380), .ZN(U_dsdc_n124) );
  INV_X1 U_dsdc_U199 ( .A(U_dsdc_DP_OP_1642_126_2028_n28), .ZN(U_dsdc_n123) );
  NAND2_X1 U_dsdc_U197 ( .A1(U_dsdc_N1762), .A2(U_dsdc_n1381), .ZN(U_dsdc_n121) );
  AOI21_X1 U_dsdc_U196 ( .B1(U_dsdc_data_cnt_0_), .B2(U_dsdc_n1444), .A(
        U_dsdc_n1825), .ZN(U_dsdc_n120) );
  OAI21_X1 U_dsdc_U195 ( .B1(U_dsdc_n116), .B2(U_dsdc_n118), .A(U_dsdc_n119), 
        .ZN(U_dsdc_n278) );
  OAI21_X1 U_dsdc_U194 ( .B1(U_dsdc_n116), .B2(U_dsdc_n113), .A(s_cke), .ZN(
        U_dsdc_n119) );
  NOR2_X1 U_dsdc_U193 ( .A1(U_dsdc_n2061), .A2(U_dsdc_n117), .ZN(U_dsdc_n118)
         );
  INV_X1 U_dsdc_U192 ( .A(U_dsdc_n2060), .ZN(U_dsdc_n117) );
  OR3_X1 U_dsdc_U191 ( .A1(U_dsdc_n2055), .A2(U_dsdc_n114), .A3(U_dsdc_n115), 
        .ZN(U_dsdc_n116) );
  OAI211_X1 U_dsdc_U190 ( .C1(U_dsdc_n2056), .C2(U_dsdc_n2057), .A(
        U_dsdc_n2058), .B(U_dsdc_n2059), .ZN(U_dsdc_n115) );
  NAND4_X1 U_dsdc_U189 ( .A1(U_dsdc_n2051), .A2(U_dsdc_n2052), .A3(
        U_dsdc_n2053), .A4(U_dsdc_n2054), .ZN(U_dsdc_n114) );
  OAI211_X1 U_dsdc_U188 ( .C1(U_dsdc_n2066), .C2(U_dsdc_n111), .A(U_dsdc_n2065), .B(U_dsdc_n112), .ZN(U_dsdc_n113) );
  NAND2_X1 U_dsdc_U187 ( .A1(U_dsdc_n2063), .A2(U_dsdc_n2064), .ZN(U_dsdc_n112) );
  INV_X1 U_dsdc_U186 ( .A(U_dsdc_n2062), .ZN(U_dsdc_n111) );
  AOI22_X1 U_dsdc_U185 ( .A1(U_dsdc_n310), .A2(U_dsdc_n109), .B1(U_cr_n128), 
        .B2(U_dsdc_n108), .ZN(U_dsdc_N4415) );
  AOI22_X1 U_dsdc_U183 ( .A1(U_dsdc_bm_ras_cnt_2__2_), .A2(U_dsdc_n1210), .B1(
        U_dsdc_bm_ras_cnt_2__3_), .B2(U_dsdc_n1214), .ZN(U_dsdc_n109) );
  AOI22_X1 U_dsdc_U182 ( .A1(U_dsdc_n310), .A2(U_dsdc_n107), .B1(n96), .B2(
        U_dsdc_n108), .ZN(U_dsdc_N4428) );
  INV_X1 U_dsdc_U181 ( .A(U_dsdc_n310), .ZN(U_dsdc_n108) );
  AOI22_X1 U_dsdc_U180 ( .A1(U_dsdc_bm_rc_cnt_2__2_), .A2(U_dsdc_n1203), .B1(
        U_dsdc_bm_rc_cnt_2__3_), .B2(U_dsdc_n1207), .ZN(U_dsdc_n107) );
  OAI21_X1 U_dsdc_U179 ( .B1(U_dsdc_n1166), .B2(U_dsdc_n105), .A(U_dsdc_n106), 
        .ZN(U_dsdc_N4141) );
  NAND2_X1 U_dsdc_U178 ( .A1(cr_t_rcd[2]), .A2(U_dsdc_n1166), .ZN(U_dsdc_n106)
         );
  NAND2_X1 U_dsdc_U177 ( .A1(U_dsdc_n1165), .A2(U_dsdc_rcd_cnt_2_), .ZN(
        U_dsdc_n105) );
  NAND3_X1 U_dsdc_U176 ( .A1(U_dsdc_n1173), .A2(U_dsdc_n103), .A3(U_dsdc_n104), 
        .ZN(U_dsdc_N420) );
  AOI22_X1 U_dsdc_U175 ( .A1(U_dsdc_n1121), .A2(debug_ad_col_addr_0_), .B1(
        U_dsdc_N1685), .B2(U_dsdc_n1138), .ZN(U_dsdc_n104) );
  AOI22_X1 U_dsdc_U174 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_0_), .B1(
        cr_exn_mode_value[0]), .B2(U_dsdc_n102), .ZN(U_dsdc_n103) );
  INV_X1 U_dsdc_U173 ( .A(U_dsdc_n1513), .ZN(U_dsdc_n102) );
  OAI21_X1 U_dsdc_U172 ( .B1(U_dsdc_n554), .B2(U_dsdc_n1393), .A(U_dsdc_n101), 
        .ZN(U_dsdc_N4129) );
  NAND3_X1 U_dsdc_U171 ( .A1(U_dsdc_n1393), .A2(U_dsdc_n1094), .A3(
        U_dsdc_cas_latency_cnt_3_), .ZN(U_dsdc_n101) );
  AOI22_X1 U_dsdc_U170 ( .A1(U_dsdc_n99), .A2(U_dsdc_n434), .B1(U_dsdc_n98), 
        .B2(U_dsdc_n100), .ZN(U_dsdc_n231) );
  NOR2_X1 U_dsdc_U169 ( .A1(U_dsdc_n434), .A2(U_dsdc_n1971), .ZN(U_dsdc_n100)
         );
  NAND2_X1 U_dsdc_U168 ( .A1(U_dsdc_bm_bank_age_0__3_), .A2(U_dsdc_n1973), 
        .ZN(U_dsdc_n99) );
  AOI22_X1 U_dsdc_U167 ( .A1(U_dsdc_bm_bank_age_0__3_), .A2(U_dsdc_n2081), 
        .B1(U_dsdc_n1972), .B2(U_dsdc_n458), .ZN(U_dsdc_n98) );
  AOI21_X1 U_dsdc_U166 ( .B1(U_dsdc_n97), .B2(U_dsdc_n1375), .A(U_dsdc_n909), 
        .ZN(U_dsdc_N402) );
  NOR4_X1 U_dsdc_U165 ( .A1(U_dsdc_n1373), .A2(U_dsdc_n908), .A3(U_dsdc_n94), 
        .A4(U_dsdc_n96), .ZN(U_dsdc_n97) );
  OAI211_X1 U_dsdc_U164 ( .C1(U_dsdc_n994), .C2(U_dsdc_n95), .A(U_dsdc_n922), 
        .B(U_dsdc_n901), .ZN(U_dsdc_n96) );
  INV_X1 U_dsdc_U163 ( .A(U_dsdc_n917), .ZN(U_dsdc_n95) );
  NAND3_X1 U_dsdc_U162 ( .A1(U_dsdc_n920), .A2(U_dsdc_n1309), .A3(U_dsdc_n93), 
        .ZN(U_dsdc_n94) );
  NOR2_X1 U_dsdc_U161 ( .A1(U_dsdc_n907), .A2(U_dsdc_n1974), .ZN(U_dsdc_n93)
         );
  NOR3_X1 U_dsdc_U160 ( .A1(U_dsdc_row_cnt_1_), .A2(U_dsdc_row_cnt_0_), .A3(
        U_dsdc_n92), .ZN(U_dsdc_n325) );
  INV_X1 U_dsdc_U159 ( .A(U_dsdc_n1791), .ZN(U_dsdc_n92) );
  INV_X1 U_dsdc_U158 ( .A(U_dsdc_n91), .ZN(U_dsdc_n1984) );
  AOI21_X1 U_dsdc_U157 ( .B1(U_dsdc_n702), .B2(U_dsdc_n444), .A(U_dsdc_n701), 
        .ZN(U_dsdc_n91) );
  XNOR2_X1 U_dsdc_U156 ( .A(U_dsdc_n90), .B(hiu_burst_size[5]), .ZN(
        U_dsdc_N1767) );
  AOI22_X1 U_dsdc_U155 ( .A1(hiu_burst_size[4]), .A2(U_dsdc_N1991), .B1(
        U_dsdc_DP_OP_1642_126_2028_n42), .B2(U_dsdc_DP_OP_1642_126_2028_n34), 
        .ZN(U_dsdc_n90) );
  AOI21_X1 U_dsdc_U154 ( .B1(U_dsdc_n798), .B2(U_dsdc_n801), .A(U_dsdc_n89), 
        .ZN(U_dsdc_n514) );
  NOR3_X1 U_dsdc_U153 ( .A1(U_dsdc_n800), .A2(U_dsdc_n785), .A3(
        U_dsdc_bm_row_addr_0__13_), .ZN(U_dsdc_n89) );
  AOI21_X2 U_dsdc_U152 ( .B1(U_dsdc_bm_row_addr_2__14_), .B2(U_dsdc_n159), .A(
        U_dsdc_n88), .ZN(U_dsdc_n548) );
  NAND2_X2 U_dsdc_U151 ( .A1(U_dsdc_n547), .A2(U_dsdc_n87), .ZN(U_dsdc_n88) );
  AOI22_X2 U_dsdc_U150 ( .A1(U_dsdc_n998), .A2(U_dsdc_bm_row_addr_0__14_), 
        .B1(U_dsdc_n604), .B2(U_dsdc_bm_row_addr_1__14_), .ZN(U_dsdc_n87) );
  AND2_X4 U_dsdc_U149 ( .A1(U_dsdc_n799), .A2(U_dsdc_n86), .ZN(U_dsdc_n813) );
  AOI22_X1 U_dsdc_U148 ( .A1(U_dsdc_bm_row_addr_3__1_), .A2(U_dsdc_n978), .B1(
        U_dsdc_bm_row_addr_1__1_), .B2(U_dsdc_n604), .ZN(U_dsdc_n86) );
  AOI221_X1 U_dsdc_U147 ( .B1(U_dsdc_n1339), .B2(U_dsdc_n1282), .C1(
        U_dsdc_n1281), .C2(U_dsdc_n1282), .A(U_dsdc_n1340), .ZN(
        U_dsdc_cas_cnt_nxt[1]) );
  AOI22_X1 U_dsdc_U146 ( .A1(U_dsdc_n620), .A2(U_dsdc_n84), .B1(U_cr_n128), 
        .B2(U_dsdc_n621), .ZN(U_dsdc_N4368) );
  AOI22_X1 U_dsdc_U144 ( .A1(U_dsdc_bm_ras_cnt_1__2_), .A2(U_dsdc_n1196), .B1(
        U_dsdc_bm_ras_cnt_1__3_), .B2(U_dsdc_n1200), .ZN(U_dsdc_n84) );
  AOI22_X1 U_dsdc_U143 ( .A1(U_dsdc_n620), .A2(U_dsdc_n82), .B1(n96), .B2(
        U_dsdc_n621), .ZN(U_dsdc_N4381) );
  AOI22_X1 U_dsdc_U141 ( .A1(U_dsdc_bm_rc_cnt_1__2_), .A2(U_dsdc_n1189), .B1(
        U_dsdc_bm_rc_cnt_1__3_), .B2(U_dsdc_n1193), .ZN(U_dsdc_n82) );
  OAI21_X1 U_dsdc_U140 ( .B1(U_dsdc_n1166), .B2(U_dsdc_n80), .A(U_dsdc_n81), 
        .ZN(U_dsdc_N4284) );
  NAND2_X1 U_dsdc_U139 ( .A1(cr_t_ras_min[3]), .A2(U_dsdc_n1166), .ZN(
        U_dsdc_n81) );
  NAND2_X1 U_dsdc_U138 ( .A1(U_dsdc_n1161), .A2(U_dsdc_bm_ras_cnt_max_3_), 
        .ZN(U_dsdc_n80) );
  NAND3_X1 U_dsdc_U137 ( .A1(U_dsdc_n1171), .A2(U_dsdc_n78), .A3(U_dsdc_n79), 
        .ZN(U_dsdc_N418) );
  AOI22_X1 U_dsdc_U136 ( .A1(U_dsdc_n1121), .A2(debug_ad_col_addr_2_), .B1(
        U_dsdc_n1810), .B2(U_dsdc_n1138), .ZN(U_dsdc_n79) );
  AOI22_X1 U_dsdc_U135 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_2_), .B1(
        cr_exn_mode_value[2]), .B2(U_dsdc_n1671), .ZN(U_dsdc_n78) );
  OAI211_X1 U_dsdc_U131 ( .C1(U_dsdc_n1382), .C2(U_dsdc_n72), .A(U_dsdc_n73), 
        .B(U_dsdc_n75), .ZN(U_dsdc_n290) );
  OAI211_X1 U_dsdc_U130 ( .C1(U_dsdc_DP_OP_1642_126_2028_n3), .C2(
        U_dsdc_DP_OP_1642_126_2028_n13), .A(U_dsdc_n1380), .B(U_dsdc_n74), 
        .ZN(U_dsdc_n75) );
  NAND2_X1 U_dsdc_U129 ( .A1(U_dsdc_DP_OP_1642_126_2028_n3), .A2(
        U_dsdc_DP_OP_1642_126_2028_n13), .ZN(U_dsdc_n74) );
  NAND2_X1 U_dsdc_U128 ( .A1(U_dsdc_n1381), .A2(U_dsdc_N1766), .ZN(U_dsdc_n73)
         );
  AOI21_X1 U_dsdc_U127 ( .B1(U_dsdc_data_cnt_4_), .B2(U_dsdc_n1820), .A(
        U_dsdc_n762), .ZN(U_dsdc_n72) );
  NOR2_X1 U_dsdc_U126 ( .A1(U_dsdc_n71), .A2(U_dsdc_n945), .ZN(U_dsdc_n972) );
  AOI211_X1 U_dsdc_U125 ( .C1(U_dsdc_n1041), .C2(U_dsdc_n1428), .A(
        U_dsdc_n2014), .B(debug_ref_req), .ZN(U_dsdc_n71) );
  INV_X1 U_dsdc_U124 ( .A(U_dsdc_n70), .ZN(U_dsdc_n494) );
  AOI22_X1 U_dsdc_U123 ( .A1(U_dsdc_n800), .A2(U_dsdc_bm_row_addr_0__13_), 
        .B1(U_dsdc_n814), .B2(U_dsdc_bm_row_addr_0__1_), .ZN(U_dsdc_n70) );
  AOI22_X1 U_dsdc_U122 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__12_), 
        .B1(U_dsdc_n998), .B2(U_dsdc_bm_row_addr_0__12_), .ZN(U_dsdc_n515) );
  OAI211_X1 U_dsdc_U121 ( .C1(U_dsdc_n457), .C2(U_dsdc_n63), .A(U_dsdc_n66), 
        .B(U_dsdc_n69), .ZN(U_dsdc_term_cnt_nxt[4]) );
  OAI211_X1 U_dsdc_U120 ( .C1(U_dsdc_N1991), .C2(U_dsdc_n67), .A(U_dsdc_n1379), 
        .B(U_dsdc_n68), .ZN(U_dsdc_n69) );
  NAND2_X1 U_dsdc_U119 ( .A1(U_dsdc_N1991), .A2(U_dsdc_n67), .ZN(U_dsdc_n68)
         );
  AND2_X1 U_dsdc_U118 ( .A1(U_dsdc_N1990), .A2(U_dsdc_DP_OP_1642_126_2028_n30), 
        .ZN(U_dsdc_n67) );
  AOI222_X1 U_dsdc_U117 ( .A1(n89), .A2(U_dsdc_N1991), .B1(U_dsdc_n65), .B2(
        U_dsdc_n1649), .C1(U_dsdc_n1424), .C2(U_dsdc_n1648), .ZN(U_dsdc_n66)
         );
  NOR3_X1 U_dsdc_U116 ( .A1(U_dsdc_term_cnt_3_), .A2(U_dsdc_term_cnt_4_), .A3(
        U_dsdc_term_cnt_2_), .ZN(U_dsdc_n65) );
  AOI21_X1 U_dsdc_U114 ( .B1(U_dsdc_term_cnt_3_), .B2(U_dsdc_n62), .A(
        U_dsdc_n1647), .ZN(U_dsdc_n63) );
  INV_X1 U_dsdc_U113 ( .A(U_dsdc_n1646), .ZN(U_dsdc_n62) );
  AOI22_X1 U_dsdc_U112 ( .A1(n83), .A2(U_dsdc_n60), .B1(U_cr_n128), .B2(
        U_dsdc_n59), .ZN(U_dsdc_N4321) );
  AOI22_X1 U_dsdc_U110 ( .A1(U_dsdc_bm_ras_cnt_0__2_), .A2(U_dsdc_n1182), .B1(
        U_dsdc_bm_ras_cnt_0__3_), .B2(U_dsdc_n1186), .ZN(U_dsdc_n60) );
  AOI22_X1 U_dsdc_U109 ( .A1(n83), .A2(U_dsdc_n58), .B1(n96), .B2(U_dsdc_n59), 
        .ZN(U_dsdc_N4334) );
  INV_X1 U_dsdc_U108 ( .A(n83), .ZN(U_dsdc_n59) );
  AOI22_X1 U_dsdc_U107 ( .A1(U_dsdc_bm_rc_cnt_0__2_), .A2(U_dsdc_n1175), .B1(
        U_dsdc_bm_rc_cnt_0__3_), .B2(U_dsdc_n1179), .ZN(U_dsdc_n58) );
  NAND3_X1 U_dsdc_U106 ( .A1(U_dsdc_n1170), .A2(U_dsdc_n56), .A3(U_dsdc_n57), 
        .ZN(U_dsdc_N417) );
  AOI22_X1 U_dsdc_U105 ( .A1(U_dsdc_n1121), .A2(debug_ad_col_addr_3_), .B1(
        U_dsdc_n1399), .B2(U_dsdc_n1138), .ZN(U_dsdc_n57) );
  AOI22_X1 U_dsdc_U104 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_3_), .B1(
        cr_exn_mode_value[3]), .B2(U_dsdc_n1671), .ZN(U_dsdc_n56) );
  XOR2_X1 U_dsdc_U100 ( .A(U_dsdc_n1462), .B(s_read_pipe[1]), .Z(U_dsdc_n1085)
         );
  OR4_X1 U_dsdc_U99 ( .A1(U_dsdc_bm_bank_status_3_), .A2(
        U_dsdc_bm_bank_status_2_), .A3(U_dsdc_bm_bank_status_1_), .A4(
        U_dsdc_bm_bank_status_0_), .ZN(U_dsdc_n1483) );
  AOI222_X1 U_dsdc_U98 ( .A1(U_dsdc_cas_cnt_1_), .A2(U_dsdc_n1268), .B1(
        U_dsdc_r_burst_size_1_), .B2(U_dsdc_n1269), .C1(hiu_burst_size[1]), 
        .C2(U_dsdc_n1270), .ZN(U_dsdc_n1281) );
  NOR3_X2 U_dsdc_U97 ( .A1(U_dsdc_data_cnt_0_), .A2(U_dsdc_data_cnt_1_), .A3(
        U_dsdc_n53), .ZN(U_dsdc_n740) );
  OR4_X1 U_dsdc_U96 ( .A1(U_dsdc_data_cnt_5_), .A2(U_dsdc_data_cnt_3_), .A3(
        U_dsdc_data_cnt_2_), .A4(U_dsdc_data_cnt_4_), .ZN(U_dsdc_n53) );
  INV_X1 U_dsdc_U95 ( .A(U_dsdc_n52), .ZN(U_dsdc_n477) );
  AOI222_X1 U_dsdc_U94 ( .A1(U_dsdc_n1840), .A2(U_dsdc_bm_bank_age_2__2_), 
        .B1(U_dsdc_bm_bank_age_1__2_), .B2(U_dsdc_n1839), .C1(
        U_dsdc_bm_bank_age_3__2_), .C2(U_dsdc_n476), .ZN(U_dsdc_n52) );
  AOI22_X2 U_dsdc_U92 ( .A1(debug_ad_row_addr[15]), .A2(U_dsdc_n805), .B1(
        debug_ad_row_addr[9]), .B2(U_dsdc_n802), .ZN(U_dsdc_n51) );
  AOI22_X1 U_dsdc_U91 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__2_), .B1(
        U_dsdc_n998), .B2(U_dsdc_bm_row_addr_0__2_), .ZN(U_dsdc_n562) );
  NAND3_X1 U_dsdc_U90 ( .A1(U_dsdc_n1150), .A2(U_dsdc_n49), .A3(U_dsdc_n50), 
        .ZN(U_dsdc_N413) );
  AOI22_X1 U_dsdc_U89 ( .A1(U_dsdc_n1121), .A2(debug_ad_col_addr_7_), .B1(
        U_dsdc_n1400), .B2(U_dsdc_n1138), .ZN(U_dsdc_n50) );
  AOI22_X1 U_dsdc_U88 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_7_), .B1(
        cr_exn_mode_value[7]), .B2(U_dsdc_n1671), .ZN(U_dsdc_n49) );
  OAI21_X1 U_dsdc_U87 ( .B1(U_dsdc_n1643), .B2(U_dsdc_n200), .A(U_dsdc_n48), 
        .ZN(U_dsdc_term_cnt_nxt[2]) );
  AOI21_X1 U_dsdc_U86 ( .B1(U_dsdc_N1989), .B2(n89), .A(U_dsdc_n47), .ZN(
        U_dsdc_n48) );
  OAI21_X1 U_dsdc_U85 ( .B1(U_dsdc_n1645), .B2(U_dsdc_term_cnt_2_), .A(
        U_dsdc_n46), .ZN(U_dsdc_n47) );
  AOI22_X1 U_dsdc_U84 ( .A1(U_dsdc_r_cas_latency_2_), .A2(U_dsdc_n770), .B1(
        U_dsdc_n1379), .B2(U_dsdc_n45), .ZN(U_dsdc_n46) );
  XOR2_X1 U_dsdc_U83 ( .A(U_dsdc_N1989), .B(U_dsdc_DP_OP_1642_126_2028_n31), 
        .Z(U_dsdc_n45) );
  INV_X4 U_dsdc_U82 ( .A(U_dsdc_n44), .ZN(U_dsdc_n291) );
  AOI222_X2 U_dsdc_U81 ( .A1(U_dsdc_C880_DATA5_5), .A2(U_dsdc_n1380), .B1(
        U_dsdc_N1767), .B2(U_dsdc_n1381), .C1(U_dsdc_n764), .C2(U_dsdc_n43), 
        .ZN(U_dsdc_n44) );
  XOR2_X1 U_dsdc_U80 ( .A(U_dsdc_data_cnt_5_), .B(U_dsdc_n762), .Z(U_dsdc_n43)
         );
  OAI22_X1 U_dsdc_U79 ( .A1(U_dsdc_n2073), .A2(U_dsdc_n41), .B1(U_dsdc_n42), 
        .B2(U_dsdc_n440), .ZN(U_dsdc_n281) );
  AND3_X1 U_dsdc_U78 ( .A1(U_dsdc_n2072), .A2(U_dsdc_n2071), .A3(U_dsdc_n2075), 
        .ZN(U_dsdc_n42) );
  AOI221_X1 U_dsdc_U77 ( .B1(U_dsdc_n1872), .B2(U_dsdc_n721), .C1(U_dsdc_n39), 
        .C2(U_dsdc_n721), .A(U_dsdc_n40), .ZN(U_dsdc_n41) );
  INV_X1 U_dsdc_U76 ( .A(U_dsdc_n974), .ZN(U_dsdc_n40) );
  NAND2_X1 U_dsdc_U75 ( .A1(U_dsdc_n2069), .A2(U_dsdc_n991), .ZN(U_dsdc_n39)
         );
  NOR3_X1 U_dsdc_U74 ( .A1(U_dsdc_n2064), .A2(U_dsdc_n1526), .A3(U_dsdc_n38), 
        .ZN(U_dsdc_n930) );
  NAND3_X1 U_dsdc_U73 ( .A1(U_dsdc_n2054), .A2(U_dsdc_n2060), .A3(U_dsdc_n37), 
        .ZN(U_dsdc_n38) );
  OAI21_X1 U_dsdc_U72 ( .B1(U_dsdc_n1428), .B2(U_dsdc_n896), .A(U_dsdc_n1499), 
        .ZN(U_dsdc_n37) );
  NAND3_X1 U_dsdc_U71 ( .A1(U_dsdc_n36), .A2(U_dsdc_n34), .A3(U_dsdc_n35), 
        .ZN(U_dsdc_n979) );
  NAND2_X1 U_dsdc_U70 ( .A1(U_dsdc_n1181), .A2(U_dsdc_n998), .ZN(U_dsdc_n36)
         );
  AOI22_X1 U_dsdc_U69 ( .A1(U_dsdc_n159), .A2(U_dsdc_n1209), .B1(U_dsdc_n978), 
        .B2(U_dsdc_n1237), .ZN(U_dsdc_n35) );
  AOI21_X1 U_dsdc_U68 ( .B1(U_dsdc_n1195), .B2(U_dsdc_n604), .A(U_dsdc_n1294), 
        .ZN(U_dsdc_n34) );
  INV_X1 U_dsdc_U67 ( .A(U_dsdc_n33), .ZN(U_dsdc_n495) );
  AOI22_X1 U_dsdc_U66 ( .A1(U_dsdc_n806), .A2(U_dsdc_bm_row_addr_0__15_), .B1(
        U_addrdec_n231), .B2(U_dsdc_bm_row_addr_0__11_), .ZN(U_dsdc_n33) );
  NAND3_X1 U_dsdc_U65 ( .A1(U_dsdc_n1147), .A2(U_dsdc_n31), .A3(U_dsdc_n32), 
        .ZN(U_dsdc_N411) );
  AOI22_X1 U_dsdc_U64 ( .A1(U_dsdc_n1121), .A2(debug_ad_col_addr_9_), .B1(
        U_dsdc_n1402), .B2(U_dsdc_n1138), .ZN(U_dsdc_n32) );
  AOI22_X1 U_dsdc_U63 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_9_), .B1(
        cr_exn_mode_value[9]), .B2(U_dsdc_n1671), .ZN(U_dsdc_n31) );
  NAND3_X1 U_dsdc_U62 ( .A1(U_dsdc_n1645), .A2(U_dsdc_n28), .A3(U_dsdc_n30), 
        .ZN(U_dsdc_term_cnt_nxt[1]) );
  AOI22_X1 U_dsdc_U61 ( .A1(U_dsdc_term_cnt_1_), .A2(U_dsdc_n29), .B1(
        U_dsdc_N1988), .B2(n89), .ZN(U_dsdc_n30) );
  OAI22_X1 U_dsdc_U60 ( .A1(U_dsdc_n1637), .A2(U_dsdc_n1636), .B1(U_dsdc_n1646), .B2(U_dsdc_n463), .ZN(U_dsdc_n29) );
  AOI22_X1 U_dsdc_U59 ( .A1(U_dsdc_r_cas_latency_1_), .A2(U_dsdc_n770), .B1(
        U_dsdc_n1379), .B2(U_dsdc_n27), .ZN(U_dsdc_n28) );
  XOR2_X1 U_dsdc_U58 ( .A(U_dsdc_N1987), .B(U_dsdc_N1988), .Z(U_dsdc_n27) );
  INV_X1 U_dsdc_U57 ( .A(U_dsdc_n26), .ZN(U_dsdc_n1093) );
  AOI22_X1 U_dsdc_U56 ( .A1(U_dsdc_n1084), .A2(U_dsdc_n1085), .B1(
        s_read_pipe[1]), .B2(U_dsdc_n1462), .ZN(U_dsdc_n26) );
  AOI222_X1 U_dsdc_U55 ( .A1(U_dsdc_cas_cnt_3_), .A2(U_dsdc_n1268), .B1(
        U_dsdc_r_burst_size_3_), .B2(U_dsdc_n1269), .C1(hiu_burst_size[3]), 
        .C2(U_dsdc_n1270), .ZN(U_dsdc_n1276) );
  OAI22_X1 U_dsdc_U54 ( .A1(U_dsdc_DP_OP_1642_126_2028_n28), .A2(U_dsdc_n25), 
        .B1(U_dsdc_n162), .B2(U_dsdc_n601), .ZN(U_dsdc_n163) );
  INV_X1 U_dsdc_U53 ( .A(U_dsdc_DP_OP_1642_126_2028_n11), .ZN(U_dsdc_n25) );
  NAND2_X1 U_dsdc_U52 ( .A1(U_dsdc_n937), .A2(U_dsdc_n24), .ZN(U_dsdc_n716) );
  AOI21_X1 U_dsdc_U51 ( .B1(U_dsdc_n672), .B2(U_dsdc_n759), .A(U_dsdc_n683), 
        .ZN(U_dsdc_n24) );
  AND2_X1 U_dsdc_U50 ( .A1(U_dsdc_n22), .A2(U_dsdc_n23), .ZN(U_dsdc_n884) );
  AOI22_X1 U_dsdc_U49 ( .A1(U_dsdc_n998), .A2(U_dsdc_bm_bank_status_0_), .B1(
        U_dsdc_n978), .B2(U_dsdc_bm_bank_status_3_), .ZN(U_dsdc_n23) );
  AOI22_X1 U_dsdc_U48 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_bank_status_1_), .B1(
        U_dsdc_n159), .B2(U_dsdc_bm_bank_status_2_), .ZN(U_dsdc_n22) );
  NOR4_X1 U_dsdc_U47 ( .A1(cr_do_initialize), .A2(cr_exn_mode_reg_update), 
        .A3(cr_do_self_ref_rp), .A4(cr_mode_reg_update), .ZN(U_dsdc_n1428) );
  OAI211_X1 U_dsdc_U45 ( .C1(U_dsdc_n605), .C2(U_dsdc_n1986), .A(U_dsdc_n19), 
        .B(U_dsdc_n20), .ZN(U_dsdc_N408) );
  AOI21_X1 U_dsdc_U44 ( .B1(U_dsdc_n1121), .B2(debug_ad_col_addr_11_), .A(
        U_dsdc_n1143), .ZN(U_dsdc_n20) );
  AOI22_X1 U_dsdc_U43 ( .A1(U_dsdc_n619), .A2(U_dsdc_r_col_addr_11_), .B1(
        cr_exn_mode_value[12]), .B2(U_dsdc_n1671), .ZN(U_dsdc_n19) );
  OAI221_X1 U_dsdc_U42 ( .B1(U_dsdc_n355), .B2(U_dsdc_n2069), .C1(U_dsdc_n355), 
        .C2(U_dsdc_n1417), .A(U_dsdc_n18), .ZN(U_dsdc_n[2090]) );
  NOR4_X1 U_dsdc_U41 ( .A1(U_dsdc_n1344), .A2(U_dsdc_n1412), .A3(U_dsdc_n1363), 
        .A4(U_dsdc_n17), .ZN(U_dsdc_n18) );
  OAI211_X1 U_dsdc_U40 ( .C1(U_dsdc_n2071), .C2(U_dsdc_n1805), .A(U_dsdc_n1979), .B(U_dsdc_n16), .ZN(U_dsdc_n17) );
  OR2_X1 U_dsdc_U39 ( .A1(U_dsdc_n1650), .A2(U_dsdc_n1496), .ZN(U_dsdc_n16) );
  NAND3_X1 U_dsdc_U38 ( .A1(U_dsdc_n699), .A2(U_dsdc_i_col_addr_5_), .A3(
        U_dsdc_i_col_addr_4_), .ZN(U_dsdc_n681) );
  XNOR2_X1 U_dsdc_U37 ( .A(U_dsdc_n15), .B(U_dsdc_DP_OP_1642_126_2028_n85), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n20) );
  NAND2_X1 U_dsdc_U36 ( .A1(U_dsdc_r_cas_latency_2_), .A2(U_dsdc_n753), .ZN(
        U_dsdc_n15) );
  OAI211_X1 U_dsdc_U35 ( .C1(U_dsdc_n785), .C2(U_dsdc_n800), .A(U_dsdc_n572), 
        .B(U_dsdc_n14), .ZN(U_dsdc_n492) );
  NAND2_X1 U_dsdc_U34 ( .A1(U_dsdc_n810), .A2(debug_ad_row_addr[11]), .ZN(
        U_dsdc_n14) );
  OAI211_X1 U_dsdc_U32 ( .C1(U_dsdc_term_cnt_0_), .C2(U_dsdc_n8), .A(
        U_dsdc_n11), .B(U_dsdc_n12), .ZN(U_dsdc_term_cnt_nxt[0]) );
  NAND2_X1 U_dsdc_U31 ( .A1(U_dsdc_N1987), .A2(n89), .ZN(U_dsdc_n12) );
  AOI222_X1 U_dsdc_U30 ( .A1(U_dsdc_n9), .A2(U_dsdc_n1379), .B1(
        U_dsdc_term_cnt_0_), .B2(U_dsdc_n10), .C1(U_dsdc_r_cas_latency_0_), 
        .C2(U_dsdc_n770), .ZN(U_dsdc_n11) );
  NOR2_X1 U_dsdc_U29 ( .A1(U_dsdc_n1636), .A2(U_dsdc_n1637), .ZN(U_dsdc_n10)
         );
  INV_X1 U_dsdc_U28 ( .A(U_dsdc_N1987), .ZN(U_dsdc_n9) );
  AOI21_X1 U_dsdc_U27 ( .B1(U_dsdc_n1637), .B2(U_dsdc_n1642), .A(U_dsdc_n1639), 
        .ZN(U_dsdc_n8) );
  NAND2_X1 U_dsdc_U26 ( .A1(U_dsdc_n1043), .A2(U_dsdc_n7), .ZN(U_dsdc_n1320)
         );
  NAND2_X1 U_dsdc_U25 ( .A1(U_dsdc_n6), .A2(U_dsdc_n1286), .ZN(U_dsdc_n7) );
  NAND3_X1 U_dsdc_U24 ( .A1(U_dsdc_n1041), .A2(U_dsdc_n1042), .A3(U_dsdc_n1411), .ZN(U_dsdc_n6) );
  NAND3_X2 U_dsdc_U23 ( .A1(U_dsdc_n3), .A2(U_dsdc_n717), .A3(U_dsdc_n5), .ZN(
        U_dsdc_n2007) );
  AOI211_X1 U_dsdc_U22 ( .C1(U_dsdc_n1061), .C2(U_dsdc_n1412), .A(U_dsdc_n4), 
        .B(U_dsdc_n716), .ZN(U_dsdc_n5) );
  AOI21_X1 U_dsdc_U21 ( .B1(U_dsdc_n181), .B2(U_dsdc_n1980), .A(U_dsdc_n1064), 
        .ZN(U_dsdc_n4) );
  AOI21_X1 U_dsdc_U20 ( .B1(U_dsdc_n881), .B2(U_dsdc_n2), .A(U_dsdc_n2012), 
        .ZN(U_dsdc_n3) );
  INV_X1 U_dsdc_U19 ( .A(U_dsdc_n1299), .ZN(U_dsdc_n2) );
  XNOR2_X1 U_dsdc_U18 ( .A(U_dsdc_n1), .B(U_dsdc_DP_OP_1642_126_2028_n85), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n21) );
  NAND2_X1 U_dsdc_U17 ( .A1(U_dsdc_r_cas_latency_1_), .A2(U_dsdc_n753), .ZN(
        U_dsdc_n1) );
  NOR2_X2 U_dsdc_U15 ( .A1(U_dsdc_n1124), .A2(U_dsdc_n1364), .ZN(U_dsdc_n1393)
         );
  AOI222_X1 U_dsdc_U13 ( .A1(U_dsdc_n1380), .A2(U_dsdc_C880_DATA5_3), .B1(
        U_dsdc_n1821), .B2(U_dsdc_n764), .C1(U_dsdc_n1381), .C2(U_dsdc_N1765), 
        .ZN(U_dsdc_n763) );
  AOI222_X1 U_dsdc_U12 ( .A1(U_dsdc_n1380), .A2(U_dsdc_C880_DATA5_1), .B1(
        U_dsdc_n1824), .B2(U_dsdc_n764), .C1(U_dsdc_n1381), .C2(U_dsdc_N1763), 
        .ZN(U_dsdc_n765) );
  NAND2_X2 U_dsdc_U11 ( .A1(U_dsdc_n900), .A2(U_dsdc_n983), .ZN(U_dsdc_n1286)
         );
  INV_X4 U_dsdc_U10 ( .A(U_dsdc_n621), .ZN(U_dsdc_n620) );
  AOI22_X2 U_dsdc_U9 ( .A1(U_dsdc_DP_OP_1642_126_2028_n9), .A2(U_dsdc_n163), 
        .B1(U_dsdc_DP_OP_1642_126_2028_n58), .B2(
        U_dsdc_DP_OP_1642_126_2028_n21), .ZN(U_dsdc_DP_OP_1642_126_2028_n8) );
  NAND2_X2 U_dsdc_U5 ( .A1(U_dsdc_n887), .A2(U_dsdc_n818), .ZN(U_dsdc_n914) );
  INV_X4 U_dsdc_U4 ( .A(U_dsdc_n483), .ZN(U_dsdc_n887) );
  DFFR_X2 U_dsdc_term_cnt_reg_0_ ( .D(U_dsdc_term_cnt_nxt[0]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_term_cnt_0_), .QN(U_dsdc_n463) );
  DFFR_X2 U_dsdc_r_row_addr_reg_0_ ( .D(U_dsdc_n255), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_0_), .QN(U_dsdc_n453) );
  DFFR_X2 U_dsdc_r_row_addr_reg_1_ ( .D(U_dsdc_n262), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_1_), .QN(U_dsdc_n452) );
  DFFR_X2 U_dsdc_r_row_addr_reg_2_ ( .D(U_dsdc_n263), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_2_), .QN(U_dsdc_n451) );
  DFFR_X2 U_dsdc_r_row_addr_reg_3_ ( .D(U_dsdc_n264), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_3_), .QN(U_dsdc_n450) );
  DFFR_X2 U_dsdc_r_row_addr_reg_7_ ( .D(U_dsdc_n268), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_7_), .QN(U_dsdc_n449) );
  DFFR_X2 U_dsdc_r_row_addr_reg_9_ ( .D(U_dsdc_n270), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_9_), .QN(U_dsdc_n448) );
  DFFR_X2 U_dsdc_r_row_addr_reg_11_ ( .D(U_dsdc_n257), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_11_), .QN(U_dsdc_n447) );
  DFFR_X2 U_dsdc_r_row_addr_reg_13_ ( .D(U_dsdc_n259), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_13_), .QN(U_dsdc_n454) );
  DFFR_X2 U_dsdc_r_row_addr_reg_14_ ( .D(U_dsdc_n260), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_14_), .QN(U_dsdc_n455) );
  DFFR_X2 U_dsdc_r_row_addr_reg_15_ ( .D(U_dsdc_n261), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_15_), .QN(U_dsdc_n456) );
  DFFR_X2 U_dsdc_r_burst_size_reg_3_ ( .D(U_dsdc_n274), .CK(hclk), .RN(hresetn), .Q(U_dsdc_r_burst_size_3_), .QN(U_dsdc_n299) );
  DFFR_X2 U_dsdc_r_burst_size_reg_4_ ( .D(U_dsdc_n275), .CK(hclk), .RN(hresetn), .Q(U_dsdc_r_burst_size_4_), .QN(U_dsdc_n301) );
  DFFR_X2 U_dsdc_r_burst_size_reg_5_ ( .D(U_dsdc_n276), .CK(hclk), .RN(hresetn), .Q(U_dsdc_r_burst_size_5_), .QN(U_dsdc_n172) );
  DFFR_X2 U_dsdc_r_burst_size_reg_0_ ( .D(U_dsdc_n271), .CK(hclk), .RN(hresetn), .Q(U_dsdc_r_burst_size_0_), .QN(U_dsdc_n182) );
  DFFR_X2 U_dsdc_access_cs_reg_2_ ( .D(U_dsdc_n[2090]), .CK(hclk), .RN(hresetn), .Q(U_dsdc_access_cs_2_), .QN(U_dsdc_n355) );
  DFFR_X2 U_dsdc_r_wrapped_burst_reg ( .D(U_dsdc_n277), .CK(hclk), .RN(hresetn), .Q(U_dsdc_r_wrapped_burst), .QN(U_dsdc_n328) );
  DFFR_X2 U_dsdc_i_col_addr_reg_1_ ( .D(U_dsdc_n319), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_i_col_addr_1_), .QN(U_dsdc_n354) );
  DFFR_X2 U_dsdc_i_col_addr_reg_13_ ( .D(U_dsdc_i_col_addr_nxt[13]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_i_col_addr_13_), .QN(U_dsdc_n446) );
  DFFR_X2 U_dsdc_delta_delay_reg_0_ ( .D(U_dsdc_n216), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_delta_delay_0_), .QN(U_dsdc_n461) );
  DFFR_X2 U_dsdc_early_term_flag_reg ( .D(U_dsdc_n282), .CK(hclk), .RN(hresetn), .Q(U_dsdc_early_term_flag), .QN(U_dsdc_n306) );
  DFFR_X2 U_dsdc_data_flag_reg ( .D(U_dsdc_n281), .CK(hclk), .RN(hresetn), .Q(
        U_dsdc_data_flag), .QN(U_dsdc_n440) );
  DFFR_X2 U_dsdc_rcar_cnt2_reg_3_ ( .D(U_dsdc_rcar_cnt2_nxt[3]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_rcar_cnt2_3_), .QN(U_dsdc_n430) );
  DFFR_X2 U_dsdc_mrd_cnt_reg_0_ ( .D(U_dsdc_N4174), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_mrd_cnt_0_), .QN(U_dsdc_n199) );
  DFFR_X2 U_dsdc_mrd_cnt_reg_1_ ( .D(U_dsdc_n423), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_mrd_cnt_1_), .QN(U_dsdc_n429) );
  DFFR_X2 U_dsdc_num_init_ref_cnt_reg_2_ ( .D(U_dsdc_num_init_ref_cnt_nxt[2]), 
        .CK(hclk), .RN(hresetn), .Q(U_dsdc_num_init_ref_cnt_2_), .QN(
        U_dsdc_n473) );
  DFFR_X2 U_dsdc_rp_cnt1_reg_0_ ( .D(U_dsdc_rp_cnt1_nxt[0]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_rp_cnt1_0_), .QN(U_dsdc_n169) );
  DFFR_X2 U_dsdc_rp_cnt1_reg_2_ ( .D(U_dsdc_rp_cnt1_nxt[2]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_rp_cnt1_2_), .QN(U_dsdc_n427) );
  DFFR_X2 U_dsdc_rp_cnt1_reg_1_ ( .D(U_dsdc_rp_cnt1_nxt[1]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_rp_cnt1_1_), .QN(U_dsdc_n198) );
  DFFR_X2 U_dsdc_r_cas_latency_reg_0_ ( .D(U_dsdc_add_x_2600_1_n8), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_r_cas_latency_0_), .QN(U_dsdc_n342) );
  DFFR_X2 U_dsdc_bm_num_open_bank_reg_3_ ( .D(U_dsdc_n296), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_num_open_bank_3_), .QN(U_dsdc_n179) );
  DFFR_X2 U_dsdc_operation_cs_reg_3_ ( .D(U_dsdc_n2094), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_operation_cs_3_), .QN(U_dsdc_n196) );
  DFFR_X2 U_dsdc_row_cnt_reg_12_ ( .D(U_dsdc_n369), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_12_), .QN(U_dsdc_n203) );
  DFFR_X2 U_dsdc_bm_bank_age_reg_0__0_ ( .D(U_dsdc_n283), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_0__0_), .QN(U_dsdc_n201) );
  DFFR_X2 U_dsdc_bm_bank_age_reg_2__2_ ( .D(U_dsdc_n211), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_2__2_), .QN(U_dsdc_n336) );
  DFFR_X2 U_dsdc_data_cnt_reg_1_ ( .D(U_dsdc_n287), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_data_cnt_1_), .QN(U_dsdc_n436) );
  DFFR_X2 U_dsdc_bm_bank_age_reg_2__0_ ( .D(U_dsdc_n209), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_2__0_), .QN(U_dsdc_n353) );
  DFFR_X2 U_dsdc_bm_bank_age_reg_1__0_ ( .D(U_dsdc_n223), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_1__0_), .QN(U_dsdc_n352) );
  DFFR_X2 U_dsdc_wrapped_pop_flag_reg ( .D(U_dsdc_wrapped_pop_flag_nxt), .CK(
        hclk), .RN(hresetn), .Q(U_dsdc_wrapped_pop_flag) );
  DFFR_X2 U_dsdc_num_init_ref_cnt_reg_0_ ( .D(U_dsdc_num_init_ref_cnt_nxt[0]), 
        .CK(hclk), .RN(hresetn), .Q(U_dsdc_num_init_ref_cnt_0_) );
  DFFR_X2 U_dsdc_s_rd_end_reg ( .D(U_dsdc_s_rd_end_nxt), .CK(hclk), .RN(
        hresetn), .Q(s_rd_end) );
  DFFR_X2 U_dsdc_num_init_ref_cnt_reg_1_ ( .D(U_dsdc_num_init_ref_cnt_nxt[1]), 
        .CK(hclk), .RN(hresetn), .Q(U_dsdc_num_init_ref_cnt_1_) );
  DFFR_X2 U_dsdc_dout_valid_flag_reg ( .D(U_dsdc_n232), .CK(hclk), .RN(hresetn), .QN(U_dsdc_n466) );
  DFFR_X2 U_dsdc_rp_cnt2_reg_0_ ( .D(U_dsdc_rp_cnt2_nxt[0]), .CK(hclk), .RN(
        hresetn), .QN(U_dsdc_n171) );
  DFFR_X2 U_dsdc_write_start_reg ( .D(U_dsdc_write_start_nxt), .CK(hclk), .RN(
        hresetn), .QN(U_dsdc_n433) );
  DFFR_X2 U_dsdc_rcd_cnt_reg_1_ ( .D(U_dsdc_N4140), .CK(hclk), .RN(hresetn), 
        .QN(U_dsdc_n326) );
  DFFR_X2 U_dsdc_wtr_cnt_reg_1_ ( .D(U_dsdc_wtr_cnt_nxt[1]), .CK(hclk), .RN(
        hresetn), .QN(U_dsdc_n194) );
  DFFR_X2 U_dsdc_cas_cnt_reg_0_ ( .D(U_dsdc_cas_cnt_nxt[0]), .CK(hclk), .RN(
        hresetn), .QN(U_dsdc_n327) );
  DFFR_X2 U_dsdc_i_col_addr_reg_3_ ( .D(U_dsdc_n321), .CK(hclk), .RN(hresetn), 
        .QN(U_dsdc_n443) );
  DFFR_X2 U_dsdc_i_col_addr_reg_10_ ( .D(U_dsdc_n316), .CK(hclk), .RN(hresetn), 
        .QN(U_dsdc_n444) );
  DFFR_X2 U_dsdc_xsr_cnt_reg_6_ ( .D(U_dsdc_n392), .CK(hclk), .RN(hresetn), 
        .QN(U_dsdc_n359) );
  DFFR_X2 U_dsdc_terminate_reg ( .D(hiu_terminate), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_n165), .QN(U_dsdc_n181) );
  XOR2_X1 U_dsdc_DP_OP_1642_126_2028_U42 ( .A(U_dsdc_DP_OP_1642_126_2028_n30), 
        .B(U_dsdc_N1990), .Z(U_dsdc_N2002) );
  AND2_X2 U_dsdc_DP_OP_1642_126_2028_U45 ( .A1(U_dsdc_N1989), .A2(
        U_dsdc_DP_OP_1642_126_2028_n31), .ZN(U_dsdc_DP_OP_1642_126_2028_n30)
         );
  AND2_X2 U_dsdc_DP_OP_1642_126_2028_U47 ( .A1(U_dsdc_N1988), .A2(U_dsdc_N1987), .ZN(U_dsdc_DP_OP_1642_126_2028_n31) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U1 ( .A(U_dsdc_DP_OP_1642_126_2028_n1), 
        .B(U_dsdc_DP_OP_1642_126_2028_n12), .Z(U_dsdc_C880_DATA5_5) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U2 ( .A(U_dsdc_DP_OP_1642_126_2028_n85), 
        .B(U_dsdc_DP_OP_1642_126_2028_n62), .Z(U_dsdc_DP_OP_1642_126_2028_n1)
         );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U6 ( .A(U_dsdc_DP_OP_1642_126_2028_n85), 
        .B(U_dsdc_DP_OP_1642_126_2028_n61), .Z(U_dsdc_DP_OP_1642_126_2028_n3)
         );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U7 ( .A(U_dsdc_DP_OP_1642_126_2028_n14), 
        .B(U_dsdc_DP_OP_1642_126_2028_n5), .Z(U_dsdc_C880_DATA5_3) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U10 ( .A(U_dsdc_DP_OP_1642_126_2028_n19), 
        .B(U_dsdc_DP_OP_1642_126_2028_n60), .Z(U_dsdc_DP_OP_1642_126_2028_n5)
         );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U14 ( .A(U_dsdc_DP_OP_1642_126_2028_n20), 
        .B(U_dsdc_DP_OP_1642_126_2028_n59), .Z(U_dsdc_DP_OP_1642_126_2028_n7)
         );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U15 ( .A(U_dsdc_n163), .B(
        U_dsdc_DP_OP_1642_126_2028_n9), .Z(U_dsdc_C880_DATA5_1) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U18 ( .A(U_dsdc_DP_OP_1642_126_2028_n21), 
        .B(U_dsdc_DP_OP_1642_126_2028_n58), .Z(U_dsdc_DP_OP_1642_126_2028_n9)
         );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U51 ( .A(U_dsdc_DP_OP_1642_126_2028_n34), 
        .B(U_dsdc_DP_OP_1642_126_2028_n42), .Z(U_dsdc_N1766) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U54 ( .A(hiu_burst_size[4]), .B(
        U_dsdc_N1991), .Z(U_dsdc_DP_OP_1642_126_2028_n34) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U55 ( .A(U_dsdc_DP_OP_1642_126_2028_n36), 
        .B(U_dsdc_DP_OP_1642_126_2028_n43), .Z(U_dsdc_N1765) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U58 ( .A(hiu_burst_size[3]), .B(
        U_dsdc_N1990), .Z(U_dsdc_DP_OP_1642_126_2028_n36) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U59 ( .A(U_dsdc_DP_OP_1642_126_2028_n44), 
        .B(U_dsdc_DP_OP_1642_126_2028_n38), .Z(U_dsdc_N1764) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U62 ( .A(hiu_burst_size[2]), .B(
        U_dsdc_N1989), .Z(U_dsdc_DP_OP_1642_126_2028_n38) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U63 ( .A(U_dsdc_DP_OP_1642_126_2028_n45), 
        .B(U_dsdc_DP_OP_1642_126_2028_n40), .Z(U_dsdc_N1763) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U66 ( .A(hiu_burst_size[1]), .B(
        U_dsdc_N1988), .Z(U_dsdc_DP_OP_1642_126_2028_n40) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U67 ( .A(hiu_burst_size[0]), .B(
        U_dsdc_N1987), .Z(U_dsdc_N1762) );
  AND2_X4 U_dsdc_DP_OP_1642_126_2028_U68 ( .A1(U_dsdc_N1987), .A2(
        hiu_burst_size[0]), .ZN(U_dsdc_DP_OP_1642_126_2028_n45) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U69 ( .A(U_dsdc_r_cas_latency_3_), .B(
        U_dsdc_DP_OP_1642_126_2028_n50), .Z(U_dsdc_N1990) );
  AND2_X4 U_dsdc_DP_OP_1642_126_2028_U70 ( .A1(U_dsdc_DP_OP_1642_126_2028_n50), 
        .A2(U_dsdc_r_cas_latency_3_), .ZN(U_dsdc_N1991) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U71 ( .A(U_dsdc_DP_OP_1642_126_2028_n47), 
        .B(U_dsdc_DP_OP_1642_126_2028_n51), .Z(U_dsdc_N1989) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U74 ( .A(U_dsdc_delta_delay_2_), .B(
        U_dsdc_r_cas_latency_2_), .Z(U_dsdc_DP_OP_1642_126_2028_n47) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U75 ( .A(U_dsdc_DP_OP_1642_126_2028_n52), 
        .B(U_dsdc_DP_OP_1642_126_2028_n49), .Z(U_dsdc_N1988) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U78 ( .A(U_dsdc_delta_delay_1_), .B(
        U_dsdc_r_cas_latency_1_), .Z(U_dsdc_DP_OP_1642_126_2028_n49) );
  XOR2_X2 U_dsdc_DP_OP_1642_126_2028_U79 ( .A(U_dsdc_delta_delay_0_), .B(
        U_dsdc_r_cas_latency_0_), .Z(U_dsdc_N1987) );
  AND2_X4 U_dsdc_DP_OP_1642_126_2028_U80 ( .A1(U_dsdc_r_cas_latency_0_), .A2(
        U_dsdc_delta_delay_0_), .ZN(U_dsdc_DP_OP_1642_126_2028_n52) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U77 ( .A1(U_dsdc_DP_OP_1642_126_2028_n49), .A2(U_dsdc_DP_OP_1642_126_2028_n52), .B1(U_dsdc_r_cas_latency_1_), .B2(
        U_dsdc_delta_delay_1_), .ZN(U_dsdc_DP_OP_1642_126_2028_n48) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U76 ( .A(U_dsdc_DP_OP_1642_126_2028_n48), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n51) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U65 ( .A1(U_dsdc_DP_OP_1642_126_2028_n40), .A2(U_dsdc_DP_OP_1642_126_2028_n45), .B1(U_dsdc_N1988), .B2(
        hiu_burst_size[1]), .ZN(U_dsdc_DP_OP_1642_126_2028_n39) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U64 ( .A(U_dsdc_DP_OP_1642_126_2028_n39), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n44) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U61 ( .A1(U_dsdc_DP_OP_1642_126_2028_n38), .A2(U_dsdc_DP_OP_1642_126_2028_n44), .B1(U_dsdc_N1989), .B2(
        hiu_burst_size[2]), .ZN(U_dsdc_DP_OP_1642_126_2028_n37) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U60 ( .A(U_dsdc_DP_OP_1642_126_2028_n37), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n43) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U73 ( .A1(U_dsdc_DP_OP_1642_126_2028_n51), .A2(U_dsdc_DP_OP_1642_126_2028_n47), .B1(U_dsdc_r_cas_latency_2_), .B2(
        U_dsdc_delta_delay_2_), .ZN(U_dsdc_DP_OP_1642_126_2028_n46) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U72 ( .A(U_dsdc_DP_OP_1642_126_2028_n46), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n50) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U57 ( .A1(U_dsdc_DP_OP_1642_126_2028_n43), .A2(U_dsdc_DP_OP_1642_126_2028_n36), .B1(U_dsdc_N1990), .B2(
        hiu_burst_size[3]), .ZN(U_dsdc_DP_OP_1642_126_2028_n35) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U56 ( .A(U_dsdc_DP_OP_1642_126_2028_n35), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n42) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U29 ( .A1(U_dsdc_N1767), .A2(
        U_dsdc_DP_OP_1642_126_2028_I4), .B1(U_dsdc_DP_OP_1642_126_2028_I6), 
        .B2(U_dsdc_DP_OP_1642_126_2028_I5_5_), .ZN(
        U_dsdc_DP_OP_1642_126_2028_n23) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U30 ( .A(U_dsdc_DP_OP_1642_126_2028_n23), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n62) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U34 ( .A1(U_dsdc_N1765), .A2(
        U_dsdc_DP_OP_1642_126_2028_I4), .B1(U_dsdc_DP_OP_1642_126_2028_I6), 
        .B2(U_dsdc_DP_OP_1642_126_2028_I5_3_), .ZN(
        U_dsdc_DP_OP_1642_126_2028_n25) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U33 ( .A(U_dsdc_DP_OP_1642_126_2028_n25), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n60) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U36 ( .A1(U_dsdc_N1764), .A2(
        U_dsdc_DP_OP_1642_126_2028_I4), .B1(U_dsdc_DP_OP_1642_126_2028_I6), 
        .B2(U_dsdc_DP_OP_1642_126_2028_I5_2_), .ZN(
        U_dsdc_DP_OP_1642_126_2028_n26) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U35 ( .A(U_dsdc_DP_OP_1642_126_2028_n26), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n59) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U38 ( .A1(U_dsdc_N1763), .A2(
        U_dsdc_DP_OP_1642_126_2028_I4), .B1(U_dsdc_DP_OP_1642_126_2028_I6), 
        .B2(U_dsdc_DP_OP_1642_126_2028_I5_1_), .ZN(
        U_dsdc_DP_OP_1642_126_2028_n27) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U37 ( .A(U_dsdc_DP_OP_1642_126_2028_n27), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n58) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U40 ( .A1(U_dsdc_N1762), .A2(
        U_dsdc_DP_OP_1642_126_2028_I4), .B1(U_dsdc_DP_OP_1642_126_2028_I6), 
        .B2(U_dsdc_DP_OP_1642_126_2028_I5_0_), .ZN(
        U_dsdc_DP_OP_1642_126_2028_n28) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U16 ( .A(U_dsdc_DP_OP_1642_126_2028_n8), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n15) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U12 ( .A(U_dsdc_DP_OP_1642_126_2028_n6), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n14) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U8 ( .A(U_dsdc_DP_OP_1642_126_2028_n4), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n13) );
  AOI22_X2 U_dsdc_DP_OP_1642_126_2028_U32 ( .A1(U_dsdc_N1766), .A2(
        U_dsdc_DP_OP_1642_126_2028_I4), .B1(U_dsdc_DP_OP_1642_126_2028_I6), 
        .B2(U_dsdc_DP_OP_1642_126_2028_I5_4_), .ZN(
        U_dsdc_DP_OP_1642_126_2028_n24) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U31 ( .A(U_dsdc_DP_OP_1642_126_2028_n24), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n61) );
  INV_X4 U_dsdc_DP_OP_1642_126_2028_U4 ( .A(U_dsdc_DP_OP_1642_126_2028_n2), 
        .ZN(U_dsdc_DP_OP_1642_126_2028_n12) );
  DFFR_X2 U_dsdc_miu_push_n_reg ( .D(U_dsdc_n329), .CK(hclk), .RN(hresetn), 
        .Q(n82), .QN(ctl_push_n) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_2__1_ ( .D(U_dsdc_n210), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_2__1_), .QN(U_dsdc_n178) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_2__3_ ( .D(U_dsdc_n212), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_2__3_), .QN(U_dsdc_n459) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_2__4_ ( .D(U_dsdc_n213), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_2__4_), .QN(U_dsdc_n350) );
  DFFR_X1 U_dsdc_ref_ack_reg ( .D(U_dsdc_N430), .CK(hclk), .RN(hresetn), .Q(
        ctl_ref_ack) );
  DFFR_X1 U_dsdc_s_rd_pop_reg ( .D(U_dsdc_n329), .CK(hclk), .RN(hresetn), .Q(
        s_rd_pop) );
  DFFR_X1 U_dsdc_data_cnt_reg_5_ ( .D(U_dsdc_n291), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_data_cnt_5_) );
  DFFR_X1 U_dsdc_data_cnt_reg_4_ ( .D(U_dsdc_n290), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_data_cnt_4_) );
  DFFR_X1 U_dsdc_data_cnt_reg_3_ ( .D(U_dsdc_n289), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_data_cnt_3_), .QN(U_dsdc_n437) );
  DFFR_X1 U_dsdc_data_cnt_reg_2_ ( .D(U_dsdc_n288), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_data_cnt_2_) );
  DFFR_X1 U_dsdc_term_cnt_reg_1_ ( .D(U_dsdc_term_cnt_nxt[1]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_term_cnt_1_) );
  DFFR_X1 U_dsdc_term_cnt_reg_2_ ( .D(U_dsdc_term_cnt_nxt[2]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_term_cnt_2_), .QN(U_dsdc_n200) );
  DFFR_X1 U_dsdc_term_cnt_reg_3_ ( .D(U_dsdc_term_cnt_nxt[3]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_term_cnt_3_) );
  DFFS_X2 U_dsdc_s_cs_n_reg_0_ ( .D(U_dsdc_N401), .CK(hclk), .SN(hresetn), 
        .QN(ctl_chip_select_0_) );
  DFFS_X2 U_dsdc_s_ras_n_reg ( .D(U_dsdc_N402), .CK(hclk), .SN(hresetn), .Q(
        s_ras_n) );
  DFFS_X2 U_dsdc_s_we_n_reg ( .D(U_dsdc_N404), .CK(hclk), .SN(hresetn), .Q(
        s_we_n) );
  DFFS_X2 U_dsdc_s_cas_n_reg ( .D(U_dsdc_N403), .CK(hclk), .SN(hresetn), .Q(
        s_cas_n) );
  DFFS_X2 U_dsdc_miu_pop_n_reg ( .D(U_dsdc_N429), .CK(hclk), .SN(hresetn), .Q(
        ctl_pop_n) );
  DFFS_X2 U_dsdc_i_dqs_d_reg ( .D(U_dsdc_i_dqs), .CK(hclk), .SN(hresetn), .Q(
        U_dsdc_i_dqs_d) );
  DFFS_X2 U_dsdc_i_dqs_reg ( .D(U_dsdc_i_dqs_nxt), .CK(hclk), .SN(hresetn), 
        .Q(U_dsdc_i_dqs) );
  DFFS_X2 U_dsdc_pre_amble_reg ( .D(U_dsdc_pre_amble_nxt), .CK(hclk), .SN(
        hresetn), .QN(pre_amble) );
  DFFS_X2 U_dsdc_s_dout_valid_reg_1_ ( .D(U_dsdc_s_dout_valid_nxt), .CK(hclk), 
        .SN(hresetn), .Q(s_dout_valid[1]) );
  DFFS_X2 U_dsdc_s_dout_valid_reg_0_ ( .D(U_dsdc_s_dout_valid_nxt), .CK(hclk), 
        .SN(hresetn), .Q(s_dout_valid[0]) );
  DFFR_X1 U_dsdc_delta_delay_reg_2_ ( .D(U_dsdc_n214), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_delta_delay_2_), .QN(U_dsdc_n467) );
  DFFR_X1 U_dsdc_delta_delay_reg_1_ ( .D(U_dsdc_n215), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_delta_delay_1_), .QN(U_dsdc_n464) );
  DFFR_X1 U_dsdc_pre_rd_dqs_mask_reg ( .D(U_dsdc_n217), .CK(hclk), .RN(hresetn), .Q(pre_rd_dqs_mask), .QN(U_dsdc_n475) );
  DFFR_X1 U_dsdc_dqs_mask_end_reg ( .D(U_dsdc_dqs_mask_end_nxt), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_dqs_mask_end) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_3__0_ ( .D(U_dsdc_n218), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_3__0_), .QN(U_dsdc_n304) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_3__1_ ( .D(U_dsdc_n219), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_3__1_), .QN(U_dsdc_n302) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_3__2_ ( .D(U_dsdc_n220), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_3__2_), .QN(U_dsdc_n303) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_3__3_ ( .D(U_dsdc_n221), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_3__3_), .QN(U_dsdc_n284) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_3__4_ ( .D(U_dsdc_n222), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_3__4_), .QN(U_dsdc_n351) );
  DFFR_X1 U_dsdc_bm_bank_status_reg_3_ ( .D(U_dsdc_N4496), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_status_3_), .QN(U_dsdc_n396) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_1__1_ ( .D(U_dsdc_n224), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_1__1_), .QN(U_dsdc_n335) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_1__2_ ( .D(U_dsdc_n225), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_1__2_), .QN(U_dsdc_n337) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_1__3_ ( .D(U_dsdc_n226), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_1__3_), .QN(U_dsdc_n460) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_1__4_ ( .D(U_dsdc_n227), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_1__4_), .QN(U_dsdc_n349) );
  DFFR_X1 U_dsdc_bm_bank_status_reg_1_ ( .D(U_dsdc_N4402), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_status_1_), .QN(U_dsdc_n383) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_0__1_ ( .D(U_dsdc_n228), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_0__1_), .QN(U_dsdc_n435) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_0__2_ ( .D(U_dsdc_n229), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_0__2_), .QN(U_dsdc_n334) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_0__3_ ( .D(U_dsdc_n230), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_0__3_), .QN(U_dsdc_n458) );
  DFFR_X1 U_dsdc_bm_bank_age_reg_0__4_ ( .D(U_dsdc_n231), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_age_0__4_), .QN(U_dsdc_n434) );
  DFFR_X1 U_dsdc_bm_bank_status_reg_0_ ( .D(U_dsdc_N4355), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_status_0_), .QN(U_dsdc_n384) );
  DFFR_X1 U_dsdc_bm_num_open_bank_reg_0_ ( .D(U_dsdc_n293), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_num_open_bank_0_), .QN(U_dsdc_n340) );
  DFFR_X1 U_dsdc_bm_num_open_bank_reg_1_ ( .D(U_dsdc_n294), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_num_open_bank_1_), .QN(U_dsdc_n180) );
  DFFR_X1 U_dsdc_bm_num_open_bank_reg_2_ ( .D(U_dsdc_n295), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_num_open_bank_2_), .QN(U_dsdc_n338) );
  DFFR_X1 U_dsdc_bm_num_open_bank_reg_4_ ( .D(U_dsdc_n297), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_num_open_bank_4_), .QN(U_dsdc_n385) );
  DFFR_X1 U_dsdc_s_addr_reg_10_ ( .D(U_dsdc_N410), .CK(hclk), .RN(hresetn), 
        .Q(s_addr[10]) );
  DFFS_X2 U_dsdc_r_bm_close_all_reg ( .D(U_dsdc_n1394), .CK(hclk), .SN(hresetn), .QN(U_dsdc_r_bm_close_all) );
  DFFR_X1 U_dsdc_i_col_addr_reg_0_ ( .D(U_dsdc_n315), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_N1685) );
  DFFR_X1 U_dsdc_i_col_addr_reg_11_ ( .D(U_dsdc_n317), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_i_col_addr_11_) );
  DFFR_X1 U_dsdc_i_col_addr_reg_12_ ( .D(U_dsdc_i_col_addr_nxt[12]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_i_col_addr_12_) );
  DFFR_X1 U_dsdc_i_col_addr_reg_14_ ( .D(U_dsdc_i_col_addr_nxt[14]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_i_col_addr_14_) );
  DFFS_X2 U_dsdc_pre_amble_mute_reg ( .D(U_dsdc_n348), .CK(hclk), .SN(hresetn), 
        .QN(U_dsdc_pre_amble_mute) );
  DFFR_X1 U_dsdc_pre_dqm_reg_0_ ( .D(U_dsdc_N425), .CK(hclk), .RN(hresetn), 
        .Q(pre_dqm[0]) );
  DFFR_X1 U_dsdc_pre_dqm_reg_1_ ( .D(U_dsdc_N426), .CK(hclk), .RN(hresetn), 
        .Q(pre_dqm[1]) );
  DFFR_X1 U_dsdc_pre_dqm_reg_2_ ( .D(U_dsdc_N427), .CK(hclk), .RN(hresetn), 
        .Q(pre_dqm[2]) );
  DFFR_X1 U_dsdc_pre_dqm_reg_3_ ( .D(U_dsdc_N428), .CK(hclk), .RN(hresetn), 
        .Q(pre_dqm[3]) );
  DFFR_X1 U_dsdc_s_addr_reg_12_ ( .D(U_dsdc_N408), .CK(hclk), .RN(hresetn), 
        .Q(s_addr[12]) );
  DFFR_X1 U_dsdc_s_addr_reg_11_ ( .D(U_dsdc_N409), .CK(hclk), .RN(hresetn), 
        .Q(s_addr[11]) );
  DFFR_X1 U_dsdc_s_addr_reg_9_ ( .D(U_dsdc_N411), .CK(hclk), .RN(hresetn), .Q(
        s_addr[9]) );
  DFFR_X1 U_dsdc_s_addr_reg_8_ ( .D(U_dsdc_N412), .CK(hclk), .RN(hresetn), .Q(
        s_addr[8]) );
  DFFR_X1 U_dsdc_cas_latency_cnt_reg_2_ ( .D(U_dsdc_N4128), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_cas_latency_cnt_2_), .QN(U_dsdc_n331) );
  DFFR_X1 U_dsdc_cas_latency_cnt_reg_1_ ( .D(U_dsdc_N4127), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_cas_latency_cnt_1_) );
  DFFR_X1 U_dsdc_cas_latency_cnt_reg_0_ ( .D(U_dsdc_n300), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_cas_latency_cnt_0_) );
  DFFR_X1 U_dsdc_cas_latency_cnt_reg_3_ ( .D(U_dsdc_N4129), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_cas_latency_cnt_3_) );
  DFFS_X2 U_dsdc_s_rd_start_reg ( .D(U_dsdc_n1393), .CK(hclk), .SN(hresetn), 
        .QN(s_rd_start) );
  DFFR_X1 U_dsdc_s_addr_reg_7_ ( .D(U_dsdc_N413), .CK(hclk), .RN(hresetn), .Q(
        s_addr[7]) );
  DFFR_X1 U_dsdc_s_addr_reg_6_ ( .D(U_dsdc_N414), .CK(hclk), .RN(hresetn), .Q(
        s_addr[6]) );
  DFFR_X1 U_dsdc_i_col_addr_reg_6_ ( .D(U_dsdc_i_col_addr_nxt[6]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_i_col_addr_6_) );
  DFFR_X1 U_dsdc_s_addr_reg_5_ ( .D(U_dsdc_N415), .CK(hclk), .RN(hresetn), .Q(
        s_addr[5]) );
  DFFR_X1 U_dsdc_i_col_addr_reg_5_ ( .D(U_dsdc_i_col_addr_nxt[5]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_i_col_addr_5_) );
  DFFR_X1 U_dsdc_s_addr_reg_4_ ( .D(U_dsdc_N416), .CK(hclk), .RN(hresetn), .Q(
        s_addr[4]) );
  DFFR_X1 U_dsdc_i_col_addr_reg_4_ ( .D(U_dsdc_i_col_addr_nxt[4]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_i_col_addr_4_) );
  DFFR_X1 U_dsdc_s_addr_reg_3_ ( .D(U_dsdc_N417), .CK(hclk), .RN(hresetn), .Q(
        s_addr[3]) );
  DFFR_X1 U_dsdc_s_addr_reg_2_ ( .D(U_dsdc_N418), .CK(hclk), .RN(hresetn), .Q(
        s_addr[2]) );
  DFFR_X1 U_dsdc_s_addr_reg_1_ ( .D(U_dsdc_N419), .CK(hclk), .RN(hresetn), .Q(
        s_addr[1]) );
  DFFR_X1 U_dsdc_s_addr_reg_0_ ( .D(U_dsdc_N420), .CK(hclk), .RN(hresetn), .Q(
        s_addr[0]) );
  DFFR_X1 U_dsdc_s_bank_addr_reg_0_ ( .D(U_dsdc_N422), .CK(hclk), .RN(hresetn), 
        .Q(s_bank_addr[0]) );
  DFFR_X1 U_dsdc_s_bank_addr_reg_1_ ( .D(U_dsdc_s_bank_addr_nxt_a_1_), .CK(
        hclk), .RN(hresetn), .Q(s_bank_addr[1]) );
  DFFR_X1 U_dsdc_s_addr_reg_13_ ( .D(U_dsdc_s_addr_nxt_a[13]), .CK(hclk), .RN(
        hresetn), .Q(s_addr[13]) );
  DFFR_X1 U_dsdc_s_addr_reg_14_ ( .D(U_dsdc_s_addr_nxt_a[14]), .CK(hclk), .RN(
        hresetn), .Q(s_addr[14]) );
  DFFR_X1 U_dsdc_s_addr_reg_15_ ( .D(U_dsdc_s_addr_nxt_a[15]), .CK(hclk), .RN(
        hresetn), .Q(s_addr[15]) );
  DFFR_X1 U_dsdc_i_col_addr_reg_2_ ( .D(U_dsdc_n320), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_i_col_addr_2_) );
  DFFR_X1 U_dsdc_i_col_addr_reg_7_ ( .D(U_dsdc_n322), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_i_col_addr_7_) );
  DFFR_X1 U_dsdc_i_col_addr_reg_8_ ( .D(U_dsdc_n323), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_i_col_addr_8_) );
  DFFR_X1 U_dsdc_i_col_addr_reg_9_ ( .D(U_dsdc_n324), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_i_col_addr_9_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__12_ ( .D(U_dsdc_N4348), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__12_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__12_ ( .D(U_dsdc_N4395), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__12_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__12_ ( .D(U_dsdc_N4442), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__12_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__12_ ( .D(U_dsdc_N4489), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__12_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__11_ ( .D(U_dsdc_N4347), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__11_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__11_ ( .D(U_dsdc_N4394), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__11_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__11_ ( .D(U_dsdc_N4441), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__11_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__11_ ( .D(U_dsdc_N4488), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__11_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__10_ ( .D(U_dsdc_N4346), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__10_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__10_ ( .D(U_dsdc_N4393), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__10_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__10_ ( .D(U_dsdc_N4440), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__10_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__10_ ( .D(U_dsdc_N4487), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__10_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__9_ ( .D(U_dsdc_N4345), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__9_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__9_ ( .D(U_dsdc_N4392), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__9_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__9_ ( .D(U_dsdc_N4439), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__9_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__9_ ( .D(U_dsdc_N4486), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__9_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__8_ ( .D(U_dsdc_N4344), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__8_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__8_ ( .D(U_dsdc_N4391), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__8_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__8_ ( .D(U_dsdc_N4438), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__8_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__8_ ( .D(U_dsdc_N4485), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__8_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__7_ ( .D(U_dsdc_N4343), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__7_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__7_ ( .D(U_dsdc_N4390), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__7_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__7_ ( .D(U_dsdc_N4437), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__7_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__7_ ( .D(U_dsdc_N4484), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__7_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_0_ ( .D(U_dsdc_n233), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_0_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_10_ ( .D(U_dsdc_n234), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_10_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_11_ ( .D(U_dsdc_n235), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_11_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_12_ ( .D(U_dsdc_n236), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_12_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_13_ ( .D(U_dsdc_n237), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_13_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_14_ ( .D(U_dsdc_n238), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_14_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_1_ ( .D(U_dsdc_n240), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_1_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_2_ ( .D(U_dsdc_n241), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_2_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_3_ ( .D(U_dsdc_n242), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_3_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_4_ ( .D(U_dsdc_n243), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_4_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_5_ ( .D(U_dsdc_n244), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_5_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_6_ ( .D(U_dsdc_n245), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_6_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_7_ ( .D(U_dsdc_n246), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_7_) );
  DFFR_X1 U_dsdc_r_col_addr_reg_8_ ( .D(U_dsdc_n247), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_8_), .QN(U_dsdc_n445) );
  DFFR_X1 U_dsdc_r_col_addr_reg_9_ ( .D(U_dsdc_n248), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_col_addr_9_) );
  DFFR_X1 U_dsdc_bm_ras_cnt_max_reg_2_ ( .D(U_dsdc_N4283), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_max_2_), .QN(U_dsdc_n428) );
  DFFR_X1 U_dsdc_bm_ras_cnt_max_reg_1_ ( .D(U_dsdc_N4282), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_max_1_) );
  DFFR_X1 U_dsdc_bm_ras_cnt_max_reg_0_ ( .D(U_dsdc_N4281), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_max_0_) );
  DFFR_X1 U_dsdc_bm_ras_cnt_max_reg_3_ ( .D(U_dsdc_N4284), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_max_3_) );
  DFFR_X1 U_dsdc_rcd_cnt_reg_0_ ( .D(U_dsdc_N4139), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_rcd_cnt_0_), .QN(U_dsdc_n174) );
  DFFR_X1 U_dsdc_rcd_cnt_reg_2_ ( .D(U_dsdc_N4141), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_rcd_cnt_2_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__15_ ( .D(U_dsdc_N4351), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__15_), .QN(U_dsdc_n425) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__14_ ( .D(U_dsdc_N4350), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__14_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__13_ ( .D(U_dsdc_N4349), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__13_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__6_ ( .D(U_dsdc_N4342), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__6_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__5_ ( .D(U_dsdc_N4341), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__5_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__4_ ( .D(U_dsdc_N4340), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__4_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__3_ ( .D(U_dsdc_N4339), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__3_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__2_ ( .D(U_dsdc_N4338), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__2_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__1_ ( .D(U_dsdc_N4337), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__1_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_0__0_ ( .D(U_dsdc_N4336), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_0__0_) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_0__2_ ( .D(U_dsdc_N4334), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_0__2_) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_0__1_ ( .D(U_dsdc_N4333), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_0__1_), .QN(U_dsdc_n402) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_0__0_ ( .D(U_dsdc_N4332), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_0__0_), .QN(U_dsdc_n192) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_0__3_ ( .D(U_dsdc_N4335), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_0__3_), .QN(U_dsdc_n441) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_0__2_ ( .D(U_dsdc_N4321), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_0__2_) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_0__1_ ( .D(U_dsdc_N4320), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_0__1_), .QN(U_dsdc_n424) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_0__0_ ( .D(U_dsdc_N4319), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_0__0_), .QN(U_dsdc_n189) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_0__3_ ( .D(U_dsdc_N4322), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_0__3_), .QN(U_dsdc_n363) );
  DFFS_X2 U_dsdc_r_bm_open_bank_reg_0_ ( .D(n83), .CK(hclk), .SN(hresetn), .Q(
        U_dsdc_n168), .QN(U_dsdc_r_bm_open_bank[0]) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__15_ ( .D(U_dsdc_N4398), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__15_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__14_ ( .D(U_dsdc_N4397), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__14_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__13_ ( .D(U_dsdc_N4396), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__13_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__6_ ( .D(U_dsdc_N4389), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__6_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__5_ ( .D(U_dsdc_N4388), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__5_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__4_ ( .D(U_dsdc_N4387), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__4_), .QN(U_dsdc_n339) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__3_ ( .D(U_dsdc_N4386), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__3_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__2_ ( .D(U_dsdc_N4385), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__2_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__1_ ( .D(U_dsdc_N4384), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__1_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_1__0_ ( .D(U_dsdc_N4383), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_1__0_) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_1__2_ ( .D(U_dsdc_N4381), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_1__2_) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_1__1_ ( .D(U_dsdc_N4380), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_1__1_), .QN(U_dsdc_n419) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_1__0_ ( .D(U_dsdc_N4379), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_1__0_), .QN(U_dsdc_n193) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_1__3_ ( .D(U_dsdc_N4382), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_1__3_), .QN(U_dsdc_n438) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_1__2_ ( .D(U_dsdc_N4368), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_1__2_) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_1__1_ ( .D(U_dsdc_N4367), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_1__1_), .QN(U_dsdc_n420) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_1__0_ ( .D(U_dsdc_N4366), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_1__0_), .QN(U_dsdc_n186) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_1__3_ ( .D(U_dsdc_N4369), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_1__3_), .QN(U_dsdc_n364) );
  DFFS_X2 U_dsdc_r_bm_open_bank_reg_1_ ( .D(U_dsdc_n307), .CK(hclk), .SN(
        hresetn), .Q(U_dsdc_n356), .QN(U_dsdc_r_bm_open_bank[1]) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__15_ ( .D(U_dsdc_N4445), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__15_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__14_ ( .D(U_dsdc_N4444), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__14_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__13_ ( .D(U_dsdc_N4443), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__13_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__6_ ( .D(U_dsdc_N4436), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__6_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__5_ ( .D(U_dsdc_N4435), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__5_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__4_ ( .D(U_dsdc_N4434), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__4_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__3_ ( .D(U_dsdc_N4433), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__3_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__2_ ( .D(U_dsdc_N4432), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__2_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__1_ ( .D(U_dsdc_N4431), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__1_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_2__0_ ( .D(U_dsdc_N4430), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_2__0_) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_2__2_ ( .D(U_dsdc_N4428), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_2__2_) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_2__1_ ( .D(U_dsdc_N4427), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_2__1_), .QN(U_dsdc_n401) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_2__0_ ( .D(U_dsdc_N4426), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_2__0_), .QN(U_dsdc_n191) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_2__3_ ( .D(U_dsdc_N4429), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_2__3_), .QN(U_dsdc_n439) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_2__2_ ( .D(U_dsdc_N4415), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_2__2_) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_2__1_ ( .D(U_dsdc_N4414), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_2__1_), .QN(U_dsdc_n422) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_2__0_ ( .D(U_dsdc_N4413), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_2__0_), .QN(U_dsdc_n188) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_2__3_ ( .D(U_dsdc_N4416), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_2__3_), .QN(U_dsdc_n365) );
  DFFS_X2 U_dsdc_r_bm_open_bank_reg_2_ ( .D(U_dsdc_n310), .CK(hclk), .SN(
        hresetn), .Q(U_dsdc_n164) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__15_ ( .D(U_dsdc_N4492), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__15_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__14_ ( .D(U_dsdc_N4491), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__14_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__13_ ( .D(U_dsdc_N4490), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__13_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__6_ ( .D(U_dsdc_N4483), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__6_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__5_ ( .D(U_dsdc_N4482), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__5_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__4_ ( .D(U_dsdc_N4481), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__4_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__3_ ( .D(U_dsdc_N4480), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__3_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__2_ ( .D(U_dsdc_N4479), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__2_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__1_ ( .D(U_dsdc_N4478), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__1_) );
  DFFR_X1 U_dsdc_bm_row_addr_reg_3__0_ ( .D(U_dsdc_N4477), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_row_addr_3__0_) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_3__2_ ( .D(U_dsdc_N4475), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_3__2_) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_3__1_ ( .D(U_dsdc_N4474), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_3__1_), .QN(U_dsdc_n400) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_3__0_ ( .D(U_dsdc_N4473), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_3__0_), .QN(U_dsdc_n190) );
  DFFR_X1 U_dsdc_bm_rc_cnt_reg_3__3_ ( .D(U_dsdc_N4476), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_rc_cnt_3__3_), .QN(U_dsdc_n442) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_3__2_ ( .D(U_dsdc_N4462), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_3__2_) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_3__1_ ( .D(U_dsdc_N4461), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_3__1_), .QN(U_dsdc_n421) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_3__0_ ( .D(U_dsdc_N4460), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_3__0_), .QN(U_dsdc_n187) );
  DFFR_X1 U_dsdc_bm_ras_cnt_reg_3__3_ ( .D(U_dsdc_N4463), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_ras_cnt_3__3_), .QN(U_dsdc_n382) );
  DFFS_X2 U_dsdc_r_bm_open_bank_reg_3_ ( .D(U_dsdc_n313), .CK(hclk), .SN(
        hresetn), .Q(U_dsdc_n185), .QN(U_dsdc_r_bm_open_bank[3]) );
  DFFR_X1 U_dsdc_rcar_cnt2_reg_2_ ( .D(U_dsdc_rcar_cnt2_nxt[2]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_rcar_cnt2_2_) );
  DFFR_X1 U_dsdc_rcar_cnt2_reg_1_ ( .D(U_dsdc_rcar_cnt2_nxt[1]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_rcar_cnt2_1_) );
  DFFR_X1 U_dsdc_rcar_cnt2_reg_0_ ( .D(U_dsdc_rcar_cnt2_nxt[0]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_rcar_cnt2_0_) );
  DFFR_X1 U_dsdc_wtr_cnt_reg_2_ ( .D(U_dsdc_wtr_cnt_nxt[2]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_wtr_cnt_2_) );
  DFFR_X1 U_dsdc_wtr_cnt_reg_0_ ( .D(U_dsdc_wtr_cnt_nxt[0]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_wtr_cnt_0_), .QN(U_dsdc_n398) );
  DFFR_X1 U_dsdc_r_data_mask_reg_0_ ( .D(U_dsdc_n249), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_data_mask[0]), .QN(U_dsdc_n469) );
  DFFR_X1 U_dsdc_r_data_mask_reg_1_ ( .D(U_dsdc_n250), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_data_mask[1]), .QN(U_dsdc_n470) );
  DFFR_X1 U_dsdc_r_data_mask_reg_2_ ( .D(U_dsdc_n251), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_data_mask[2]), .QN(U_dsdc_n471) );
  DFFR_X1 U_dsdc_r_data_mask_reg_3_ ( .D(U_dsdc_n252), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_data_mask[3]), .QN(U_dsdc_n472) );
  DFFR_X1 U_dsdc_r_bank_addr_reg_0_ ( .D(U_dsdc_n253), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_bank_addr_0_) );
  DFFR_X1 U_dsdc_r_bank_addr_reg_1_ ( .D(U_dsdc_n254), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_bank_addr_1_) );
  DFFR_X1 U_dsdc_r_row_addr_reg_10_ ( .D(U_dsdc_n256), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_10_) );
  DFFR_X1 U_dsdc_r_row_addr_reg_12_ ( .D(U_dsdc_n258), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_12_) );
  DFFR_X1 U_dsdc_r_row_addr_reg_4_ ( .D(U_dsdc_n265), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_4_) );
  DFFR_X1 U_dsdc_r_row_addr_reg_5_ ( .D(U_dsdc_n266), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_5_) );
  DFFR_X1 U_dsdc_r_row_addr_reg_6_ ( .D(U_dsdc_n267), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_6_) );
  DFFR_X1 U_dsdc_r_row_addr_reg_8_ ( .D(U_dsdc_n269), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_row_addr_8_) );
  DFFR_X1 U_dsdc_cas_cnt_reg_5_ ( .D(U_dsdc_cas_cnt_nxt[5]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_cas_cnt_5_) );
  DFFR_X1 U_dsdc_cas_cnt_reg_4_ ( .D(U_dsdc_cas_cnt_nxt[4]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_cas_cnt_4_) );
  DFFR_X1 U_dsdc_cas_cnt_reg_3_ ( .D(U_dsdc_cas_cnt_nxt[3]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_cas_cnt_3_) );
  DFFR_X1 U_dsdc_cas_cnt_reg_2_ ( .D(U_dsdc_cas_cnt_nxt[2]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_cas_cnt_2_) );
  DFFR_X1 U_dsdc_cas_cnt_reg_1_ ( .D(U_dsdc_cas_cnt_nxt[1]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_cas_cnt_1_) );
  DFFR_X1 U_dsdc_r_burst_size_reg_1_ ( .D(U_dsdc_n272), .CK(hclk), .RN(hresetn), .Q(U_dsdc_r_burst_size_1_) );
  DFFR_X1 U_dsdc_r_burst_size_reg_2_ ( .D(U_dsdc_n273), .CK(hclk), .RN(hresetn), .Q(U_dsdc_r_burst_size_2_) );
  DFFR_X1 U_dsdc_r_close_bank_addr_reg_0_ ( .D(U_dsdc_close_bank_addr_0_), 
        .CK(hclk), .RN(hresetn), .Q(U_dsdc_r_close_bank_addr_0_), .QN(
        U_dsdc_n292) );
  DFFR_X1 U_dsdc_r_bm_close_bank_reg_1_ ( .D(U_dsdc_bm_close_bank_1_), .CK(
        hclk), .RN(hresetn), .Q(U_dsdc_r_bm_close_bank_1_) );
  DFFR_X1 U_dsdc_r_bm_close_bank_reg_0_ ( .D(U_dsdc_bm_close_bank_0_), .CK(
        hclk), .RN(hresetn), .Q(U_dsdc_r_bm_close_bank_0_) );
  DFFR_X1 U_dsdc_r_bm_close_bank_reg_3_ ( .D(U_dsdc_bm_close_bank_3_), .CK(
        hclk), .RN(hresetn), .Q(U_dsdc_r_bm_close_bank_3_) );
  DFFR_X1 U_dsdc_r_close_bank_addr_reg_1_ ( .D(U_dsdc_close_bank_addr_1_), 
        .CK(hclk), .RN(hresetn), .Q(U_dsdc_r_close_bank_addr_1_) );
  DFFR_X1 U_dsdc_auto_ref_en_reg ( .D(U_dsdc_auto_ref_en_nxt), .CK(hclk), .RN(
        hresetn), .Q(ctl_auto_ref_en), .QN(n94) );
  DFFR_X1 U_dsdc_s_cke_reg ( .D(U_dsdc_n278), .CK(hclk), .RN(hresetn), .Q(
        s_cke) );
  DFFR_X1 U_dsdc_init_cnt_reg_15_ ( .D(U_dsdc_n418), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_15_) );
  DFFR_X1 U_dsdc_init_cnt_reg_14_ ( .D(U_dsdc_n417), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_14_) );
  DFFR_X1 U_dsdc_init_cnt_reg_13_ ( .D(U_dsdc_n416), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_13_) );
  DFFR_X1 U_dsdc_init_cnt_reg_12_ ( .D(U_dsdc_n415), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_12_) );
  DFFR_X1 U_dsdc_init_cnt_reg_11_ ( .D(U_dsdc_n414), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_11_) );
  DFFR_X1 U_dsdc_init_cnt_reg_10_ ( .D(U_dsdc_n413), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_10_) );
  DFFR_X1 U_dsdc_init_cnt_reg_9_ ( .D(U_dsdc_n412), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_9_) );
  DFFR_X1 U_dsdc_init_cnt_reg_8_ ( .D(U_dsdc_n411), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_8_) );
  DFFR_X1 U_dsdc_init_cnt_reg_7_ ( .D(U_dsdc_n410), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_7_) );
  DFFR_X1 U_dsdc_init_cnt_reg_6_ ( .D(U_dsdc_n409), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_6_) );
  DFFR_X1 U_dsdc_init_cnt_reg_5_ ( .D(U_dsdc_n408), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_5_) );
  DFFR_X1 U_dsdc_init_cnt_reg_4_ ( .D(U_dsdc_n407), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_4_) );
  DFFR_X1 U_dsdc_init_cnt_reg_3_ ( .D(U_dsdc_n406), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_3_) );
  DFFR_X1 U_dsdc_init_cnt_reg_2_ ( .D(U_dsdc_n405), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_2_), .QN(U_dsdc_n468) );
  DFFR_X1 U_dsdc_init_cnt_reg_1_ ( .D(U_dsdc_n404), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_1_) );
  DFFR_X1 U_dsdc_init_cnt_reg_0_ ( .D(U_dsdc_n403), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_init_cnt_0_) );
  DFFR_X1 U_dsdc_row_cnt_reg_0_ ( .D(U_dsdc_n366), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_0_), .QN(U_dsdc_n462) );
  DFFR_X1 U_dsdc_row_cnt_reg_10_ ( .D(U_dsdc_n367), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_10_), .QN(U_dsdc_n208) );
  DFFR_X1 U_dsdc_row_cnt_reg_11_ ( .D(U_dsdc_n368), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_11_) );
  DFFR_X1 U_dsdc_row_cnt_reg_13_ ( .D(U_dsdc_n370), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_13_), .QN(U_dsdc_n197) );
  DFFR_X1 U_dsdc_row_cnt_reg_14_ ( .D(U_dsdc_n371), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_14_), .QN(U_dsdc_n202) );
  DFFR_X1 U_dsdc_row_cnt_reg_15_ ( .D(U_dsdc_n372), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_15_), .QN(U_dsdc_n426) );
  DFFR_X1 U_dsdc_row_cnt_reg_1_ ( .D(U_dsdc_n373), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_1_), .QN(U_dsdc_n465) );
  DFFR_X1 U_dsdc_row_cnt_reg_2_ ( .D(U_dsdc_n374), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_2_), .QN(U_dsdc_n204) );
  DFFR_X1 U_dsdc_row_cnt_reg_3_ ( .D(U_dsdc_n375), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_3_) );
  DFFR_X1 U_dsdc_row_cnt_reg_4_ ( .D(U_dsdc_n376), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_4_), .QN(U_dsdc_n207) );
  DFFR_X1 U_dsdc_row_cnt_reg_5_ ( .D(U_dsdc_n377), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_5_) );
  DFFR_X1 U_dsdc_row_cnt_reg_6_ ( .D(U_dsdc_n378), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_6_), .QN(U_dsdc_n206) );
  DFFR_X1 U_dsdc_row_cnt_reg_7_ ( .D(U_dsdc_n379), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_7_) );
  DFFR_X1 U_dsdc_row_cnt_reg_8_ ( .D(U_dsdc_n380), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_8_), .QN(U_dsdc_n205) );
  DFFR_X1 U_dsdc_row_cnt_reg_9_ ( .D(U_dsdc_n381), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_row_cnt_9_) );
  DFFR_X1 U_dsdc_rcar_cnt1_reg_3_ ( .D(U_dsdc_rcar_cnt1_nxt[3]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_rcar_cnt1_3_) );
  DFFR_X1 U_dsdc_rcar_cnt1_reg_2_ ( .D(U_dsdc_rcar_cnt1_nxt[2]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_rcar_cnt1_2_) );
  DFFR_X1 U_dsdc_rcar_cnt1_reg_1_ ( .D(U_dsdc_rcar_cnt1_nxt[1]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_rcar_cnt1_1_) );
  DFFR_X1 U_dsdc_rcar_cnt1_reg_0_ ( .D(U_dsdc_rcar_cnt1_nxt[0]), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_rcar_cnt1_0_) );
  DFFR_X1 U_dsdc_xsr_cnt_reg_0_ ( .D(U_dsdc_n386), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_xsr_cnt_0_) );
  DFFR_X1 U_dsdc_xsr_cnt_reg_1_ ( .D(U_dsdc_n387), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_xsr_cnt_1_) );
  DFFR_X1 U_dsdc_xsr_cnt_reg_2_ ( .D(U_dsdc_n388), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_xsr_cnt_2_) );
  DFFR_X1 U_dsdc_xsr_cnt_reg_3_ ( .D(U_dsdc_n389), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_xsr_cnt_3_) );
  DFFR_X1 U_dsdc_xsr_cnt_reg_4_ ( .D(U_dsdc_n390), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_xsr_cnt_4_) );
  DFFR_X1 U_dsdc_xsr_cnt_reg_5_ ( .D(U_dsdc_n391), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_xsr_cnt_5_) );
  DFFR_X1 U_dsdc_xsr_cnt_reg_7_ ( .D(U_dsdc_n393), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_xsr_cnt_7_) );
  DFFR_X1 U_dsdc_xsr_cnt_reg_8_ ( .D(U_dsdc_n394), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_xsr_cnt_8_) );
  DFFR_X1 U_dsdc_operation_cs_reg_2_ ( .D(U_dsdc_n2095), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_operation_cs_2_), .QN(U_dsdc_n341) );
  DFFR_X1 U_dsdc_operation_cs_reg_4_ ( .D(U_dsdc_n2093), .CK(hclk), .RN(
        hresetn), .QN(U_dsdc_n432) );
  DFFR_X1 U_dsdc_num_init_ref_cnt_reg_3_ ( .D(U_dsdc_n431), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_num_init_ref_cnt_3_) );
  DFFR_X1 U_dsdc_operation_cs_reg_0_ ( .D(U_dsdc_n2097), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_operation_cs_0_), .QN(U_dsdc_n344) );
  DFFR_X1 U_dsdc_operation_cs_reg_1_ ( .D(U_dsdc_n2096), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_operation_cs_1_), .QN(U_dsdc_n343) );
  DFFR_X1 U_dsdc_t_xp_cnt_reg_1_ ( .D(U_dsdc_N4229), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_t_xp_cnt_1_), .QN(U_dsdc_n474) );
  DFFR_X1 U_dsdc_t_xp_cnt_reg_0_ ( .D(U_dsdc_N4228), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_t_xp_cnt_0_), .QN(U_dsdc_n239) );
  DFFR_X1 U_dsdc_access_cs_reg_4_ ( .D(U_dsdc_n[2088]), .CK(hclk), .RN(hresetn), .Q(U_dsdc_access_cs_4_), .QN(U_dsdc_n167) );
  DFFR_X1 U_dsdc_wr_cnt_reg_2_ ( .D(U_dsdc_wr_cnt_nxt[2]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_wr_cnt_2_) );
  DFFR_X1 U_dsdc_wr_cnt_reg_1_ ( .D(U_dsdc_wr_cnt_nxt[1]), .CK(hclk), .RN(
        hresetn), .QN(U_dsdc_n195) );
  DFFR_X1 U_dsdc_wr_cnt_reg_0_ ( .D(U_dsdc_wr_cnt_nxt[0]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_wr_cnt_0_), .QN(U_dsdc_n397) );
  DFFR_X1 U_dsdc_access_cs_reg_3_ ( .D(U_dsdc_n[2089]), .CK(hclk), .RN(hresetn), .Q(U_dsdc_access_cs_3_), .QN(U_dsdc_n173) );
  DFFR_X1 U_dsdc_rp_cnt2_reg_2_ ( .D(U_dsdc_rp_cnt2_nxt[2]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_rp_cnt2_2_) );
  DFFR_X1 U_dsdc_rp_cnt2_reg_1_ ( .D(U_dsdc_rp_cnt2_nxt[1]), .CK(hclk), .RN(
        hresetn), .QN(U_dsdc_n309) );
  DFFS_X2 U_dsdc_r_rw_reg ( .D(U_dsdc_n279), .CK(hclk), .SN(hresetn), .Q(
        U_dsdc_r_rw), .QN(U_dsdc_n166) );
  DFFR_X1 U_dsdc_r_chip_slct_reg_0_ ( .D(U_dsdc_n280), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_r_chip_slct_0_), .QN(U_dsdc_n361) );
  DFFR_X1 U_dsdc_access_cs_reg_0_ ( .D(U_dsdc_n[2092]), .CK(hclk), .RN(hresetn), .Q(U_dsdc_access_cs_0_), .QN(U_dsdc_n170) );
  DFFR_X1 U_dsdc_term_cnt_reg_4_ ( .D(U_dsdc_term_cnt_nxt[4]), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_term_cnt_4_), .QN(U_dsdc_n457) );
  DFFR_X1 U_dsdc_data_cnt_reg_0_ ( .D(U_dsdc_n286), .CK(hclk), .RN(hresetn), 
        .Q(U_dsdc_data_cnt_0_), .QN(U_dsdc_n347) );
  DFFR_X1 U_dsdc_access_cs_reg_1_ ( .D(U_dsdc_n[2091]), .CK(hclk), .RN(hresetn), .Q(U_dsdc_access_cs_1_), .QN(U_dsdc_n298) );
  DFFR_X1 U_dsdc_bm_bank_status_reg_2_ ( .D(U_dsdc_N4449), .CK(hclk), .RN(
        hresetn), .Q(U_dsdc_bm_bank_status_2_), .QN(U_dsdc_n395) );
  DFFR_X1 U_dsdc_r_bm_close_bank_reg_2_ ( .D(U_dsdc_bm_close_bank_2_), .CK(
        hclk), .RN(hresetn), .Q(U_dsdc_r_bm_close_bank_2_) );
  DFFR_X1 U_dsdc_r_cas_latency_reg_1_ ( .D(U_dsdc_cas_latency_1_), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_r_cas_latency_1_) );
  DFFR_X1 U_dsdc_r_cas_latency_reg_2_ ( .D(U_dsdc_cas_latency_2_), .CK(hclk), 
        .RN(hresetn), .Q(U_dsdc_r_cas_latency_2_) );
  DFFS_X2 U_dsdc_r_cas_latency_reg_3_ ( .D(U_dsdc_n554), .CK(hclk), .SN(
        hresetn), .QN(U_dsdc_r_cas_latency_3_) );
  XNOR2_X1 U_ddrwr_U59 ( .A(hclk_2x), .B(scan_mode), .ZN(
        U_ddrwr_hclk_2x_scan_clk) );
  NOR2_X2 U_ddrwr_U58 ( .A1(U_ddrwr_n27), .A2(cr_s_data_width_early_0_), .ZN(
        U_ddrwr_n52) );
  OAI221_X2 U_ddrwr_U56 ( .B1(s_cas_latency[1]), .B2(pre_rd_dqs_mask), .C1(n93), .C2(U_ddrwr_rd_dqs_mask_d_3_), .A(s_cas_latency[0]), .ZN(U_ddrwr_n32) );
  OAI221_X2 U_ddrwr_U55 ( .B1(s_cas_latency[1]), .B2(U_ddrwr_rd_dqs_mask_d_3_), 
        .C1(n93), .C2(U_ddrwr_rd_dqs_mask_d_1_), .A(n90), .ZN(U_ddrwr_n31) );
  AOI22_X2 U_ddrwr_U54 ( .A1(s_cas_latency[1]), .A2(U_ddrwr_rd_dqs_mask_d_2_), 
        .B1(U_ddrwr_rd_dqs_mask_d_5_), .B2(n93), .ZN(U_ddrwr_n28) );
  OAI221_X2 U_ddrwr_U53 ( .B1(s_cas_latency[1]), .B2(U_ddrwr_rd_dqs_mask_d_0_), 
        .C1(n93), .C2(U_ddrwr_rd_dqs_mask_d_4_), .A(s_cas_latency[0]), .ZN(
        U_ddrwr_n26) );
  OAI21_X2 U_ddrwr_U52 ( .B1(s_cas_latency[0]), .B2(U_ddrwr_n28), .A(
        U_ddrwr_n26), .ZN(U_ddrwr_n29) );
  NAND2_X2 U_ddrwr_U51 ( .A1(U_ddrwr_n29), .A2(s_cas_latency[2]), .ZN(
        U_ddrwr_n30) );
  OAI21_X2 U_ddrwr_U48 ( .B1(n88), .B2(U_ddrwr_r_pre_dqs_hclk_2x), .A(
        U_ddrwr_r_dqs), .ZN(U_ddrwr_n33) );
  NOR2_X2 U_ddrwr_U47 ( .A1(pre_amble), .A2(U_ddrwr_n33), .ZN(U_ddrwr_i_dqs_1_) );
  NAND2_X2 U_ddrwr_U46 ( .A1(U_ddrwr_r_dqs), .A2(n88), .ZN(U_ddrwr_N44) );
  AOI222_X1 U_ddrwr_U43 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_7_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_23_), .C1(U_ddrwr_n52), .C2(
        U_ddrwr_r_wr_data_15_), .ZN(U_ddrwr_n45) );
  AOI222_X1 U_ddrwr_U42 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_3_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_19_), .C1(U_ddrwr_n52), .C2(
        U_ddrwr_r_wr_data_11_), .ZN(U_ddrwr_n49) );
  AOI222_X1 U_ddrwr_U41 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_2_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_18_), .C1(U_ddrwr_n52), .C2(
        U_ddrwr_r_wr_data_10_), .ZN(U_ddrwr_n50) );
  AOI222_X1 U_ddrwr_U40 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_1_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_17_), .C1(U_ddrwr_n52), .C2(
        U_ddrwr_r_wr_data_9_), .ZN(U_ddrwr_n51) );
  AOI222_X1 U_ddrwr_U39 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_5_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_21_), .C1(U_ddrwr_n52), .C2(
        U_ddrwr_r_wr_data_13_), .ZN(U_ddrwr_n47) );
  AOI222_X1 U_ddrwr_U38 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_6_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_22_), .C1(U_ddrwr_n52), .C2(
        U_ddrwr_r_wr_data_14_), .ZN(U_ddrwr_n46) );
  AOI222_X1 U_ddrwr_U37 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_pre_dqm_0_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_pre_dqm_2_), .C1(U_ddrwr_n52), .C2(
        U_ddrwr_r_pre_dqm_1_), .ZN(U_ddrwr_n36) );
  AOI222_X1 U_ddrwr_U36 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_0_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_16_), .C1(U_ddrwr_n52), .C2(
        U_ddrwr_r_wr_data_8_), .ZN(U_ddrwr_n54) );
  AOI222_X1 U_ddrwr_U35 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_4_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_20_), .C1(U_ddrwr_n52), .C2(
        U_ddrwr_r_wr_data_12_), .ZN(U_ddrwr_n48) );
  OAI221_X1 U_ddrwr_U34 ( .B1(s_cas_latency[2]), .B2(U_ddrwr_n32), .C1(
        s_cas_latency[2]), .C2(U_ddrwr_n31), .A(U_ddrwr_n30), .ZN(U_ddrwr_N41)
         );
  NOR2_X2 U_ddrwr_U33 ( .A1(U_ddrwr_n27), .A2(n85), .ZN(U_ddrwr_n53) );
  AOI22_X1 U_ddrwr_U29 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_11_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_27_), .ZN(U_ddrwr_n41) );
  AOI22_X1 U_ddrwr_U28 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_10_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_26_), .ZN(U_ddrwr_n42) );
  AOI22_X1 U_ddrwr_U27 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_12_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_28_), .ZN(U_ddrwr_n40) );
  AOI22_X1 U_ddrwr_U26 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_9_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_25_), .ZN(U_ddrwr_n43) );
  AOI22_X1 U_ddrwr_U25 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_13_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_29_), .ZN(U_ddrwr_n39) );
  AOI22_X1 U_ddrwr_U24 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_14_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_30_), .ZN(U_ddrwr_n38) );
  AOI22_X1 U_ddrwr_U23 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_15_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_31_), .ZN(U_ddrwr_n37) );
  AOI22_X1 U_ddrwr_U22 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_wr_data_8_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_wr_data_24_), .ZN(U_ddrwr_n44) );
  AOI22_X1 U_ddrwr_U21 ( .A1(U_ddrwr_n27), .A2(U_ddrwr_r_pre_dqm_1_), .B1(
        U_ddrwr_n53), .B2(U_ddrwr_r_pre_dqm_3_), .ZN(U_ddrwr_n35) );
  INV_X2 U_ddrwr_U20 ( .A(U_ddrwr_n50), .ZN(U_ddrwr_n3) );
  INV_X2 U_ddrwr_U19 ( .A(U_ddrwr_n54), .ZN(U_ddrwr_n1) );
  INV_X2 U_ddrwr_U18 ( .A(U_ddrwr_n51), .ZN(U_ddrwr_n2) );
  INV_X2 U_ddrwr_U17 ( .A(U_ddrwr_n49), .ZN(U_ddrwr_n4) );
  INV_X2 U_ddrwr_U16 ( .A(U_ddrwr_n48), .ZN(U_ddrwr_n5) );
  INV_X2 U_ddrwr_U15 ( .A(U_ddrwr_n35), .ZN(U_ddrwr_n18) );
  INV_X2 U_ddrwr_U14 ( .A(U_ddrwr_n47), .ZN(U_ddrwr_n6) );
  INV_X2 U_ddrwr_U13 ( .A(U_ddrwr_n46), .ZN(U_ddrwr_n7) );
  INV_X2 U_ddrwr_U12 ( .A(U_ddrwr_n40), .ZN(U_ddrwr_n13) );
  INV_X2 U_ddrwr_U11 ( .A(U_ddrwr_n36), .ZN(U_ddrwr_n17) );
  INV_X2 U_ddrwr_U10 ( .A(U_ddrwr_n45), .ZN(U_ddrwr_n8) );
  INV_X2 U_ddrwr_U9 ( .A(U_ddrwr_n37), .ZN(U_ddrwr_n16) );
  INV_X2 U_ddrwr_U8 ( .A(U_ddrwr_n44), .ZN(U_ddrwr_n9) );
  INV_X2 U_ddrwr_U7 ( .A(U_ddrwr_n38), .ZN(U_ddrwr_n15) );
  INV_X2 U_ddrwr_U6 ( .A(U_ddrwr_n43), .ZN(U_ddrwr_n10) );
  INV_X2 U_ddrwr_U5 ( .A(U_ddrwr_n42), .ZN(U_ddrwr_n11) );
  INV_X2 U_ddrwr_U4 ( .A(U_ddrwr_n39), .ZN(U_ddrwr_n14) );
  INV_X2 U_ddrwr_U3 ( .A(U_ddrwr_n41), .ZN(U_ddrwr_n12) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_7_ ( .D(hiu_wr_data[7]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_7_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_0_ ( .D(hiu_wr_data[0]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_0_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_1_ ( .D(hiu_wr_data[1]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_1_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_27_ ( .D(hiu_wr_data[27]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_27_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_28_ ( .D(hiu_wr_data[28]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_28_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_29_ ( .D(hiu_wr_data[29]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_29_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_30_ ( .D(hiu_wr_data[30]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_30_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_31_ ( .D(hiu_wr_data[31]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_31_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_26_ ( .D(hiu_wr_data[26]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_26_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_24_ ( .D(hiu_wr_data[24]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_24_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_25_ ( .D(hiu_wr_data[25]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_25_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_17_ ( .D(hiu_wr_data[17]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_17_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_18_ ( .D(hiu_wr_data[18]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_18_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_19_ ( .D(hiu_wr_data[19]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_19_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_20_ ( .D(hiu_wr_data[20]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_20_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_21_ ( .D(hiu_wr_data[21]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_21_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_22_ ( .D(hiu_wr_data[22]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_22_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_16_ ( .D(hiu_wr_data[16]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_16_) );
  DFFR_X2 U_ddrwr_r_wr_data_reg_23_ ( .D(hiu_wr_data[23]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_23_) );
  DFFR_X2 U_ddrwr_r_pre_dqm_reg_0_ ( .D(pre_dqm[0]), .CK(hclk), .RN(hresetn), 
        .Q(U_ddrwr_r_pre_dqm_0_) );
  DFFR_X2 U_ddrwr_r_pre_dqm_reg_1_ ( .D(pre_dqm[1]), .CK(hclk), .RN(hresetn), 
        .Q(U_ddrwr_r_pre_dqm_1_) );
  DFFR_X2 U_ddrwr_r_pre_dqm_reg_2_ ( .D(pre_dqm[2]), .CK(hclk), .RN(hresetn), 
        .Q(U_ddrwr_r_pre_dqm_2_) );
  DFFR_X2 U_ddrwr_r_pre_dqm_reg_3_ ( .D(pre_dqm[3]), .CK(hclk), .RN(hresetn), 
        .Q(U_ddrwr_r_pre_dqm_3_) );
  MUX2_X2 U_ddrwr_U49 ( .A(hclk), .B(U_ddrwr_r_dqs), .S(scan_mode), .Z(
        U_ddrwr_n27) );
  DFFR_X1 U_ddrwr_s_dqm_reg_0_ ( .D(U_ddrwr_ddr_dqm[0]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_dqm[0]) );
  DFFR_X1 U_ddrwr_s_dqm_reg_1_ ( .D(U_ddrwr_ddr_dqm[1]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_dqm[1]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_0_ ( .D(U_ddrwr_ddr_wr_data[0]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[0]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_1_ ( .D(U_ddrwr_ddr_wr_data[1]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[1]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_2_ ( .D(U_ddrwr_ddr_wr_data[2]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[2]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_3_ ( .D(U_ddrwr_ddr_wr_data[3]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[3]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_4_ ( .D(U_ddrwr_ddr_wr_data[4]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[4]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_5_ ( .D(U_ddrwr_ddr_wr_data[5]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[5]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_6_ ( .D(U_ddrwr_ddr_wr_data[6]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[6]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_7_ ( .D(U_ddrwr_ddr_wr_data[7]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[7]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_8_ ( .D(U_ddrwr_ddr_wr_data[8]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[8]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_9_ ( .D(U_ddrwr_ddr_wr_data[9]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[9]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_10_ ( .D(U_ddrwr_ddr_wr_data[10]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[10]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_11_ ( .D(U_ddrwr_ddr_wr_data[11]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[11]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_12_ ( .D(U_ddrwr_ddr_wr_data[12]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[12]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_13_ ( .D(U_ddrwr_ddr_wr_data[13]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[13]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_14_ ( .D(U_ddrwr_ddr_wr_data[14]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[14]) );
  DFFR_X1 U_ddrwr_s_wr_data_reg_15_ ( .D(U_ddrwr_ddr_wr_data[15]), .CK(
        U_ddrwr_hclk_2x_scan_clk), .RN(hresetn), .Q(s_wr_data[15]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_0_ ( .D(U_ddrwr_n1), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[0]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_1_ ( .D(U_ddrwr_n2), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[1]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_2_ ( .D(U_ddrwr_n3), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[2]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_3_ ( .D(U_ddrwr_n4), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[3]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_4_ ( .D(U_ddrwr_n5), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[4]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_5_ ( .D(U_ddrwr_n6), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[5]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_6_ ( .D(U_ddrwr_n7), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[6]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_7_ ( .D(U_ddrwr_n8), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[7]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_8_ ( .D(U_ddrwr_n9), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[8]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_9_ ( .D(U_ddrwr_n10), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[9]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_10_ ( .D(U_ddrwr_n11), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[10]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_11_ ( .D(U_ddrwr_n12), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[11]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_12_ ( .D(U_ddrwr_n13), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[12]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_13_ ( .D(U_ddrwr_n14), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[13]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_14_ ( .D(U_ddrwr_n15), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[14]) );
  DFFR_X1 U_ddrwr_ddr_wr_data_reg_15_ ( .D(U_ddrwr_n16), .CK(hclk_2x), .RN(
        hresetn), .Q(U_ddrwr_ddr_wr_data[15]) );
  DFFR_X1 U_ddrwr_ddr_dqm_reg_0_ ( .D(U_ddrwr_n17), .CK(hclk_2x), .RN(hresetn), 
        .Q(U_ddrwr_ddr_dqm[0]) );
  DFFR_X1 U_ddrwr_ddr_dqm_reg_1_ ( .D(U_ddrwr_n18), .CK(hclk_2x), .RN(hresetn), 
        .Q(U_ddrwr_ddr_dqm[1]) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_2_ ( .D(hiu_wr_data[2]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_2_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_3_ ( .D(hiu_wr_data[3]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_3_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_4_ ( .D(hiu_wr_data[4]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_4_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_5_ ( .D(hiu_wr_data[5]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_5_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_6_ ( .D(hiu_wr_data[6]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_6_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_8_ ( .D(hiu_wr_data[8]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_8_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_9_ ( .D(hiu_wr_data[9]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_9_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_10_ ( .D(hiu_wr_data[10]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_10_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_11_ ( .D(hiu_wr_data[11]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_11_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_12_ ( .D(hiu_wr_data[12]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_12_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_13_ ( .D(hiu_wr_data[13]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_13_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_14_ ( .D(hiu_wr_data[14]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_14_) );
  DFFR_X1 U_ddrwr_r_wr_data_reg_15_ ( .D(hiu_wr_data[15]), .CK(hclk), .RN(
        hresetn), .Q(U_ddrwr_r_wr_data_15_) );
  DFFS_X2 U_ddrwr_s_dqs_reg_0_ ( .D(U_ddrwr_i2_dqs[0]), .CK(hclk_2x), .SN(
        hresetn), .Q(s_dqs[0]) );
  DFFS_X2 U_ddrwr_s_dqs_reg_1_ ( .D(U_ddrwr_i2_dqs[1]), .CK(hclk_2x), .SN(
        hresetn), .Q(s_dqs[1]) );
  DFFS_X2 U_ddrwr_i2_dqs_reg_0_ ( .D(U_ddrwr_i_dqs_1_), .CK(hclk_2x), .SN(
        hresetn), .Q(U_ddrwr_i2_dqs[0]) );
  DFFS_X2 U_ddrwr_i2_dqs_reg_1_ ( .D(U_ddrwr_i_dqs_1_), .CK(hclk_2x), .SN(
        hresetn), .Q(U_ddrwr_i2_dqs[1]) );
  DFFS_X2 U_ddrwr_r_dqs_reg ( .D(U_ddrwr_N44), .CK(hclk_2x), .SN(hresetn), .Q(
        U_ddrwr_r_dqs) );
  DFFR_X1 U_ddrwr_r_pre_dqs_hclk_2x_reg ( .D(n88), .CK(hclk_2x), .RN(hresetn), 
        .QN(U_ddrwr_r_pre_dqs_hclk_2x) );
  DFFR_X1 U_ddrwr_s_rd_dqs_mask_reg ( .D(U_ddrwr_N41), .CK(hclk_2x), .RN(
        hresetn), .Q(s_rd_dqs_mask) );
  DFFR_X1 U_ddrwr_rd_dqs_mask_d_reg_5_ ( .D(U_ddrwr_rd_dqs_mask_d_4_), .CK(
        hclk_2x), .RN(hresetn), .Q(U_ddrwr_rd_dqs_mask_d_5_) );
  DFFR_X1 U_ddrwr_rd_dqs_mask_d_reg_4_ ( .D(U_ddrwr_rd_dqs_mask_d_3_), .CK(
        hclk_2x), .RN(hresetn), .Q(U_ddrwr_rd_dqs_mask_d_4_) );
  DFFR_X1 U_ddrwr_rd_dqs_mask_d_reg_3_ ( .D(U_ddrwr_rd_dqs_mask_d_2_), .CK(
        hclk_2x), .RN(hresetn), .Q(U_ddrwr_rd_dqs_mask_d_3_) );
  DFFR_X1 U_ddrwr_rd_dqs_mask_d_reg_2_ ( .D(U_ddrwr_rd_dqs_mask_d_1_), .CK(
        hclk_2x), .RN(hresetn), .Q(U_ddrwr_rd_dqs_mask_d_2_) );
  DFFR_X1 U_ddrwr_rd_dqs_mask_d_reg_1_ ( .D(U_ddrwr_rd_dqs_mask_d_0_), .CK(
        hclk_2x), .RN(hresetn), .Q(U_ddrwr_rd_dqs_mask_d_1_) );
  DFFR_X1 U_ddrwr_rd_dqs_mask_d_reg_0_ ( .D(pre_rd_dqs_mask), .CK(hclk_2x), 
        .RN(hresetn), .Q(U_ddrwr_rd_dqs_mask_d_0_) );
  OAI22_X1 U_cr_U595 ( .A1(n27), .A2(U_cr_n531), .B1(U_cr_n519), .B2(U_cr_n17), 
        .ZN(U_cr_n507) );
  NAND2_X1 U_cr_U594 ( .A1(U_cr_n17), .A2(hiu_rw), .ZN(U_cr_n504) );
  AOI22_X1 U_cr_U593 ( .A1(U_cr_n422), .A2(s_read_pipe[0]), .B1(U_cr_n407), 
        .B2(cr_row_addr_width[1]), .ZN(U_cr_n387) );
  INV_X4 U_cr_U591 ( .A(U_cr_n487), .ZN(U_cr_n204) );
  INV_X4 U_cr_U590 ( .A(U_cr_n492), .ZN(U_cr_n203) );
  NAND3_X2 U_cr_U589 ( .A1(U_cr_n180), .A2(U_cr_n185), .A3(U_cr_n179), .ZN(
        U_cr_n182) );
  NOR2_X2 U_cr_U588 ( .A1(hiu_haddr[2]), .A2(U_cr_n308), .ZN(U_cr_n424) );
  NAND3_X2 U_cr_U587 ( .A1(U_cr_n227), .A2(U_cr_n320), .A3(U_cr_n283), .ZN(
        U_cr_n416) );
  OR2_X4 U_cr_U586 ( .A1(hiu_haddr[2]), .A2(U_cr_n263), .ZN(U_cr_n25) );
  NAND3_X2 U_cr_U585 ( .A1(U_cr_n283), .A2(hiu_haddr[2]), .A3(U_cr_n227), .ZN(
        U_cr_n391) );
  INV_X4 U_cr_U584 ( .A(U_cr_n391), .ZN(U_cr_n430) );
  AOI221_X2 U_cr_U583 ( .B1(ad_cr_data_mask[0]), .B2(big_endian), .C1(
        ad_cr_data_mask[3]), .C2(U_addrdec_n40), .A(U_cr_n237), .ZN(U_cr_n239)
         );
  NOR2_X2 U_cr_U582 ( .A1(big_endian), .A2(U_cr_n241), .ZN(U_cr_n258) );
  NOR2_X2 U_cr_U581 ( .A1(U_cr_n242), .A2(U_cr_n241), .ZN(U_cr_n259) );
  NOR2_X2 U_cr_U580 ( .A1(U_cr_n526), .A2(U_cr_n416), .ZN(U_cr_n215) );
  INV_X4 U_cr_U579 ( .A(U_cr_n230), .ZN(U_cr_n229) );
  INV_X4 U_cr_U578 ( .A(U_cr_n313), .ZN(U_cr_n312) );
  INV_X4 U_cr_U577 ( .A(U_cr_n536), .ZN(U_cr_n538) );
  INV_X4 U_cr_U576 ( .A(U_cr_n305), .ZN(U_cr_n304) );
  INV_X4 U_cr_U575 ( .A(U_cr_n289), .ZN(U_cr_n288) );
  NAND3_X1 U_cr_U574 ( .A1(U_cr_n194), .A2(U_cr_n17), .A3(U_cr_n23), .ZN(
        U_cr_n174) );
  NOR2_X2 U_cr_U573 ( .A1(U_cr_n182), .A2(U_addrdec_n40), .ZN(U_cr_n499) );
  INV_X4 U_cr_U572 ( .A(U_cr_n268), .ZN(U_cr_n267) );
  AND2_X4 U_cr_U571 ( .A1(n27), .A2(U_cr_n223), .ZN(U_cr_n511) );
  NOR2_X2 U_cr_U570 ( .A1(U_cr_n544), .A2(U_cr_n416), .ZN(U_cr_n221) );
  NOR2_X2 U_cr_U569 ( .A1(U_cr_n544), .A2(U_cr_n358), .ZN(U_cr_n307) );
  NOR2_X2 U_cr_U568 ( .A1(U_cr_n544), .A2(U_cr_n334), .ZN(U_cr_n542) );
  INV_X4 U_cr_U567 ( .A(U_cr_n294), .ZN(U_cr_n292) );
  INV_X4 U_cr_U566 ( .A(U_cr_n270), .ZN(U_cr_n269) );
  NAND3_X1 U_cr_U565 ( .A1(hiu_reg_req), .A2(U_cr_n194), .A3(n27), .ZN(
        U_cr_n195) );
  XNOR2_X2 U_cr_U564 ( .A(U_cr_sctlr_16_), .B(U_cr_n210), .ZN(U_cr_N574) );
  XNOR2_X2 U_cr_U563 ( .A(U_cr_stmg0r_26), .B(U_cr_n282), .ZN(U_cr_N577) );
  INV_X4 U_cr_U562 ( .A(U_cr_n236), .ZN(U_cr_n205) );
  INV_X4 U_cr_U561 ( .A(U_cr_n422), .ZN(U_cr_n396) );
  AOI222_X2 U_cr_U560 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[3]), .B1(U_cr_n168), .B2(hiu_wr_data[27]), .C1(hiu_wr_data[11]), .C2(U_cr_n319), .ZN(U_cr_n531)
         );
  INV_X4 U_cr_U559 ( .A(U_cr_n424), .ZN(U_cr_n334) );
  NAND3_X2 U_cr_U558 ( .A1(U_cr_n284), .A2(hiu_addr[4]), .A3(U_cr_n283), .ZN(
        U_cr_n315) );
  INV_X4 U_cr_U557 ( .A(U_cr_n423), .ZN(U_cr_n358) );
  NAND2_X2 U_cr_U556 ( .A1(U_cr_n182), .A2(big_endian), .ZN(U_cr_n487) );
  NAND2_X2 U_cr_U555 ( .A1(U_cr_n182), .A2(U_addrdec_n40), .ZN(U_cr_n492) );
  AOI221_X2 U_cr_U554 ( .B1(U_addrdec_n40), .B2(ad_cr_data_mask[2]), .C1(
        big_endian), .C2(ad_cr_data_mask[1]), .A(U_cr_n205), .ZN(U_cr_n223) );
  INV_X4 U_cr_U553 ( .A(U_cr_n232), .ZN(U_cr_n231) );
  AOI21_X2 U_cr_U552 ( .B1(hiu_rw), .B2(U_cr_cr_cs_1_), .A(U_cr_cr_cs_0_), 
        .ZN(U_cr_n187) );
  INV_X4 U_cr_U551 ( .A(U_cr_n190), .ZN(U_cr_n199) );
  OAI211_X2 U_cr_U550 ( .C1(U_cr_n187), .C2(U_cr_n24), .A(U_cr_n186), .B(
        U_cr_n199), .ZN(cr_pop_n) );
  AOI222_X2 U_cr_U548 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[8]), .B1(U_cr_n168), .B2(hiu_wr_data[16]), .C1(hiu_wr_data[0]), .C2(U_cr_n319), .ZN(U_cr_n548) );
  NOR3_X2 U_cr_U547 ( .A1(hiu_burst_size[3]), .A2(hiu_burst_size[5]), .A3(
        hiu_burst_size[0]), .ZN(U_cr_n212) );
  NAND3_X2 U_cr_U546 ( .A1(hiu_burst_size[1]), .A2(U_cr_n212), .A3(U_cr_n211), 
        .ZN(U_cr_n550) );
  NAND2_X2 U_cr_U545 ( .A1(hiu_haddr[1]), .A2(U_cr_n550), .ZN(U_cr_n318) );
  NOR4_X2 U_cr_U544 ( .A1(hiu_addr[5]), .A2(hiu_addr[7]), .A3(hiu_addr[6]), 
        .A4(hiu_addr[4]), .ZN(U_cr_n227) );
  NAND2_X2 U_cr_U543 ( .A1(U_cr_n202), .A2(U_cr_n200), .ZN(U_cr_n236) );
  NAND2_X2 U_cr_U542 ( .A1(U_cr_n238), .A2(U_cr_n239), .ZN(U_cr_n262) );
  NAND2_X2 U_cr_U541 ( .A1(U_cr_n239), .A2(n27), .ZN(U_cr_n241) );
  NAND2_X2 U_cr_U540 ( .A1(U_cr_n240), .A2(U_cr_n239), .ZN(U_cr_n257) );
  AOI22_X2 U_cr_U539 ( .A1(hiu_wr_data[24]), .A2(U_cr_n258), .B1(cr_t_rc[2]), 
        .B2(U_cr_n257), .ZN(U_cr_n244) );
  AOI222_X2 U_cr_U538 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[9]), .B1(U_cr_n168), .B2(hiu_wr_data[17]), .C1(hiu_wr_data[1]), .C2(U_cr_n319), .ZN(U_cr_n546) );
  AOI22_X2 U_cr_U537 ( .A1(hiu_wr_data[25]), .A2(U_cr_n258), .B1(cr_t_rc[3]), 
        .B2(U_cr_n257), .ZN(U_cr_n246) );
  OAI211_X2 U_cr_U536 ( .C1(U_cr_n546), .C2(U_cr_n262), .A(U_cr_n246), .B(
        U_cr_n245), .ZN(U_cr_N414) );
  AOI222_X2 U_cr_U535 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[10]), .B1(
        U_cr_n168), .B2(hiu_wr_data[18]), .C1(hiu_wr_data[2]), .C2(U_cr_n319), 
        .ZN(U_cr_n545) );
  AOI22_X2 U_cr_U534 ( .A1(hiu_wr_data[26]), .A2(U_cr_n258), .B1(
        U_cr_stmg0r_26), .B2(U_cr_n257), .ZN(U_cr_n248) );
  OAI211_X2 U_cr_U533 ( .C1(U_cr_n545), .C2(U_cr_n262), .A(U_cr_n248), .B(
        U_cr_n247), .ZN(U_cr_N415) );
  AOI22_X2 U_cr_U532 ( .A1(hiu_wr_data[28]), .A2(U_cr_n258), .B1(cr_t_xsr[5]), 
        .B2(U_cr_n257), .ZN(U_cr_n252) );
  AOI22_X2 U_cr_U531 ( .A1(hiu_wr_data[27]), .A2(U_cr_n258), .B1(cr_t_xsr[4]), 
        .B2(U_cr_n257), .ZN(U_cr_n250) );
  AOI22_X2 U_cr_U530 ( .A1(hiu_wr_data[29]), .A2(U_cr_n258), .B1(cr_t_xsr[6]), 
        .B2(U_cr_n257), .ZN(U_cr_n254) );
  AOI22_X2 U_cr_U529 ( .A1(hiu_wr_data[31]), .A2(U_cr_n258), .B1(cr_t_xsr[8]), 
        .B2(U_cr_n257), .ZN(U_cr_n261) );
  AOI22_X2 U_cr_U528 ( .A1(hiu_wr_data[30]), .A2(U_cr_n258), .B1(cr_t_xsr[7]), 
        .B2(U_cr_n257), .ZN(U_cr_n256) );
  INV_X4 U_cr_U527 ( .A(U_cr_n318), .ZN(U_cr_n317) );
  AOI221_X2 U_cr_U526 ( .B1(big_endian), .B2(ad_cr_data_mask[3]), .C1(
        U_addrdec_n40), .C2(ad_cr_data_mask[0]), .A(U_cr_n205), .ZN(U_cr_n213)
         );
  AOI222_X2 U_cr_U525 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[5]), .B1(U_cr_n168), .B2(hiu_wr_data[29]), .C1(hiu_wr_data[13]), .C2(U_cr_n319), .ZN(U_cr_n529)
         );
  INV_X4 U_cr_U524 ( .A(U_cr_n215), .ZN(U_cr_n214) );
  AOI22_X2 U_cr_U523 ( .A1(U_cr_n215), .A2(U_cr_n529), .B1(U_cr_n21), .B2(
        U_cr_n214), .ZN(U_cr_N300) );
  AOI222_X2 U_cr_U522 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[4]), .B1(U_cr_n168), .B2(hiu_wr_data[28]), .C1(hiu_wr_data[12]), .C2(U_cr_n319), .ZN(U_cr_n530)
         );
  AOI22_X2 U_cr_U521 ( .A1(U_cr_n215), .A2(U_cr_n530), .B1(U_cr_n66), .B2(
        U_cr_n214), .ZN(U_cr_N299) );
  AOI222_X2 U_cr_U520 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[6]), .B1(U_cr_n168), .B2(hiu_wr_data[30]), .C1(hiu_wr_data[14]), .C2(U_cr_n319), .ZN(U_cr_n528)
         );
  AOI22_X2 U_cr_U519 ( .A1(U_cr_n215), .A2(U_cr_n528), .B1(U_cr_n42), .B2(
        U_cr_n214), .ZN(U_cr_N301) );
  NAND2_X2 U_cr_U518 ( .A1(hiu_haddr[3]), .A2(U_cr_n227), .ZN(U_cr_n263) );
  INV_X4 U_cr_U517 ( .A(U_cr_n273), .ZN(U_cr_n272) );
  AOI22_X2 U_cr_U516 ( .A1(U_cr_n273), .A2(U_cr_n530), .B1(U_cr_n139), .B2(
        U_cr_n272), .ZN(U_cr_N554) );
  AOI22_X2 U_cr_U515 ( .A1(U_cr_n273), .A2(U_cr_n529), .B1(U_cr_n132), .B2(
        U_cr_n272), .ZN(U_cr_N555) );
  AOI22_X2 U_cr_U514 ( .A1(U_cr_n273), .A2(U_cr_n528), .B1(U_cr_n40), .B2(
        U_cr_n272), .ZN(U_cr_N556) );
  AOI221_X2 U_cr_U513 ( .B1(U_cr_n516), .B2(U_cr_n273), .C1(U_cr_n39), .C2(
        U_cr_n272), .A(clear_sr_dp), .ZN(U_cr_N551) );
  AOI22_X2 U_cr_U512 ( .A1(U_cr_n230), .A2(U_cr_n516), .B1(U_cr_n43), .B2(
        U_cr_n229), .ZN(U_cr_N390) );
  AOI222_X2 U_cr_U511 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[7]), .B1(U_cr_n168), .B2(hiu_wr_data[31]), .C1(hiu_wr_data[15]), .C2(U_cr_n319), .ZN(U_cr_n527)
         );
  AOI22_X2 U_cr_U510 ( .A1(U_cr_n230), .A2(U_cr_n527), .B1(U_cr_n133), .B2(
        U_cr_n229), .ZN(U_cr_N396) );
  AOI22_X2 U_cr_U509 ( .A1(U_cr_n230), .A2(U_cr_n531), .B1(U_cr_n120), .B2(
        U_cr_n229), .ZN(U_cr_N392) );
  AOI22_X2 U_cr_U508 ( .A1(U_cr_n230), .A2(U_cr_n529), .B1(U_cr_n54), .B2(
        U_cr_n229), .ZN(U_cr_N394) );
  AOI22_X2 U_cr_U507 ( .A1(U_cr_n313), .A2(U_cr_n531), .B1(U_cr_n156), .B2(
        U_cr_n312), .ZN(U_cr_N736) );
  NOR3_X2 U_cr_U506 ( .A1(U_cr_n320), .A2(U_cr_n316), .A3(U_cr_n315), .ZN(
        U_cr_n525) );
  INV_X4 U_cr_U505 ( .A(U_cr_n525), .ZN(U_cr_n543) );
  AOI22_X2 U_cr_U504 ( .A1(U_cr_n536), .A2(U_cr_n530), .B1(U_cr_n152), .B2(
        U_cr_n538), .ZN(U_cr_n83) );
  AOI22_X2 U_cr_U503 ( .A1(U_cr_n313), .A2(U_cr_n527), .B1(U_cr_n159), .B2(
        U_cr_n312), .ZN(U_cr_N740) );
  AOI22_X2 U_cr_U502 ( .A1(U_cr_n305), .A2(U_cr_n529), .B1(U_cr_n124), .B2(
        U_cr_n304), .ZN(U_cr_N693) );
  AOI22_X2 U_cr_U501 ( .A1(U_cr_n536), .A2(U_cr_n528), .B1(U_cr_n119), .B2(
        U_cr_n538), .ZN(U_cr_n81) );
  AOI22_X2 U_cr_U500 ( .A1(U_cr_n536), .A2(U_cr_n529), .B1(U_cr_n110), .B2(
        U_cr_n538), .ZN(U_cr_n82) );
  AOI22_X2 U_cr_U499 ( .A1(U_cr_n305), .A2(U_cr_n531), .B1(U_cr_n97), .B2(
        U_cr_n304), .ZN(U_cr_N691) );
  NOR3_X2 U_cr_U498 ( .A1(hiu_haddr[2]), .A2(hiu_addr[6]), .A3(U_cr_n315), 
        .ZN(U_cr_n429) );
  INV_X4 U_cr_U497 ( .A(U_cr_n429), .ZN(U_cr_n170) );
  AOI22_X2 U_cr_U496 ( .A1(U_cr_n289), .A2(U_cr_n527), .B1(U_cr_n113), .B2(
        U_cr_n288), .ZN(U_cr_N639) );
  AOI22_X2 U_cr_U495 ( .A1(U_cr_n536), .A2(U_cr_n527), .B1(U_cr_n167), .B2(
        U_cr_n538), .ZN(U_cr_n80) );
  AOI22_X2 U_cr_U494 ( .A1(U_cr_n289), .A2(U_cr_n529), .B1(U_cr_n112), .B2(
        U_cr_n288), .ZN(U_cr_N637) );
  AOI22_X2 U_cr_U493 ( .A1(U_cr_n305), .A2(U_cr_n528), .B1(U_cr_n125), .B2(
        U_cr_n304), .ZN(U_cr_N694) );
  AOI22_X2 U_cr_U492 ( .A1(U_cr_n305), .A2(U_cr_n530), .B1(U_cr_n26), .B2(
        U_cr_n304), .ZN(U_cr_N692) );
  AOI22_X2 U_cr_U491 ( .A1(U_cr_n313), .A2(U_cr_n530), .B1(U_cr_n164), .B2(
        U_cr_n312), .ZN(U_cr_N737) );
  AOI22_X2 U_cr_U490 ( .A1(U_cr_n305), .A2(U_cr_n527), .B1(U_cr_n100), .B2(
        U_cr_n304), .ZN(U_cr_N695) );
  AOI22_X2 U_cr_U489 ( .A1(U_cr_n313), .A2(U_cr_n529), .B1(U_cr_n157), .B2(
        U_cr_n312), .ZN(U_cr_N738) );
  AOI22_X2 U_cr_U488 ( .A1(U_cr_n289), .A2(U_cr_n528), .B1(U_cr_n121), .B2(
        U_cr_n288), .ZN(U_cr_N638) );
  AOI22_X2 U_cr_U487 ( .A1(U_cr_n289), .A2(U_cr_n531), .B1(U_cr_n69), .B2(
        U_cr_n288), .ZN(U_cr_N635) );
  AOI22_X2 U_cr_U486 ( .A1(U_cr_n313), .A2(U_cr_n528), .B1(U_cr_n158), .B2(
        U_cr_n312), .ZN(U_cr_N739) );
  AOI22_X2 U_cr_U485 ( .A1(U_cr_n215), .A2(U_cr_n531), .B1(U_cr_n36), .B2(
        U_cr_n214), .ZN(U_cr_N298) );
  AOI22_X2 U_cr_U484 ( .A1(U_cr_n215), .A2(U_cr_n527), .B1(U_cr_n55), .B2(
        U_cr_n214), .ZN(U_cr_N302) );
  AOI22_X2 U_cr_U483 ( .A1(U_cr_n273), .A2(U_cr_n531), .B1(U_cr_n58), .B2(
        U_cr_n272), .ZN(U_cr_N553) );
  AOI22_X2 U_cr_U482 ( .A1(U_cr_n273), .A2(U_cr_n527), .B1(U_cr_n59), .B2(
        U_cr_n272), .ZN(U_cr_N557) );
  AOI221_X2 U_cr_U481 ( .B1(U_cr_n514), .B2(U_cr_n273), .C1(U_cr_n56), .C2(
        U_cr_n272), .A(ctl_init_done), .ZN(U_cr_N550) );
  INV_X4 U_cr_U480 ( .A(U_cr_n518), .ZN(U_cr_n532) );
  INV_X4 U_cr_U479 ( .A(U_cr_n514), .ZN(U_cr_n537) );
  AOI22_X2 U_cr_U478 ( .A1(U_cr_n230), .A2(U_cr_n514), .B1(U_cr_n20), .B2(
        U_cr_n229), .ZN(U_cr_N389) );
  AOI22_X2 U_cr_U477 ( .A1(U_cr_n230), .A2(U_cr_n530), .B1(U_cr_n128), .B2(
        U_cr_n229), .ZN(U_cr_N393) );
  AOI22_X2 U_cr_U476 ( .A1(U_cr_n230), .A2(U_cr_n528), .B1(U_cr_n149), .B2(
        U_cr_n229), .ZN(U_cr_N395) );
  INV_X4 U_cr_U475 ( .A(U_cr_n25), .ZN(U_cr_n171) );
  INV_X4 U_cr_U474 ( .A(U_cr_n416), .ZN(U_cr_n407) );
  NOR2_X2 U_cr_U473 ( .A1(U_cr_n316), .A2(U_cr_n359), .ZN(U_cr_n321) );
  NAND2_X2 U_cr_U472 ( .A1(hiu_haddr[3]), .A2(U_cr_n321), .ZN(U_cr_n412) );
  AOI21_X2 U_cr_U471 ( .B1(U_cr_n171), .B2(cr_t_wtr[0]), .A(U_cr_n356), .ZN(
        U_cr_n467) );
  NAND2_X2 U_cr_U470 ( .A1(U_cr_n318), .A2(big_endian), .ZN(U_cr_n176) );
  NOR2_X2 U_cr_U469 ( .A1(U_cr_n188), .A2(U_cr_n174), .ZN(U_cr_n177) );
  NAND3_X2 U_cr_U468 ( .A1(U_cr_n176), .A2(U_cr_n177), .A3(U_cr_n175), .ZN(
        U_cr_n180) );
  NOR2_X2 U_cr_U467 ( .A1(U_cr_n182), .A2(big_endian), .ZN(U_cr_n497) );
  NOR2_X2 U_cr_U466 ( .A1(U_cr_n412), .A2(hiu_haddr[2]), .ZN(U_cr_n421) );
  INV_X4 U_cr_U465 ( .A(U_cr_n421), .ZN(U_cr_n431) );
  NAND2_X2 U_cr_U464 ( .A1(U_cr_n357), .A2(U_cr_n431), .ZN(U_cr_n465) );
  OAI22_X2 U_cr_U463 ( .A1(U_cr_n360), .A2(U_cr_n359), .B1(U_cr_n358), .B2(
        U_cr_n26), .ZN(U_cr_n365) );
  AOI22_X2 U_cr_U462 ( .A1(U_cr_n407), .A2(cr_bank_addr_width[1]), .B1(
        U_cr_n169), .B2(cr_t_ref[4]), .ZN(U_cr_n362) );
  NAND3_X2 U_cr_U461 ( .A1(U_cr_n363), .A2(U_cr_n362), .A3(U_cr_n361), .ZN(
        U_cr_n364) );
  AOI211_X2 U_cr_U460 ( .C1(U_cr_n525), .C2(U_cr_n554), .A(U_cr_n365), .B(
        U_cr_n364), .ZN(U_cr_n463) );
  INV_X4 U_cr_U459 ( .A(U_cr_n499), .ZN(U_cr_n469) );
  AOI22_X2 U_cr_U458 ( .A1(U_cr_n407), .A2(n[23]), .B1(U_cr_n430), .B2(
        cr_t_wr[0]), .ZN(U_cr_n368) );
  AOI22_X2 U_cr_U457 ( .A1(U_cr_n422), .A2(U_cr_sctlr_12_), .B1(U_cr_n169), 
        .B2(cr_t_ref[12]), .ZN(U_cr_n367) );
  NAND3_X2 U_cr_U456 ( .A1(U_cr_n368), .A2(U_cr_n367), .A3(U_cr_n366), .ZN(
        U_cr_n369) );
  AOI211_X2 U_cr_U455 ( .C1(U_cr_n171), .C2(cr_t_init[12]), .A(U_cr_n421), .B(
        U_cr_n369), .ZN(U_cr_n462) );
  OAI22_X2 U_cr_U454 ( .A1(U_cr_n463), .A2(U_cr_n469), .B1(U_cr_n462), .B2(
        U_cr_n492), .ZN(U_cr_n370) );
  AOI21_X2 U_cr_U453 ( .B1(U_cr_n497), .B2(U_cr_n465), .A(U_cr_n370), .ZN(
        U_cr_n371) );
  OAI21_X2 U_cr_U452 ( .B1(U_cr_n467), .B2(U_cr_n487), .A(U_cr_n371), .ZN(
        cr_reg_data_out[12]) );
  INV_X4 U_cr_U451 ( .A(U_cr_n497), .ZN(U_cr_n485) );
  OAI22_X2 U_cr_U450 ( .A1(U_cr_n463), .A2(U_cr_n492), .B1(U_cr_n462), .B2(
        U_cr_n469), .ZN(U_cr_n464) );
  AOI21_X2 U_cr_U449 ( .B1(U_cr_n204), .B2(U_cr_n465), .A(U_cr_n464), .ZN(
        U_cr_n466) );
  OAI21_X2 U_cr_U448 ( .B1(U_cr_n467), .B2(U_cr_n485), .A(U_cr_n466), .ZN(
        cr_reg_data_out[4]) );
  AOI22_X2 U_cr_U447 ( .A1(U_cr_n289), .A2(U_cr_n530), .B1(U_cr_n130), .B2(
        U_cr_n288), .ZN(U_cr_N636) );
  AOI22_X2 U_cr_U446 ( .A1(U_cr_n536), .A2(U_cr_n531), .B1(U_cr_n165), .B2(
        U_cr_n538), .ZN(U_cr_n84) );
  AOI22_X2 U_cr_U445 ( .A1(U_cr_n169), .A2(gpo[2]), .B1(U_cr_n171), .B2(
        cr_num_init_ref[2]), .ZN(U_cr_n331) );
  AOI21_X2 U_cr_U444 ( .B1(U_cr_n422), .B2(cr_exn_mode_reg_update), .A(
        U_cr_n333), .ZN(U_cr_n450) );
  AOI22_X2 U_cr_U443 ( .A1(U_cr_n169), .A2(cr_t_ref[10]), .B1(U_cr_n171), .B2(
        cr_t_init[10]), .ZN(U_cr_n339) );
  AOI22_X2 U_cr_U442 ( .A1(U_cr_n407), .A2(n[25]), .B1(U_cr_n430), .B2(
        cr_t_rp[1]), .ZN(U_cr_n338) );
  NAND2_X2 U_cr_U441 ( .A1(U_cr_n321), .A2(U_cr_n320), .ZN(U_cr_n378) );
  AOI211_X2 U_cr_U440 ( .C1(U_cr_n525), .C2(U_cr_n551), .A(U_cr_n393), .B(
        U_cr_n335), .ZN(U_cr_n336) );
  NAND4_X2 U_cr_U439 ( .A1(U_cr_n339), .A2(U_cr_n338), .A3(U_cr_n337), .A4(
        U_cr_n336), .ZN(U_cr_n448) );
  AOI22_X2 U_cr_U438 ( .A1(U_cr_n169), .A2(cr_t_ref[2]), .B1(U_cr_n171), .B2(
        cr_t_init[2]), .ZN(U_cr_n342) );
  NAND3_X2 U_cr_U437 ( .A1(U_cr_n342), .A2(U_cr_n341), .A3(U_cr_n340), .ZN(
        U_cr_n343) );
  AOI211_X2 U_cr_U436 ( .C1(U_cr_n525), .C2(U_cr_n556), .A(U_cr_n393), .B(
        U_cr_n343), .ZN(U_cr_n446) );
  NOR2_X2 U_cr_U435 ( .A1(U_cr_n320), .A2(U_cr_n412), .ZN(U_cr_n392) );
  AOI211_X2 U_cr_U434 ( .C1(U_cr_n169), .C2(U_cr_srefr[26]), .A(U_cr_n344), 
        .B(U_cr_n392), .ZN(U_cr_n445) );
  OAI22_X2 U_cr_U433 ( .A1(U_cr_n446), .A2(U_cr_n469), .B1(U_cr_n445), .B2(
        U_cr_n485), .ZN(U_cr_n345) );
  AOI21_X2 U_cr_U432 ( .B1(U_cr_n203), .B2(U_cr_n448), .A(U_cr_n345), .ZN(
        U_cr_n346) );
  OAI22_X2 U_cr_U431 ( .A1(U_cr_n446), .A2(U_cr_n492), .B1(U_cr_n445), .B2(
        U_cr_n487), .ZN(U_cr_n447) );
  AOI21_X2 U_cr_U430 ( .B1(U_cr_n499), .B2(U_cr_n448), .A(U_cr_n447), .ZN(
        U_cr_n449) );
  OAI21_X2 U_cr_U429 ( .B1(U_cr_n450), .B2(U_cr_n485), .A(U_cr_n449), .ZN(
        cr_reg_data_out[2]) );
  INV_X4 U_cr_U428 ( .A(U_cr_n516), .ZN(U_cr_n534) );
  OAI22_X2 U_cr_U427 ( .A1(U_cr_n391), .A2(U_cr_n34), .B1(U_cr_n170), .B2(
        U_cr_n19), .ZN(U_cr_n372) );
  AOI211_X2 U_cr_U426 ( .C1(U_cr_n171), .C2(cr_t_wtr[1]), .A(U_cr_n421), .B(
        U_cr_n372), .ZN(U_cr_n474) );
  NAND2_X2 U_cr_U425 ( .A1(U_cr_n373), .A2(U_cr_n431), .ZN(U_cr_n472) );
  NAND2_X2 U_cr_U424 ( .A1(U_cr_n375), .A2(U_cr_n374), .ZN(U_cr_n376) );
  AOI211_X2 U_cr_U423 ( .C1(U_cr_n169), .C2(cr_t_ref[13]), .A(U_cr_n377), .B(
        U_cr_n376), .ZN(U_cr_n470) );
  AOI22_X2 U_cr_U422 ( .A1(U_cr_n430), .A2(cr_t_ras_min[3]), .B1(U_cr_n423), 
        .B2(cr_exn_mode_value[5]), .ZN(U_cr_n379) );
  NAND4_X2 U_cr_U421 ( .A1(U_cr_n381), .A2(U_cr_n380), .A3(U_cr_n379), .A4(
        U_cr_n378), .ZN(U_cr_n382) );
  AOI211_X2 U_cr_U420 ( .C1(U_cr_n422), .C2(cr_ref_all_after_sr), .A(U_cr_n383), .B(U_cr_n382), .ZN(U_cr_n468) );
  OAI22_X2 U_cr_U419 ( .A1(U_cr_n470), .A2(U_cr_n492), .B1(U_cr_n468), .B2(
        U_cr_n469), .ZN(U_cr_n384) );
  AOI21_X2 U_cr_U418 ( .B1(U_cr_n497), .B2(U_cr_n472), .A(U_cr_n384), .ZN(
        U_cr_n385) );
  OAI22_X2 U_cr_U417 ( .A1(U_cr_n470), .A2(U_cr_n469), .B1(U_cr_n468), .B2(
        U_cr_n492), .ZN(U_cr_n471) );
  AOI21_X2 U_cr_U416 ( .B1(U_cr_n204), .B2(U_cr_n472), .A(U_cr_n471), .ZN(
        U_cr_n473) );
  OAI21_X2 U_cr_U415 ( .B1(U_cr_n474), .B2(U_cr_n485), .A(U_cr_n473), .ZN(
        cr_reg_data_out[5]) );
  AOI22_X2 U_cr_U414 ( .A1(U_cr_n430), .A2(cr_t_ras_min[1]), .B1(U_cr_n423), 
        .B2(cr_exn_mode_value[3]), .ZN(U_cr_n347) );
  NAND4_X2 U_cr_U413 ( .A1(U_cr_n349), .A2(U_cr_n348), .A3(U_cr_n347), .A4(
        U_cr_n378), .ZN(U_cr_n350) );
  AOI211_X2 U_cr_U412 ( .C1(U_cr_n422), .C2(cr_delayed_precharge), .A(
        U_cr_n351), .B(U_cr_n350), .ZN(U_cr_n461) );
  AOI22_X2 U_cr_U411 ( .A1(U_cr_n430), .A2(cr_t_xsr[4]), .B1(U_cr_n169), .B2(
        U_cr_srefr[27]), .ZN(U_cr_n457) );
  AOI22_X2 U_cr_U410 ( .A1(big_endian), .A2(U_cr_n461), .B1(U_cr_n457), .B2(
        U_addrdec_n40), .ZN(U_cr_n442) );
  AOI22_X2 U_cr_U409 ( .A1(U_cr_n422), .A2(U_cr_n572), .B1(U_cr_n171), .B2(
        cr_num_init_ref[3]), .ZN(U_cr_n352) );
  OAI211_X2 U_cr_U408 ( .C1(U_cr_n391), .C2(U_cr_n32), .A(U_cr_n353), .B(
        U_cr_n352), .ZN(U_cr_n459) );
  AOI22_X2 U_cr_U407 ( .A1(U_cr_n442), .A2(U_cr_n181), .B1(U_cr_n204), .B2(
        U_cr_n459), .ZN(U_cr_n354) );
  AOI22_X2 U_cr_U406 ( .A1(U_cr_n268), .A2(U_cr_n528), .B1(U_cr_n135), .B2(
        U_cr_n267), .ZN(U_cr_N470) );
  AOI22_X2 U_cr_U405 ( .A1(U_cr_n268), .A2(U_cr_n530), .B1(U_cr_n134), .B2(
        U_cr_n267), .ZN(U_cr_N468) );
  AOI22_X2 U_cr_U404 ( .A1(U_cr_n268), .A2(U_cr_n527), .B1(U_cr_n142), .B2(
        U_cr_n267), .ZN(U_cr_N471) );
  AOI22_X2 U_cr_U403 ( .A1(U_cr_n268), .A2(U_cr_n529), .B1(U_cr_n141), .B2(
        U_cr_n267), .ZN(U_cr_N469) );
  AOI22_X2 U_cr_U402 ( .A1(U_cr_n268), .A2(U_cr_n531), .B1(U_cr_n150), .B2(
        U_cr_n267), .ZN(U_cr_N467) );
  OAI22_X2 U_cr_U401 ( .A1(U_cr_n457), .A2(U_cr_n487), .B1(U_cr_n456), .B2(
        U_cr_n469), .ZN(U_cr_n458) );
  AOI21_X2 U_cr_U400 ( .B1(U_cr_n497), .B2(U_cr_n459), .A(U_cr_n458), .ZN(
        U_cr_n460) );
  AOI221_X2 U_cr_U399 ( .B1(big_endian), .B2(ad_cr_data_mask[2]), .C1(
        U_addrdec_n40), .C2(ad_cr_data_mask[1]), .A(U_cr_n205), .ZN(U_cr_n216)
         );
  NOR2_X2 U_cr_U398 ( .A1(U_cr_n396), .A2(U_cr_n544), .ZN(U_cr_n275) );
  INV_X4 U_cr_U397 ( .A(U_cr_n275), .ZN(U_cr_n274) );
  AOI22_X2 U_cr_U396 ( .A1(U_cr_n275), .A2(U_cr_n291), .B1(U_cr_n35), .B2(
        U_cr_n274), .ZN(U_cr_N563) );
  AOI22_X2 U_cr_U395 ( .A1(U_cr_n275), .A2(U_cr_n293), .B1(U_cr_n44), .B2(
        U_cr_n274), .ZN(U_cr_N564) );
  AOI22_X2 U_cr_U394 ( .A1(U_cr_n275), .A2(U_cr_n548), .B1(U_cr_n41), .B2(
        U_cr_n274), .ZN(U_cr_N558) );
  AOI22_X2 U_cr_U393 ( .A1(U_cr_n275), .A2(U_cr_n545), .B1(U_cr_n155), .B2(
        U_cr_n274), .ZN(U_cr_N560) );
  AOI221_X2 U_cr_U392 ( .B1(U_cr_n546), .B2(U_cr_n275), .C1(U_cr_n61), .C2(
        U_cr_n274), .A(ctl_mode_reg_done), .ZN(U_cr_N559) );
  AOI22_X2 U_cr_U391 ( .A1(U_cr_n168), .A2(hiu_wr_data[10]), .B1(
        hiu_wr_data[18]), .B2(U_addrdec_n40), .ZN(U_cr_n517) );
  NAND2_X2 U_cr_U390 ( .A1(U_cr_n223), .A2(U_cr_n240), .ZN(U_cr_n512) );
  NOR2_X2 U_cr_U389 ( .A1(U_cr_n396), .A2(U_cr_n512), .ZN(U_cr_n506) );
  INV_X4 U_cr_U388 ( .A(U_cr_n506), .ZN(U_cr_n508) );
  NAND2_X2 U_cr_U387 ( .A1(U_cr_n238), .A2(U_cr_n223), .ZN(U_cr_n276) );
  NOR2_X2 U_cr_U386 ( .A1(U_cr_n276), .A2(U_cr_n396), .ZN(U_cr_n279) );
  AOI22_X2 U_cr_U385 ( .A1(cr_exn_mode_reg_update), .A2(U_cr_n508), .B1(
        U_cr_n279), .B2(U_cr_n532), .ZN(U_cr_n281) );
  NAND2_X2 U_cr_U384 ( .A1(U_cr_n422), .A2(U_cr_n511), .ZN(U_cr_n280) );
  AOI221_X2 U_cr_U383 ( .B1(U_cr_n517), .B2(U_cr_n281), .C1(U_cr_n280), .C2(
        U_cr_n281), .A(ctl_ext_mode_reg_done), .ZN(U_cr_N567) );
  NAND4_X2 U_cr_U382 ( .A1(U_cr_n411), .A2(U_cr_n410), .A3(U_cr_n409), .A4(
        U_cr_n408), .ZN(U_cr_n495) );
  NAND2_X2 U_cr_U381 ( .A1(U_cr_n13), .A2(big_endian), .ZN(U_cr_n453) );
  AOI21_X2 U_cr_U380 ( .B1(U_cr_n422), .B2(cr_s_ready_valid), .A(U_cr_n414), 
        .ZN(U_cr_n415) );
  OAI21_X2 U_cr_U379 ( .B1(U_cr_n416), .B2(U_cr_n31), .A(U_cr_n415), .ZN(
        U_cr_n494) );
  NAND2_X2 U_cr_U378 ( .A1(U_cr_n13), .A2(U_addrdec_n40), .ZN(U_cr_n451) );
  OAI22_X2 U_cr_U377 ( .A1(U_cr_n418), .A2(U_cr_n453), .B1(U_cr_n417), .B2(
        U_cr_n451), .ZN(cr_reg_data_out[17]) );
  AOI22_X2 U_cr_U376 ( .A1(U_cr_n430), .A2(cr_t_xsr[8]), .B1(U_cr_n429), .B2(
        U_cr_srefr[31]), .ZN(U_cr_n484) );
  NAND4_X2 U_cr_U375 ( .A1(U_cr_n402), .A2(U_cr_n401), .A3(U_cr_n400), .A4(
        U_cr_n399), .ZN(U_cr_n481) );
  AOI22_X2 U_cr_U374 ( .A1(U_cr_n407), .A2(s_sa[0]), .B1(U_cr_n169), .B2(
        cr_t_ref[15]), .ZN(U_cr_n405) );
  NAND2_X2 U_cr_U373 ( .A1(U_cr_n405), .A2(U_cr_n404), .ZN(U_cr_n406) );
  AOI21_X2 U_cr_U372 ( .B1(U_cr_sctlr_15_), .B2(U_cr_n422), .A(U_cr_n406), 
        .ZN(U_cr_n438) );
  AOI22_X2 U_cr_U371 ( .A1(U_cr_n430), .A2(cr_t_rc[1]), .B1(U_cr_n169), .B2(
        gpo[7]), .ZN(U_cr_n437) );
  AOI22_X2 U_cr_U370 ( .A1(big_endian), .A2(U_cr_n438), .B1(U_cr_n437), .B2(
        U_addrdec_n40), .ZN(U_cr_n482) );
  AOI22_X2 U_cr_U369 ( .A1(U_cr_n481), .A2(U_cr_n203), .B1(U_cr_n181), .B2(
        U_cr_n482), .ZN(U_cr_n483) );
  AOI22_X2 U_cr_U368 ( .A1(hiu_wr_data[8]), .A2(U_cr_n168), .B1(
        hiu_wr_data[16]), .B2(U_addrdec_n40), .ZN(U_cr_n513) );
  AOI22_X2 U_cr_U367 ( .A1(U_cr_n279), .A2(U_cr_n537), .B1(U_cr_sctlr_16_), 
        .B2(U_cr_n508), .ZN(U_cr_n277) );
  OAI21_X2 U_cr_U366 ( .B1(U_cr_n513), .B2(U_cr_n280), .A(U_cr_n277), .ZN(
        U_cr_N565) );
  AOI22_X2 U_cr_U365 ( .A1(hiu_wr_data[9]), .A2(U_cr_n168), .B1(
        hiu_wr_data[17]), .B2(U_addrdec_n40), .ZN(U_cr_n515) );
  AOI22_X2 U_cr_U364 ( .A1(U_cr_n279), .A2(U_cr_n534), .B1(cr_s_ready_valid), 
        .B2(U_cr_n508), .ZN(U_cr_n278) );
  OAI21_X2 U_cr_U363 ( .B1(U_cr_n515), .B2(U_cr_n280), .A(U_cr_n278), .ZN(
        U_cr_N566) );
  AOI22_X2 U_cr_U362 ( .A1(hiu_wr_data[11]), .A2(U_cr_n168), .B1(
        hiu_wr_data[19]), .B2(U_addrdec_n40), .ZN(U_cr_n519) );
  OAI22_X2 U_cr_U361 ( .A1(U_cr_n508), .A2(U_cr_n507), .B1(U_cr_n572), .B2(
        U_cr_n506), .ZN(U_cr_n509) );
  INV_X4 U_cr_U360 ( .A(U_cr_n509), .ZN(U_cr_n73) );
  AOI22_X2 U_cr_U359 ( .A1(big_endian), .A2(U_cr_n481), .B1(U_cr_n403), .B2(
        U_addrdec_n40), .ZN(U_cr_n455) );
  AOI22_X2 U_cr_U358 ( .A1(U_cr_n275), .A2(U_cr_n314), .B1(U_cr_n18), .B2(
        U_cr_n274), .ZN(U_cr_N561) );
  AOI22_X2 U_cr_U357 ( .A1(U_cr_n275), .A2(U_cr_n290), .B1(U_cr_n27), .B2(
        U_cr_n274), .ZN(U_cr_N562) );
  AOI21_X2 U_cr_U356 ( .B1(cr_do_initialize), .B2(U_cr_n422), .A(U_cr_n393), 
        .ZN(U_cr_n323) );
  NAND4_X2 U_cr_U355 ( .A1(U_cr_n325), .A2(U_cr_n324), .A3(U_cr_n323), .A4(
        U_cr_n322), .ZN(U_cr_n490) );
  AOI22_X2 U_cr_U354 ( .A1(U_cr_n169), .A2(gpo[0]), .B1(U_cr_n171), .B2(
        cr_num_init_ref[0]), .ZN(U_cr_n326) );
  AOI21_X2 U_cr_U353 ( .B1(U_cr_n422), .B2(U_cr_sctlr_16_), .A(U_cr_n328), 
        .ZN(U_cr_n488) );
  OAI22_X2 U_cr_U352 ( .A1(U_cr_n488), .A2(U_cr_n487), .B1(U_cr_n486), .B2(
        U_cr_n485), .ZN(U_cr_n489) );
  AOI21_X2 U_cr_U351 ( .B1(U_cr_n499), .B2(U_cr_n490), .A(U_cr_n489), .ZN(
        U_cr_n491) );
  OAI22_X2 U_cr_U350 ( .A1(U_cr_n488), .A2(U_cr_n485), .B1(U_cr_n486), .B2(
        U_cr_n487), .ZN(U_cr_n329) );
  AOI21_X2 U_cr_U349 ( .B1(U_cr_n203), .B2(U_cr_n490), .A(U_cr_n329), .ZN(
        U_cr_n330) );
  OAI21_X2 U_cr_U348 ( .B1(U_cr_n493), .B2(U_cr_n469), .A(U_cr_n330), .ZN(
        cr_reg_data_out[0]) );
  INV_X4 U_cr_U347 ( .A(U_cr_n221), .ZN(U_cr_n220) );
  AOI22_X2 U_cr_U346 ( .A1(U_cr_n221), .A2(U_cr_n541), .B1(U_cr_n38), .B2(
        U_cr_n220), .ZN(U_cr_N306) );
  AOI22_X2 U_cr_U345 ( .A1(U_cr_n221), .A2(U_cr_n293), .B1(U_cr_n52), .B2(
        U_cr_n220), .ZN(U_cr_N310) );
  INV_X4 U_cr_U344 ( .A(U_cr_n276), .ZN(U_cr_n510) );
  NAND2_X2 U_cr_U343 ( .A1(U_cr_n510), .A2(U_cr_n430), .ZN(U_cr_n233) );
  NAND2_X2 U_cr_U342 ( .A1(U_cr_n511), .A2(U_cr_n430), .ZN(U_cr_n235) );
  NOR2_X2 U_cr_U341 ( .A1(U_cr_n512), .A2(U_cr_n391), .ZN(U_cr_n234) );
  OAI222_X2 U_cr_U340 ( .A1(U_cr_n233), .A2(U_cr_n531), .B1(U_cr_n235), .B2(
        U_cr_n519), .C1(U_cr_n32), .C2(U_cr_n234), .ZN(U_cr_N408) );
  AOI22_X2 U_cr_U339 ( .A1(hiu_wr_data[14]), .A2(U_cr_n168), .B1(
        hiu_wr_data[22]), .B2(U_addrdec_n40), .ZN(U_cr_n295) );
  OAI222_X2 U_cr_U338 ( .A1(U_cr_n235), .A2(U_cr_n295), .B1(U_cr_n64), .B2(
        U_cr_n234), .C1(U_cr_n233), .C2(U_cr_n528), .ZN(U_cr_N411) );
  OAI222_X2 U_cr_U337 ( .A1(U_cr_n233), .A2(U_cr_n514), .B1(U_cr_n235), .B2(
        U_cr_n513), .C1(U_cr_n104), .C2(U_cr_n234), .ZN(U_cr_N405) );
  AOI22_X2 U_cr_U336 ( .A1(U_cr_n221), .A2(U_cr_n545), .B1(U_cr_n22), .B2(
        U_cr_n220), .ZN(U_cr_N305) );
  AOI22_X2 U_cr_U335 ( .A1(U_cr_n221), .A2(U_cr_n546), .B1(U_cr_n63), .B2(
        U_cr_n220), .ZN(U_cr_N304) );
  AOI22_X2 U_cr_U334 ( .A1(U_cr_n221), .A2(U_cr_n548), .B1(U_cr_n70), .B2(
        U_cr_n220), .ZN(U_cr_N303) );
  AOI22_X2 U_cr_U333 ( .A1(U_cr_n221), .A2(U_cr_n314), .B1(U_cr_n65), .B2(
        U_cr_n220), .ZN(U_cr_N307) );
  NAND2_X2 U_cr_U332 ( .A1(U_cr_n510), .A2(U_cr_n169), .ZN(U_cr_n299) );
  NAND2_X2 U_cr_U331 ( .A1(U_cr_n511), .A2(U_cr_n169), .ZN(U_cr_n298) );
  NOR2_X2 U_cr_U330 ( .A1(U_cr_n512), .A2(U_cr_n170), .ZN(U_cr_n296) );
  OAI222_X2 U_cr_U329 ( .A1(U_cr_n299), .A2(U_cr_n531), .B1(U_cr_n298), .B2(
        U_cr_n519), .C1(U_cr_n49), .C2(U_cr_n296), .ZN(U_cr_N651) );
  AOI22_X2 U_cr_U328 ( .A1(hiu_wr_data[12]), .A2(U_cr_n168), .B1(
        hiu_wr_data[20]), .B2(U_addrdec_n40), .ZN(U_cr_n520) );
  OAI222_X2 U_cr_U327 ( .A1(U_cr_n299), .A2(U_cr_n530), .B1(U_cr_n298), .B2(
        U_cr_n520), .C1(U_cr_n50), .C2(U_cr_n296), .ZN(U_cr_N652) );
  AOI22_X2 U_cr_U326 ( .A1(hiu_wr_data[13]), .A2(U_cr_n168), .B1(
        hiu_wr_data[21]), .B2(U_addrdec_n40), .ZN(U_cr_n522) );
  OAI222_X2 U_cr_U325 ( .A1(U_cr_n235), .A2(U_cr_n522), .B1(U_cr_n34), .B2(
        U_cr_n234), .C1(U_cr_n233), .C2(U_cr_n529), .ZN(U_cr_N410) );
  AOI22_X2 U_cr_U324 ( .A1(hiu_wr_data[15]), .A2(U_cr_n168), .B1(
        hiu_wr_data[23]), .B2(U_addrdec_n40), .ZN(U_cr_n297) );
  OAI222_X2 U_cr_U323 ( .A1(U_cr_n235), .A2(U_cr_n297), .B1(U_cr_n106), .B2(
        U_cr_n234), .C1(U_cr_n233), .C2(U_cr_n527), .ZN(U_cr_N412) );
  OAI222_X2 U_cr_U322 ( .A1(U_cr_n299), .A2(U_cr_n529), .B1(U_cr_n298), .B2(
        U_cr_n522), .C1(U_cr_n19), .C2(U_cr_n296), .ZN(U_cr_N653) );
  OAI222_X2 U_cr_U321 ( .A1(U_cr_n233), .A2(U_cr_n530), .B1(U_cr_n235), .B2(
        U_cr_n520), .C1(U_cr_n33), .C2(U_cr_n234), .ZN(U_cr_N409) );
  OAI222_X2 U_cr_U320 ( .A1(U_cr_n299), .A2(U_cr_n527), .B1(U_cr_n298), .B2(
        U_cr_n297), .C1(U_cr_n51), .C2(U_cr_n296), .ZN(U_cr_N655) );
  OAI222_X2 U_cr_U319 ( .A1(U_cr_n299), .A2(U_cr_n528), .B1(U_cr_n298), .B2(
        U_cr_n295), .C1(U_cr_n46), .C2(U_cr_n296), .ZN(U_cr_N654) );
  OAI222_X2 U_cr_U318 ( .A1(U_cr_n299), .A2(U_cr_n516), .B1(U_cr_n298), .B2(
        U_cr_n515), .C1(U_cr_n29), .C2(U_cr_n296), .ZN(U_cr_N649) );
  OAI222_X2 U_cr_U317 ( .A1(U_cr_n299), .A2(U_cr_n514), .B1(U_cr_n298), .B2(
        U_cr_n513), .C1(U_cr_n47), .C2(U_cr_n296), .ZN(U_cr_N648) );
  INV_X4 U_cr_U316 ( .A(U_cr_n307), .ZN(U_cr_n306) );
  AOI22_X2 U_cr_U315 ( .A1(U_cr_n307), .A2(U_cr_n546), .B1(U_cr_n101), .B2(
        U_cr_n306), .ZN(U_cr_N697) );
  INV_X4 U_cr_U314 ( .A(U_cr_n542), .ZN(U_cr_n540) );
  AOI22_X2 U_cr_U313 ( .A1(U_cr_n542), .A2(U_cr_n541), .B1(U_cr_n163), .B2(
        U_cr_n540), .ZN(U_cr_n91) );
  AOI22_X2 U_cr_U312 ( .A1(U_cr_n307), .A2(U_cr_n545), .B1(U_cr_n71), .B2(
        U_cr_n306), .ZN(U_cr_N698) );
  AOI22_X2 U_cr_U311 ( .A1(U_cr_n307), .A2(U_cr_n541), .B1(U_cr_n102), .B2(
        U_cr_n306), .ZN(U_cr_N699) );
  AOI22_X2 U_cr_U310 ( .A1(U_cr_n307), .A2(U_cr_n548), .B1(U_cr_n126), .B2(
        U_cr_n306), .ZN(U_cr_N696) );
  AOI22_X2 U_cr_U309 ( .A1(U_cr_n542), .A2(U_cr_n546), .B1(U_cr_n162), .B2(
        U_cr_n540), .ZN(U_cr_n89) );
  AOI22_X2 U_cr_U308 ( .A1(U_cr_n542), .A2(U_cr_n545), .B1(U_cr_n37), .B2(
        U_cr_n540), .ZN(U_cr_n90) );
  AOI22_X2 U_cr_U307 ( .A1(U_cr_n307), .A2(U_cr_n314), .B1(U_cr_n103), .B2(
        U_cr_n306), .ZN(U_cr_N700) );
  AOI22_X2 U_cr_U306 ( .A1(U_cr_n542), .A2(U_cr_n548), .B1(U_cr_n161), .B2(
        U_cr_n540), .ZN(U_cr_n88) );
  AOI22_X2 U_cr_U305 ( .A1(U_cr_n542), .A2(U_cr_n314), .B1(U_cr_n160), .B2(
        U_cr_n540), .ZN(U_cr_N745) );
  OAI222_X2 U_cr_U304 ( .A1(U_cr_n233), .A2(U_cr_n516), .B1(U_cr_n235), .B2(
        U_cr_n515), .C1(U_cr_n72), .C2(U_cr_n234), .ZN(U_cr_N406) );
  OAI222_X2 U_cr_U303 ( .A1(U_cr_n299), .A2(U_cr_n518), .B1(U_cr_n298), .B2(
        U_cr_n517), .C1(U_cr_n48), .C2(U_cr_n296), .ZN(U_cr_N650) );
  NAND2_X2 U_cr_U302 ( .A1(U_cr_n511), .A2(U_cr_n407), .ZN(U_cr_n226) );
  NOR2_X2 U_cr_U301 ( .A1(U_cr_n512), .A2(U_cr_n416), .ZN(U_cr_n225) );
  NAND2_X2 U_cr_U300 ( .A1(U_cr_n510), .A2(U_cr_n407), .ZN(U_cr_n224) );
  OAI222_X2 U_cr_U299 ( .A1(U_cr_n226), .A2(U_cr_n519), .B1(U_cr_n62), .B2(
        U_cr_n225), .C1(U_cr_n224), .C2(U_cr_n531), .ZN(U_cr_N314) );
  AOI22_X2 U_cr_U298 ( .A1(U_cr_n499), .A2(U_cr_n495), .B1(U_cr_n497), .B2(
        U_cr_n494), .ZN(U_cr_n434) );
  NAND4_X2 U_cr_U297 ( .A1(U_cr_n428), .A2(U_cr_n427), .A3(U_cr_n426), .A4(
        U_cr_n425), .ZN(U_cr_n498) );
  NAND2_X2 U_cr_U296 ( .A1(U_cr_n432), .A2(U_cr_n431), .ZN(U_cr_n496) );
  AOI22_X2 U_cr_U295 ( .A1(U_cr_n203), .A2(U_cr_n498), .B1(U_cr_n204), .B2(
        U_cr_n496), .ZN(U_cr_n433) );
  NAND2_X2 U_cr_U294 ( .A1(U_cr_n434), .A2(U_cr_n433), .ZN(cr_reg_data_out[1])
         );
  AOI22_X2 U_cr_U293 ( .A1(U_cr_n203), .A2(U_cr_n495), .B1(U_cr_n204), .B2(
        U_cr_n494), .ZN(U_cr_n501) );
  AOI22_X2 U_cr_U292 ( .A1(U_cr_n499), .A2(U_cr_n498), .B1(U_cr_n497), .B2(
        U_cr_n496), .ZN(U_cr_n500) );
  NAND2_X2 U_cr_U291 ( .A1(U_cr_n501), .A2(U_cr_n500), .ZN(cr_reg_data_out[9])
         );
  OAI222_X2 U_cr_U290 ( .A1(U_cr_n226), .A2(U_cr_n520), .B1(U_cr_n57), .B2(
        U_cr_n225), .C1(U_cr_n224), .C2(U_cr_n530), .ZN(U_cr_N315) );
  OAI222_X2 U_cr_U289 ( .A1(U_cr_n233), .A2(U_cr_n518), .B1(U_cr_n235), .B2(
        U_cr_n517), .C1(U_cr_n108), .C2(U_cr_n234), .ZN(U_cr_N407) );
  NAND2_X2 U_cr_U288 ( .A1(U_cr_n510), .A2(U_cr_n171), .ZN(U_cr_n524) );
  NAND2_X2 U_cr_U287 ( .A1(U_cr_n511), .A2(U_cr_n171), .ZN(U_cr_n523) );
  NOR2_X2 U_cr_U286 ( .A1(U_cr_n512), .A2(U_cr_n25), .ZN(U_cr_n521) );
  OAI222_X2 U_cr_U285 ( .A1(U_cr_n524), .A2(U_cr_n516), .B1(U_cr_n523), .B2(
        U_cr_n515), .C1(U_cr_n117), .C2(U_cr_n521), .ZN(U_cr_n75) );
  OAI222_X2 U_cr_U284 ( .A1(U_cr_n524), .A2(U_cr_n514), .B1(U_cr_n523), .B2(
        U_cr_n513), .C1(U_cr_n115), .C2(U_cr_n521), .ZN(U_cr_n74) );
  AOI22_X2 U_cr_U283 ( .A1(U_cr_n294), .A2(U_cr_n314), .B1(U_cr_n122), .B2(
        U_cr_n292), .ZN(U_cr_N644) );
  AOI22_X2 U_cr_U282 ( .A1(U_cr_n270), .A2(U_cr_n314), .B1(U_cr_n131), .B2(
        U_cr_n269), .ZN(U_cr_N476) );
  AOI22_X2 U_cr_U281 ( .A1(U_cr_n294), .A2(U_cr_n291), .B1(U_cr_n123), .B2(
        U_cr_n292), .ZN(U_cr_N646) );
  AOI22_X2 U_cr_U280 ( .A1(U_cr_n294), .A2(U_cr_n293), .B1(U_cr_n114), .B2(
        U_cr_n292), .ZN(U_cr_N647) );
  AOI22_X2 U_cr_U279 ( .A1(U_cr_n270), .A2(U_cr_n545), .B1(U_cr_n137), .B2(
        U_cr_n269), .ZN(U_cr_N474) );
  AOI22_X2 U_cr_U278 ( .A1(U_cr_n294), .A2(U_cr_n541), .B1(U_cr_n111), .B2(
        U_cr_n292), .ZN(U_cr_N643) );
  AOI22_X2 U_cr_U277 ( .A1(U_cr_n270), .A2(U_cr_n290), .B1(U_cr_n145), .B2(
        U_cr_n269), .ZN(U_cr_N477) );
  AOI22_X2 U_cr_U276 ( .A1(U_cr_n232), .A2(U_cr_n290), .B1(U_cr_n67), .B2(
        U_cr_n231), .ZN(U_cr_N402) );
  AOI22_X2 U_cr_U275 ( .A1(U_cr_n270), .A2(U_cr_n546), .B1(U_cr_n143), .B2(
        U_cr_n269), .ZN(U_cr_N473) );
  AOI22_X2 U_cr_U274 ( .A1(U_cr_n294), .A2(U_cr_n546), .B1(U_cr_n105), .B2(
        U_cr_n292), .ZN(U_cr_N641) );
  AOI22_X2 U_cr_U273 ( .A1(U_cr_n232), .A2(U_cr_n546), .B1(U_cr_n45), .B2(
        U_cr_n231), .ZN(U_cr_N398) );
  AOI22_X2 U_cr_U272 ( .A1(U_cr_n270), .A2(U_cr_n541), .B1(U_cr_n144), .B2(
        U_cr_n269), .ZN(U_cr_N475) );
  AOI22_X2 U_cr_U271 ( .A1(U_cr_n232), .A2(U_cr_n548), .B1(U_cr_n140), .B2(
        U_cr_n231), .ZN(U_cr_N397) );
  AOI22_X2 U_cr_U270 ( .A1(U_cr_n294), .A2(U_cr_n548), .B1(U_cr_n118), .B2(
        U_cr_n292), .ZN(U_cr_N640) );
  AOI22_X2 U_cr_U269 ( .A1(U_cr_n270), .A2(U_cr_n548), .B1(U_cr_n136), .B2(
        U_cr_n269), .ZN(U_cr_N472) );
  AOI22_X2 U_cr_U268 ( .A1(U_cr_n270), .A2(U_cr_n291), .B1(U_cr_n138), .B2(
        U_cr_n269), .ZN(U_cr_N478) );
  AOI22_X2 U_cr_U267 ( .A1(U_cr_n232), .A2(U_cr_n541), .B1(U_cr_n148), .B2(
        U_cr_n231), .ZN(U_cr_N400) );
  AOI22_X2 U_cr_U266 ( .A1(U_cr_n270), .A2(U_cr_n293), .B1(U_cr_n146), .B2(
        U_cr_n269), .ZN(U_cr_N479) );
  AOI22_X2 U_cr_U265 ( .A1(U_cr_n294), .A2(U_cr_n290), .B1(U_cr_n68), .B2(
        U_cr_n292), .ZN(U_cr_N645) );
  OAI222_X2 U_cr_U264 ( .A1(U_cr_n524), .A2(U_cr_n518), .B1(U_cr_n523), .B2(
        U_cr_n517), .C1(U_cr_n116), .C2(U_cr_n521), .ZN(U_cr_n76) );
  OAI222_X2 U_cr_U263 ( .A1(U_cr_n524), .A2(U_cr_n531), .B1(U_cr_n523), .B2(
        U_cr_n519), .C1(U_cr_n109), .C2(U_cr_n521), .ZN(U_cr_n77) );
  OAI222_X2 U_cr_U262 ( .A1(U_cr_n524), .A2(U_cr_n530), .B1(U_cr_n523), .B2(
        U_cr_n520), .C1(U_cr_n53), .C2(U_cr_n521), .ZN(U_cr_n78) );
  OAI222_X2 U_cr_U261 ( .A1(U_cr_n524), .A2(U_cr_n529), .B1(U_cr_n523), .B2(
        U_cr_n522), .C1(U_cr_n60), .C2(U_cr_n521), .ZN(U_cr_n79) );
  OAI22_X2 U_cr_U260 ( .A1(U_cr_n488), .A2(U_cr_n451), .B1(U_cr_n493), .B2(
        U_cr_n453), .ZN(cr_reg_data_out[16]) );
  OAI222_X2 U_cr_U259 ( .A1(U_cr_n224), .A2(U_cr_n518), .B1(U_cr_n226), .B2(
        U_cr_n517), .C1(U_cr_n30), .C2(U_cr_n225), .ZN(U_cr_N313) );
  NOR2_X2 U_cr_U258 ( .A1(U_cr_n544), .A2(U_cr_n543), .ZN(U_cr_n549) );
  INV_X4 U_cr_U257 ( .A(U_cr_n549), .ZN(U_cr_n547) );
  AOI22_X2 U_cr_U256 ( .A1(U_cr_n549), .A2(U_cr_n548), .B1(U_cr_n154), .B2(
        U_cr_n547), .ZN(U_cr_n94) );
  AOI22_X2 U_cr_U255 ( .A1(U_cr_n549), .A2(U_cr_n545), .B1(U_cr_n153), .B2(
        U_cr_n547), .ZN(U_cr_n92) );
  AOI22_X2 U_cr_U254 ( .A1(U_cr_n232), .A2(U_cr_n293), .B1(U_cr_n151), .B2(
        U_cr_n231), .ZN(U_cr_N404) );
  AOI22_X2 U_cr_U253 ( .A1(U_cr_n232), .A2(U_cr_n291), .B1(U_cr_n127), .B2(
        U_cr_n231), .ZN(U_cr_N403) );
  AOI22_X2 U_cr_U252 ( .A1(U_cr_n232), .A2(U_cr_n314), .B1(U_cr_n107), .B2(
        U_cr_n231), .ZN(U_cr_N401) );
  AOI22_X2 U_cr_U251 ( .A1(U_cr_n294), .A2(U_cr_n545), .B1(U_cr_n129), .B2(
        U_cr_n292), .ZN(U_cr_N642) );
  AOI22_X2 U_cr_U250 ( .A1(U_cr_n232), .A2(U_cr_n545), .B1(U_cr_n147), .B2(
        U_cr_n231), .ZN(U_cr_N399) );
  OAI222_X2 U_cr_U249 ( .A1(U_cr_n224), .A2(U_cr_n514), .B1(U_cr_n226), .B2(
        U_cr_n513), .C1(U_cr_n28), .C2(U_cr_n225), .ZN(U_cr_N311) );
  OAI22_X2 U_cr_U248 ( .A1(U_cr_n445), .A2(U_cr_n451), .B1(U_cr_n446), .B2(
        U_cr_n453), .ZN(cr_reg_data_out[26]) );
  OAI22_X2 U_cr_U247 ( .A1(U_cr_n419), .A2(U_cr_n453), .B1(U_cr_n450), .B2(
        U_cr_n451), .ZN(cr_reg_data_out[18]) );
  OAI222_X2 U_cr_U246 ( .A1(U_cr_n226), .A2(U_cr_n515), .B1(U_cr_n224), .B2(
        U_cr_n516), .C1(U_cr_n31), .C2(U_cr_n225), .ZN(U_cr_N312) );
  AOI21_X2 U_cr_U245 ( .B1(U_cr_n169), .B2(cr_t_ref[14]), .A(U_cr_n393), .ZN(
        U_cr_n395) );
  OAI211_X2 U_cr_U244 ( .C1(U_cr_n396), .C2(U_cr_n35), .A(U_cr_n395), .B(
        U_cr_n394), .ZN(U_cr_n478) );
  OAI22_X2 U_cr_U243 ( .A1(U_cr_n436), .A2(U_cr_n451), .B1(U_cr_n435), .B2(
        U_cr_n453), .ZN(cr_reg_data_out[22]) );
  AOI22_X2 U_cr_U242 ( .A1(U_cr_n549), .A2(U_cr_n546), .B1(U_cr_n166), .B2(
        U_cr_n547), .ZN(U_cr_n93) );
  OAI22_X2 U_cr_U241 ( .A1(U_cr_n462), .A2(U_cr_n453), .B1(U_cr_n467), .B2(
        U_cr_n451), .ZN(cr_reg_data_out[20]) );
  OAI22_X2 U_cr_U240 ( .A1(U_cr_n441), .A2(U_cr_n451), .B1(U_cr_n440), .B2(
        U_cr_n453), .ZN(cr_reg_data_out[25]) );
  OAI22_X2 U_cr_U239 ( .A1(U_cr_n486), .A2(U_cr_n451), .B1(U_cr_n439), .B2(
        U_cr_n453), .ZN(cr_reg_data_out[24]) );
  OAI22_X2 U_cr_U238 ( .A1(U_cr_n443), .A2(U_cr_n451), .B1(U_cr_n463), .B2(
        U_cr_n453), .ZN(cr_reg_data_out[28]) );
  OAI22_X2 U_cr_U237 ( .A1(U_cr_n468), .A2(U_cr_n453), .B1(U_cr_n444), .B2(
        U_cr_n451), .ZN(cr_reg_data_out[29]) );
  OAI22_X2 U_cr_U236 ( .A1(U_cr_n456), .A2(U_cr_n453), .B1(U_cr_n420), .B2(
        U_cr_n451), .ZN(cr_reg_data_out[19]) );
  NAND4_X2 U_cr_U235 ( .A1(U_cr_n389), .A2(U_cr_n388), .A3(U_cr_n387), .A4(
        U_cr_n386), .ZN(U_cr_n475) );
  AOI22_X2 U_cr_U234 ( .A1(U_cr_n499), .A2(U_cr_n475), .B1(U_cr_n204), .B2(
        U_cr_n476), .ZN(U_cr_n398) );
  AOI22_X2 U_cr_U233 ( .A1(U_cr_n497), .A2(U_cr_n477), .B1(U_cr_n203), .B2(
        U_cr_n478), .ZN(U_cr_n397) );
  NAND2_X2 U_cr_U232 ( .A1(U_cr_n398), .A2(U_cr_n397), .ZN(cr_reg_data_out[14]) );
  OAI22_X2 U_cr_U231 ( .A1(U_cr_n470), .A2(U_cr_n453), .B1(U_cr_n474), .B2(
        U_cr_n451), .ZN(cr_reg_data_out[21]) );
  AOI22_X2 U_cr_U230 ( .A1(U_cr_n497), .A2(U_cr_n476), .B1(U_cr_n203), .B2(
        U_cr_n475), .ZN(U_cr_n480) );
  AOI22_X2 U_cr_U229 ( .A1(U_cr_n499), .A2(U_cr_n478), .B1(U_cr_n204), .B2(
        U_cr_n477), .ZN(U_cr_n479) );
  NAND2_X2 U_cr_U228 ( .A1(U_cr_n480), .A2(U_cr_n479), .ZN(cr_reg_data_out[6])
         );
  OAI22_X2 U_cr_U227 ( .A1(U_cr_n454), .A2(U_cr_n453), .B1(U_cr_n452), .B2(
        U_cr_n451), .ZN(cr_reg_data_out[30]) );
  NOR2_X2 U_cr_U226 ( .A1(U_cr_n18), .A2(U_cr_n27), .ZN(U_cr_n206) );
  NAND2_X2 U_cr_U225 ( .A1(U_cr_sctlr_14_), .A2(U_cr_n206), .ZN(U_cr_n208) );
  NAND2_X2 U_cr_U224 ( .A1(U_cr_sctlr_15_), .A2(U_cr_n209), .ZN(U_cr_n210) );
  AOI22_X2 U_cr_U223 ( .A1(U_cr_sctlr_15_), .A2(U_cr_n209), .B1(U_cr_n208), 
        .B2(U_cr_n44), .ZN(U_cr_N573) );
  NAND2_X2 U_cr_U222 ( .A1(U_cr_stmg0r_0_), .A2(U_cr_stmg0r_1_), .ZN(U_cr_n282) );
  AOI21_X2 U_cr_U221 ( .B1(U_cr_n18), .B2(U_cr_n27), .A(U_cr_n206), .ZN(
        U_cr_N571) );
  INV_X4 U_cr_U219 ( .A(U_cr_n193), .ZN(U_cr_n186) );
  NOR2_X2 U_cr_U218 ( .A1(U_cr_n320), .A2(U_cr_n308), .ZN(U_cr_n423) );
  AOI22_X2 U_cr_U217 ( .A1(U_cr_n422), .A2(U_cr_n559), .B1(U_cr_n423), .B2(
        cr_exn_mode_value[10]), .ZN(U_cr_n337) );
  NOR2_X2 U_cr_U216 ( .A1(hiu_haddr[3]), .A2(U_cr_n378), .ZN(U_cr_n393) );
  AOI22_X2 U_cr_U215 ( .A1(U_cr_n422), .A2(U_cr_sctlr_13_), .B1(
        cr_s_data_width_early_0_), .B2(U_cr_n407), .ZN(U_cr_n374) );
  AOI22_X2 U_cr_U214 ( .A1(U_cr_n422), .A2(s_read_pipe[1]), .B1(U_cr_n169), 
        .B2(cr_t_ref[7]), .ZN(U_cr_n402) );
  NOR2_X2 U_cr_U213 ( .A1(n27), .A2(U_addrdec_n40), .ZN(U_cr_n319) );
  NAND2_X1 U_cr_U212 ( .A1(U_cr_n187), .A2(U_cr_cr_cs_2_), .ZN(U_cr_n202) );
  NOR2_X2 U_cr_U211 ( .A1(U_cr_n396), .A2(U_cr_n526), .ZN(U_cr_n273) );
  INV_X4 U_cr_U210 ( .A(U_cr_n170), .ZN(U_cr_n169) );
  AOI22_X2 U_cr_U209 ( .A1(U_cr_n422), .A2(cr_ref_all_before_sr), .B1(
        U_cr_n424), .B2(U_cr_n566), .ZN(U_cr_n361) );
  AOI22_X2 U_cr_U208 ( .A1(U_cr_n424), .A2(U_cr_n571), .B1(U_cr_n423), .B2(
        cr_exn_mode_value[12]), .ZN(U_cr_n366) );
  AOI22_X2 U_cr_U207 ( .A1(U_cr_n422), .A2(cr_do_power_down), .B1(U_cr_n430), 
        .B2(cr_t_ras_min[0]), .ZN(U_cr_n341) );
  AOI22_X2 U_cr_U206 ( .A1(U_cr_n424), .A2(U_cr_n568), .B1(U_cr_n423), .B2(
        cr_exn_mode_value[2]), .ZN(U_cr_n340) );
  AOI22_X2 U_cr_U205 ( .A1(U_cr_n424), .A2(U_cr_n561), .B1(U_cr_n423), .B2(
        cr_exn_mode_value[9]), .ZN(U_cr_n408) );
  AOI22_X2 U_cr_U204 ( .A1(U_cr_n424), .A2(U_cr_n563), .B1(U_cr_n423), .B2(
        cr_exn_mode_value[7]), .ZN(U_cr_n399) );
  OAI222_X2 U_cr_U203 ( .A1(U_cr_n487), .A2(U_cr_n437), .B1(U_cr_n492), .B2(
        U_cr_n438), .C1(U_cr_n182), .C2(U_cr_n455), .ZN(cr_reg_data_out[15])
         );
  AOI22_X2 U_cr_U202 ( .A1(U_cr_n424), .A2(U_cr_n570), .B1(U_cr_n423), .B2(
        cr_exn_mode_value[0]), .ZN(U_cr_n322) );
  AOI22_X2 U_cr_U201 ( .A1(U_cr_n430), .A2(cr_t_rc[2]), .B1(U_cr_n429), .B2(
        U_cr_srefr[24]), .ZN(U_cr_n486) );
  AOI22_X2 U_cr_U200 ( .A1(U_cr_n424), .A2(U_cr_n569), .B1(U_cr_n423), .B2(
        cr_exn_mode_value[1]), .ZN(U_cr_n425) );
  NOR2_X2 U_cr_U199 ( .A1(U_cr_n544), .A2(U_cr_n391), .ZN(U_cr_n232) );
  AOI22_X2 U_cr_U198 ( .A1(U_cr_n424), .A2(U_cr_n564), .B1(U_cr_n423), .B2(
        cr_exn_mode_value[6]), .ZN(U_cr_n386) );
  NOR2_X1 U_cr_U197 ( .A1(U_cr_n192), .A2(U_cr_n24), .ZN(U_cr_n201) );
  NAND3_X1 U_cr_U196 ( .A1(U_cr_n23), .A2(U_cr_cr_cs_0_), .A3(U_cr_cr_cs_2_), 
        .ZN(U_cr_n197) );
  INV_X4 U_cr_U194 ( .A(U_cr_n242), .ZN(U_cr_n168) );
  NOR2_X2 U_cr_U193 ( .A1(U_cr_n526), .A2(U_cr_n391), .ZN(U_cr_n230) );
  NOR2_X2 U_cr_U192 ( .A1(U_cr_n526), .A2(U_cr_n334), .ZN(U_cr_n313) );
  NOR2_X2 U_cr_U191 ( .A1(U_cr_n526), .A2(U_cr_n543), .ZN(U_cr_n536) );
  NOR2_X2 U_cr_U190 ( .A1(U_cr_n526), .A2(U_cr_n358), .ZN(U_cr_n305) );
  NOR2_X2 U_cr_U189 ( .A1(U_cr_n526), .A2(U_cr_n170), .ZN(U_cr_n289) );
  NOR2_X2 U_cr_U188 ( .A1(U_cr_n526), .A2(U_cr_n25), .ZN(U_cr_n268) );
  NAND2_X2 U_cr_U187 ( .A1(U_cr_n217), .A2(U_cr_n216), .ZN(U_cr_n544) );
  AOI22_X2 U_cr_U186 ( .A1(U_cr_n422), .A2(cr_mode_reg_update), .B1(U_cr_n407), 
        .B2(n[26]), .ZN(U_cr_n409) );
  NOR2_X2 U_cr_U185 ( .A1(U_cr_n544), .A2(U_cr_n170), .ZN(U_cr_n294) );
  NOR2_X2 U_cr_U184 ( .A1(U_cr_n544), .A2(U_cr_n25), .ZN(U_cr_n270) );
  NOR2_X2 U_cr_U183 ( .A1(U_cr_cr_cs_0_), .A2(U_cr_cr_cs_2_), .ZN(U_cr_n194)
         );
  NOR2_X2 U_cr_U182 ( .A1(U_cr_n178), .A2(U_cr_n23), .ZN(U_cr_n193) );
  NAND2_X1 U_cr_U181 ( .A1(U_cr_cr_cs_2_), .A2(U_cr_n16), .ZN(U_cr_n503) );
  NAND2_X2 U_cr_U180 ( .A1(U_cr_n217), .A2(U_cr_n213), .ZN(U_cr_n526) );
  NAND2_X1 U_cr_U179 ( .A1(n27), .A2(big_endian), .ZN(U_cr_n242) );
  NOR2_X2 U_cr_U178 ( .A1(U_cr_n320), .A2(U_cr_n263), .ZN(U_cr_n422) );
  AOI222_X1 U_cr_U177 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[13]), .B1(
        U_cr_n168), .B2(hiu_wr_data[21]), .C1(hiu_wr_data[5]), .C2(U_cr_n319), 
        .ZN(U_cr_n290) );
  AOI222_X1 U_cr_U176 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[12]), .B1(
        U_cr_n168), .B2(hiu_wr_data[20]), .C1(hiu_wr_data[4]), .C2(U_cr_n319), 
        .ZN(U_cr_n314) );
  AOI222_X1 U_cr_U175 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[11]), .B1(
        U_cr_n168), .B2(hiu_wr_data[19]), .C1(hiu_wr_data[3]), .C2(U_cr_n319), 
        .ZN(U_cr_n541) );
  AOI222_X1 U_cr_U174 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[15]), .B1(
        U_cr_n168), .B2(hiu_wr_data[23]), .C1(hiu_wr_data[7]), .C2(U_cr_n319), 
        .ZN(U_cr_n293) );
  AOI222_X1 U_cr_U173 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[14]), .B1(
        U_cr_n168), .B2(hiu_wr_data[22]), .C1(hiu_wr_data[6]), .C2(U_cr_n319), 
        .ZN(U_cr_n291) );
  AOI222_X1 U_cr_U172 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[1]), .B1(U_cr_n168), .B2(hiu_wr_data[25]), .C1(hiu_wr_data[9]), .C2(U_cr_n319), .ZN(U_cr_n516) );
  AOI222_X1 U_cr_U171 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[0]), .B1(U_cr_n168), .B2(hiu_wr_data[24]), .C1(hiu_wr_data[8]), .C2(U_cr_n319), .ZN(U_cr_n514) );
  NOR2_X2 U_cr_U170 ( .A1(U_cr_cr_cs_2_), .A2(U_cr_cr_cs_1_), .ZN(U_cr_n190)
         );
  MUX2_X1 U_cr_U168 ( .A(cr_s_data_width_early_0_), .B(n27), .S(U_cr_n197), 
        .Z(U_cr_n95) );
  NAND2_X2 U_cr_U167 ( .A1(U_cr_n191), .A2(U_cr_n24), .ZN(U_cr_n200) );
  INV_X1 U_cr_U166 ( .A(U_cr_n191), .ZN(U_cr_n192) );
  OAI21_X1 U_cr_U165 ( .B1(U_cr_sctlr_14_), .B2(U_cr_n206), .A(U_cr_n208), 
        .ZN(U_cr_n207) );
  INV_X2 U_cr_U164 ( .A(U_cr_n208), .ZN(U_cr_n209) );
  INV_X2 U_cr_U162 ( .A(U_cr_n207), .ZN(U_cr_N572) );
  NAND2_X1 U_cr_U161 ( .A1(U_cr_n193), .A2(U_cr_n319), .ZN(U_cr_n179) );
  NAND2_X1 U_cr_U160 ( .A1(hiu_haddr[2]), .A2(hiu_addr[6]), .ZN(U_cr_n360) );
  INV_X2 U_cr_U159 ( .A(hiu_haddr[3]), .ZN(U_cr_n283) );
  NOR2_X1 U_cr_U158 ( .A1(hiu_addr[5]), .A2(hiu_addr[7]), .ZN(U_cr_n284) );
  NOR2_X1 U_cr_U157 ( .A1(hiu_addr[6]), .A2(hiu_addr[4]), .ZN(U_cr_n300) );
  INV_X2 U_cr_U156 ( .A(hiu_haddr[2]), .ZN(U_cr_n320) );
  INV_X1 U_cr_U155 ( .A(hiu_addr[6]), .ZN(U_cr_n316) );
  NAND3_X1 U_cr_U154 ( .A1(hiu_addr[5]), .A2(hiu_addr[7]), .A3(hiu_addr[4]), 
        .ZN(U_cr_n359) );
  NAND4_X1 U_cr_U153 ( .A1(hiu_haddr[3]), .A2(hiu_addr[5]), .A3(hiu_addr[7]), 
        .A4(U_cr_n300), .ZN(U_cr_n308) );
  NOR2_X1 U_cr_U152 ( .A1(U_cr_n416), .A2(U_cr_n21), .ZN(U_cr_n383) );
  NOR2_X1 U_cr_U151 ( .A1(U_cr_n416), .A2(U_cr_n36), .ZN(U_cr_n351) );
  NAND3_X1 U_cr_U150 ( .A1(U_cr_n550), .A2(U_cr_n190), .A3(U_cr_cr_cs_0_), 
        .ZN(U_cr_n196) );
  AOI22_X1 U_cr_U149 ( .A1(U_cr_n407), .A2(U_cr_s_sda_d1), .B1(U_cr_n429), 
        .B2(gpo[3]), .ZN(U_cr_n353) );
  INV_X2 U_cr_U148 ( .A(U_cr_n412), .ZN(U_cr_n377) );
  AOI22_X1 U_cr_U147 ( .A1(U_cr_n407), .A2(cr_row_addr_width[2]), .B1(
        U_cr_n525), .B2(cr_block_size1[7]), .ZN(U_cr_n401) );
  OAI22_X1 U_cr_U146 ( .A1(U_cr_n318), .A2(U_cr_n200), .B1(U_cr_cr_cs_1_), 
        .B2(U_cr_n503), .ZN(U_cr_n222) );
  AOI21_X1 U_cr_U145 ( .B1(hiu_reg_req), .B2(U_cr_n504), .A(U_cr_cr_cs_0_), 
        .ZN(U_cr_n505) );
  AOI22_X1 U_cr_U144 ( .A1(U_cr_n424), .A2(U_cr_n565), .B1(U_cr_n171), .B2(
        cr_t_init[5]), .ZN(U_cr_n380) );
  AOI22_X1 U_cr_U143 ( .A1(U_cr_n430), .A2(cr_t_rcd[0]), .B1(U_cr_n171), .B2(
        cr_t_init[6]), .ZN(U_cr_n388) );
  OAI21_X2 U_cr_U142 ( .B1(U_cr_n200), .B2(U_cr_n317), .A(U_cr_n17), .ZN(
        U_cr_n217) );
  NAND4_X1 U_cr_U141 ( .A1(U_cr_n196), .A2(U_cr_n205), .A3(U_cr_n198), .A4(
        U_cr_n195), .ZN(U_cr_n96) );
  AOI22_X1 U_cr_U140 ( .A1(U_cr_n430), .A2(cr_t_rcd[1]), .B1(U_cr_n171), .B2(
        cr_t_init[7]), .ZN(U_cr_n400) );
  OAI21_X1 U_cr_U139 ( .B1(U_cr_n505), .B2(U_cr_n199), .A(U_cr_n198), .ZN(
        U_cr_n98) );
  INV_X2 U_cr_U138 ( .A(U_cr_n484), .ZN(U_cr_n403) );
  INV_X1 U_cr_U137 ( .A(U_cr_n188), .ZN(U_cr_n189) );
  AOI22_X1 U_cr_U136 ( .A1(U_cr_n430), .A2(cr_t_rcar[1]), .B1(U_cr_n171), .B2(
        cr_t_init[15]), .ZN(U_cr_n404) );
  AOI22_X1 U_cr_U135 ( .A1(U_cr_n430), .A2(cr_t_rcar[0]), .B1(U_cr_n171), .B2(
        cr_t_init[14]), .ZN(U_cr_n394) );
  AND2_X2 U_cr_U134 ( .A1(U_cr_n222), .A2(U_cr_n17), .ZN(U_cr_n238) );
  AOI21_X1 U_cr_U133 ( .B1(cr_do_self_ref_rp), .B2(U_cr_n422), .A(U_cr_n421), 
        .ZN(U_cr_n426) );
  AOI22_X1 U_cr_U132 ( .A1(U_cr_n424), .A2(U_cr_n567), .B1(U_cr_n171), .B2(
        cr_t_init[3]), .ZN(U_cr_n348) );
  NOR2_X1 U_cr_U131 ( .A1(U_cr_n334), .A2(U_cr_n37), .ZN(U_cr_n335) );
  AOI22_X1 U_cr_U130 ( .A1(U_cr_n430), .A2(cr_t_wr[1]), .B1(U_cr_n171), .B2(
        cr_t_init[13]), .ZN(U_cr_n375) );
  NAND2_X1 U_cr_U129 ( .A1(U_cr_n317), .A2(U_addrdec_n40), .ZN(U_cr_n175) );
  AOI21_X1 U_cr_U128 ( .B1(cr_t_xsr[0]), .B2(U_cr_n430), .A(U_cr_n377), .ZN(
        U_cr_n332) );
  AOI22_X1 U_cr_U127 ( .A1(U_cr_n430), .A2(cr_t_ras_min[2]), .B1(U_cr_n171), 
        .B2(cr_t_init[4]), .ZN(U_cr_n363) );
  AOI22_X1 U_cr_U126 ( .A1(U_cr_n169), .A2(cr_t_ref[1]), .B1(U_cr_n525), .B2(
        U_cr_n557), .ZN(U_cr_n428) );
  AND2_X2 U_cr_U125 ( .A1(U_cr_n430), .A2(U_cr_stmg0r_26), .ZN(U_cr_n344) );
  AOI22_X1 U_cr_U124 ( .A1(U_cr_n430), .A2(U_cr_stmg0r_1_), .B1(U_cr_n171), 
        .B2(cr_t_init[1]), .ZN(U_cr_n427) );
  AOI22_X1 U_cr_U123 ( .A1(U_cr_n430), .A2(cr_t_xsr[6]), .B1(U_cr_n169), .B2(
        U_cr_srefr[29]), .ZN(U_cr_n373) );
  AOI22_X1 U_cr_U122 ( .A1(U_cr_n430), .A2(U_cr_stmg0r_0_), .B1(U_cr_n171), 
        .B2(cr_t_init[0]), .ZN(U_cr_n324) );
  AOI22_X1 U_cr_U121 ( .A1(U_cr_n430), .A2(cr_t_rp[0]), .B1(U_cr_n171), .B2(
        cr_t_init[9]), .ZN(U_cr_n410) );
  AOI21_X1 U_cr_U120 ( .B1(gpo[6]), .B2(U_cr_n169), .A(U_cr_n392), .ZN(
        U_cr_n390) );
  NAND2_X1 U_cr_U119 ( .A1(U_cr_n430), .A2(U_cr_n236), .ZN(U_cr_n237) );
  AOI22_X1 U_cr_U118 ( .A1(U_cr_n169), .A2(cr_t_ref[6]), .B1(U_cr_n525), .B2(
        cr_block_size1[6]), .ZN(U_cr_n389) );
  AOI22_X1 U_cr_U117 ( .A1(U_cr_n169), .A2(cr_t_ref[9]), .B1(U_cr_n525), .B2(
        U_cr_n552), .ZN(U_cr_n411) );
  AOI21_X1 U_cr_U116 ( .B1(cr_t_rcar[2]), .B2(U_cr_n430), .A(U_cr_n377), .ZN(
        U_cr_n327) );
  OAI211_X1 U_cr_U115 ( .C1(U_cr_n29), .C2(U_cr_n170), .A(U_cr_n413), .B(
        U_cr_n412), .ZN(U_cr_n414) );
  AOI22_X1 U_cr_U114 ( .A1(U_cr_n169), .A2(cr_t_ref[0]), .B1(U_cr_n525), .B2(
        U_cr_n558), .ZN(U_cr_n325) );
  AOI22_X1 U_cr_U113 ( .A1(U_cr_n169), .A2(cr_t_ref[5]), .B1(U_cr_n525), .B2(
        cr_block_size1[5]), .ZN(U_cr_n381) );
  OAI21_X1 U_cr_U112 ( .B1(U_cr_n189), .B2(U_cr_cr_cs_1_), .A(U_cr_n194), .ZN(
        cr_push_n) );
  AOI22_X1 U_cr_U111 ( .A1(U_cr_n169), .A2(cr_t_ref[3]), .B1(U_cr_n525), .B2(
        U_cr_n555), .ZN(U_cr_n349) );
  AOI22_X1 U_cr_U110 ( .A1(U_cr_n430), .A2(cr_t_xsr[5]), .B1(U_cr_n169), .B2(
        U_cr_srefr[28]), .ZN(U_cr_n357) );
  OAI211_X1 U_cr_U109 ( .C1(U_cr_n416), .C2(U_cr_n30), .A(U_cr_n332), .B(
        U_cr_n331), .ZN(U_cr_n333) );
  OAI211_X1 U_cr_U108 ( .C1(U_cr_n416), .C2(U_cr_n28), .A(U_cr_n327), .B(
        U_cr_n326), .ZN(U_cr_n328) );
  OAI211_X1 U_cr_U107 ( .C1(U_cr_n33), .C2(U_cr_n391), .A(U_cr_n355), .B(
        U_cr_n412), .ZN(U_cr_n356) );
  INV_X2 U_cr_U106 ( .A(U_cr_n459), .ZN(U_cr_n420) );
  INV_X2 U_cr_U105 ( .A(U_cr_n498), .ZN(U_cr_n440) );
  INV_X2 U_cr_U104 ( .A(U_cr_n465), .ZN(U_cr_n443) );
  INV_X2 U_cr_U103 ( .A(U_cr_n472), .ZN(U_cr_n444) );
  INV_X2 U_cr_U102 ( .A(U_cr_n495), .ZN(U_cr_n418) );
  INV_X2 U_cr_U101 ( .A(U_cr_n478), .ZN(U_cr_n435) );
  INV_X2 U_cr_U100 ( .A(U_cr_n476), .ZN(U_cr_n436) );
  INV_X2 U_cr_U99 ( .A(U_cr_n496), .ZN(U_cr_n441) );
  INV_X2 U_cr_U98 ( .A(U_cr_n490), .ZN(U_cr_n439) );
  INV_X2 U_cr_U97 ( .A(U_cr_n448), .ZN(U_cr_n419) );
  NAND2_X1 U_cr_U96 ( .A1(U_cr_n291), .A2(U_cr_n221), .ZN(U_cr_n219) );
  INV_X2 U_cr_U95 ( .A(U_cr_n475), .ZN(U_cr_n454) );
  INV_X1 U_cr_U94 ( .A(U_cr_n182), .ZN(U_cr_n181) );
  NAND2_X1 U_cr_U93 ( .A1(U_cr_n219), .A2(cr_s_data_width_early_0_), .ZN(
        U_cr_n218) );
  NOR2_X1 U_cr_U92 ( .A1(U_cr_n455), .A2(U_cr_n185), .ZN(cr_reg_data_out[31])
         );
  INV_X2 U_cr_U91 ( .A(U_cr_n452), .ZN(U_cr_n477) );
  INV_X2 U_cr_U90 ( .A(U_cr_n494), .ZN(U_cr_n417) );
  OAI22_X1 U_cr_U89 ( .A1(U_cr_n288), .A2(U_cr_n534), .B1(cr_t_ref[1]), .B2(
        U_cr_n289), .ZN(U_cr_n286) );
  NAND2_X1 U_cr_U88 ( .A1(hiu_wr_data[3]), .A2(U_cr_n259), .ZN(U_cr_n249) );
  OAI22_X1 U_cr_U87 ( .A1(U_cr_n312), .A2(U_cr_n537), .B1(U_cr_n570), .B2(
        U_cr_n313), .ZN(U_cr_n309) );
  NAND2_X1 U_cr_U86 ( .A1(hiu_wr_data[2]), .A2(U_cr_n259), .ZN(U_cr_n247) );
  OAI22_X1 U_cr_U85 ( .A1(U_cr_n229), .A2(U_cr_n532), .B1(cr_t_ras_min[0]), 
        .B2(U_cr_n230), .ZN(U_cr_n228) );
  OAI22_X1 U_cr_U84 ( .A1(U_cr_n312), .A2(U_cr_n534), .B1(U_cr_n569), .B2(
        U_cr_n313), .ZN(U_cr_n310) );
  NAND2_X1 U_cr_U83 ( .A1(hiu_wr_data[1]), .A2(U_cr_n259), .ZN(U_cr_n245) );
  OAI22_X1 U_cr_U82 ( .A1(U_cr_n267), .A2(U_cr_n532), .B1(cr_t_init[2]), .B2(
        U_cr_n268), .ZN(U_cr_n266) );
  NAND2_X1 U_cr_U81 ( .A1(hiu_wr_data[0]), .A2(U_cr_n259), .ZN(U_cr_n243) );
  OAI22_X1 U_cr_U80 ( .A1(U_cr_n267), .A2(U_cr_n534), .B1(cr_t_init[1]), .B2(
        U_cr_n268), .ZN(U_cr_n265) );
  OAI22_X1 U_cr_U79 ( .A1(U_cr_n267), .A2(U_cr_n537), .B1(cr_t_init[0]), .B2(
        U_cr_n268), .ZN(U_cr_n264) );
  OAI22_X1 U_cr_U78 ( .A1(U_cr_n312), .A2(U_cr_n532), .B1(U_cr_n568), .B2(
        U_cr_n313), .ZN(U_cr_n311) );
  INV_X2 U_cr_U77 ( .A(U_cr_n442), .ZN(U_cr_n184) );
  OAI22_X1 U_cr_U76 ( .A1(U_cr_n538), .A2(U_cr_n532), .B1(U_cr_n556), .B2(
        U_cr_n536), .ZN(U_cr_n533) );
  OAI22_X1 U_cr_U75 ( .A1(U_cr_n538), .A2(U_cr_n534), .B1(U_cr_n557), .B2(
        U_cr_n536), .ZN(U_cr_n535) );
  OAI22_X1 U_cr_U74 ( .A1(U_cr_n538), .A2(U_cr_n537), .B1(U_cr_n558), .B2(
        U_cr_n536), .ZN(U_cr_n539) );
  AND2_X2 U_cr_U73 ( .A1(U_cr_n13), .A2(U_cr_n482), .ZN(cr_reg_data_out[23])
         );
  OAI21_X1 U_cr_U72 ( .B1(U_cr_n290), .B2(U_cr_n219), .A(U_cr_n218), .ZN(
        U_cr_N308) );
  OAI22_X1 U_cr_U71 ( .A1(U_cr_n304), .A2(U_cr_n537), .B1(cr_exn_mode_value[0]), .B2(U_cr_n305), .ZN(U_cr_n301) );
  OAI22_X1 U_cr_U70 ( .A1(U_cr_n304), .A2(U_cr_n534), .B1(cr_exn_mode_value[1]), .B2(U_cr_n305), .ZN(U_cr_n302) );
  OAI22_X1 U_cr_U69 ( .A1(U_cr_n304), .A2(U_cr_n532), .B1(cr_exn_mode_value[2]), .B2(U_cr_n305), .ZN(U_cr_n303) );
  OAI22_X1 U_cr_U68 ( .A1(U_cr_n288), .A2(U_cr_n532), .B1(cr_t_ref[2]), .B2(
        U_cr_n289), .ZN(U_cr_n287) );
  OAI22_X1 U_cr_U67 ( .A1(U_cr_n288), .A2(U_cr_n537), .B1(cr_t_ref[0]), .B2(
        U_cr_n289), .ZN(U_cr_n285) );
  NAND2_X1 U_cr_U66 ( .A1(hiu_wr_data[7]), .A2(U_cr_n259), .ZN(U_cr_n260) );
  NAND2_X1 U_cr_U65 ( .A1(hiu_wr_data[4]), .A2(U_cr_n259), .ZN(U_cr_n251) );
  NAND2_X1 U_cr_U64 ( .A1(hiu_wr_data[5]), .A2(U_cr_n259), .ZN(U_cr_n253) );
  NAND2_X1 U_cr_U63 ( .A1(hiu_wr_data[6]), .A2(U_cr_n259), .ZN(U_cr_n255) );
  OAI22_X1 U_cr_U62 ( .A1(U_cr_n272), .A2(U_cr_n532), .B1(cr_do_power_down), 
        .B2(U_cr_n273), .ZN(U_cr_n271) );
  INV_X2 U_cr_U61 ( .A(U_cr_n264), .ZN(U_cr_N464) );
  OAI211_X1 U_cr_U60 ( .C1(U_cr_n314), .C2(U_cr_n262), .A(U_cr_n252), .B(
        U_cr_n251), .ZN(U_cr_N417) );
  NOR2_X1 U_cr_U59 ( .A1(U_cr_n184), .A2(U_cr_n185), .ZN(cr_reg_data_out[27])
         );
  INV_X2 U_cr_U58 ( .A(U_cr_n271), .ZN(U_cr_N552) );
  INV_X2 U_cr_U57 ( .A(U_cr_n310), .ZN(U_cr_N734) );
  OAI211_X1 U_cr_U56 ( .C1(U_cr_n541), .C2(U_cr_n262), .A(U_cr_n250), .B(
        U_cr_n249), .ZN(U_cr_N416) );
  INV_X2 U_cr_U55 ( .A(U_cr_n539), .ZN(U_cr_n87) );
  OAI211_X1 U_cr_U54 ( .C1(U_cr_n290), .C2(U_cr_n262), .A(U_cr_n254), .B(
        U_cr_n253), .ZN(U_cr_N418) );
  INV_X2 U_cr_U53 ( .A(U_cr_n265), .ZN(U_cr_N465) );
  INV_X2 U_cr_U52 ( .A(U_cr_n287), .ZN(U_cr_N634) );
  INV_X2 U_cr_U51 ( .A(U_cr_n303), .ZN(U_cr_N690) );
  OAI211_X1 U_cr_U50 ( .C1(U_cr_n291), .C2(U_cr_n262), .A(U_cr_n256), .B(
        U_cr_n255), .ZN(U_cr_N419) );
  INV_X2 U_cr_U49 ( .A(U_cr_n228), .ZN(U_cr_N391) );
  INV_X2 U_cr_U48 ( .A(U_cr_n266), .ZN(U_cr_N466) );
  INV_X2 U_cr_U47 ( .A(U_cr_n301), .ZN(U_cr_N688) );
  OAI211_X1 U_cr_U46 ( .C1(U_cr_n293), .C2(U_cr_n262), .A(U_cr_n261), .B(
        U_cr_n260), .ZN(U_cr_N420) );
  OAI211_X1 U_cr_U45 ( .C1(U_cr_n548), .C2(U_cr_n262), .A(U_cr_n244), .B(
        U_cr_n243), .ZN(U_cr_N413) );
  INV_X2 U_cr_U44 ( .A(U_cr_n535), .ZN(U_cr_n86) );
  INV_X2 U_cr_U43 ( .A(U_cr_n309), .ZN(U_cr_N733) );
  INV_X2 U_cr_U42 ( .A(U_cr_n311), .ZN(U_cr_N735) );
  INV_X2 U_cr_U41 ( .A(U_cr_n302), .ZN(U_cr_N689) );
  INV_X2 U_cr_U40 ( .A(U_cr_n533), .ZN(U_cr_n85) );
  OAI21_X1 U_cr_U39 ( .B1(U_cr_n456), .B2(U_cr_n492), .A(U_cr_n354), .ZN(
        cr_reg_data_out[11]) );
  OAI21_X1 U_cr_U38 ( .B1(U_cr_n484), .B2(U_cr_n487), .A(U_cr_n483), .ZN(
        cr_reg_data_out[7]) );
  OAI21_X1 U_cr_U37 ( .B1(U_cr_n493), .B2(U_cr_n492), .A(U_cr_n491), .ZN(
        cr_reg_data_out[8]) );
  OAI21_X1 U_cr_U36 ( .B1(U_cr_n450), .B2(U_cr_n487), .A(U_cr_n346), .ZN(
        cr_reg_data_out[10]) );
  NOR2_X1 U_cr_U35 ( .A1(U_cr_n23), .A2(U_cr_n16), .ZN(U_cr_n191) );
  AOI22_X1 U_cr_U34 ( .A1(U_cr_stmg0r_0_), .A2(U_cr_stmg0r_1_), .B1(U_cr_n43), 
        .B2(U_cr_n20), .ZN(U_cr_N576) );
  INV_X4 U_cr_U33 ( .A(U_cr_n194), .ZN(U_cr_n178) );
  NOR2_X1 U_cr_U32 ( .A1(U_cr_n201), .A2(U_cr_n193), .ZN(U_cr_n198) );
  NAND2_X1 U_cr_U31 ( .A1(U_cr_cr_cs_1_), .A2(hiu_rw), .ZN(U_cr_n502) );
  NOR2_X1 U_cr_U30 ( .A1(hiu_burst_size[4]), .A2(hiu_burst_size[2]), .ZN(
        U_cr_n211) );
  NAND2_X1 U_cr_U29 ( .A1(hiu_reg_req), .A2(hiu_rw), .ZN(U_cr_n188) );
  OR2_X2 U_cr_U28 ( .A1(n27), .A2(U_cr_n222), .ZN(U_cr_n240) );
  AOI22_X1 U_cr_U27 ( .A1(U_cr_n430), .A2(cr_t_rcar[3]), .B1(U_cr_n171), .B2(
        cr_num_init_ref[1]), .ZN(U_cr_n413) );
  AOI22_X1 U_cr_U26 ( .A1(U_cr_n407), .A2(s_sda_oe_n), .B1(U_cr_n169), .B2(
        gpo[4]), .ZN(U_cr_n355) );
  AOI22_X1 U_cr_U25 ( .A1(U_cr_n430), .A2(cr_t_rc[3]), .B1(U_cr_n169), .B2(
        U_cr_srefr[25]), .ZN(U_cr_n432) );
  OAI21_X1 U_cr_U24 ( .B1(U_cr_n391), .B2(U_cr_n64), .A(U_cr_n390), .ZN(
        U_cr_n476) );
  OAI21_X1 U_cr_U23 ( .B1(U_cr_n474), .B2(U_cr_n487), .A(U_cr_n385), .ZN(
        cr_reg_data_out[13]) );
  OAI21_X1 U_cr_U22 ( .B1(U_cr_n461), .B2(U_cr_n492), .A(U_cr_n460), .ZN(
        cr_reg_data_out[3]) );
  INV_X1 U_cr_U21 ( .A(U_cr_n13), .ZN(U_cr_n185) );
  AOI21_X1 U_cr_U20 ( .B1(U_cr_n193), .B2(U_cr_n17), .A(U_cr_n177), .ZN(
        U_cr_n13) );
  AOI211_X1 U_cr_U19 ( .C1(U_cr_n430), .C2(cr_t_xsr[7]), .A(U_cr_n12), .B(
        U_cr_n392), .ZN(U_cr_n452) );
  AND2_X1 U_cr_U18 ( .A1(U_cr_n169), .A2(U_cr_srefr[30]), .ZN(U_cr_n12) );
  NAND3_X1 U_cr_U17 ( .A1(U_cr_n202), .A2(U_cr_n10), .A3(U_cr_n11), .ZN(
        U_cr_n99) );
  NAND4_X1 U_cr_U16 ( .A1(U_cr_n23), .A2(U_cr_n16), .A3(U_cr_n17), .A4(
        hiu_reg_req), .ZN(U_cr_n11) );
  AOI21_X1 U_cr_U15 ( .B1(U_cr_n550), .B2(U_cr_n9), .A(U_cr_n201), .ZN(
        U_cr_n10) );
  INV_X1 U_cr_U14 ( .A(U_cr_n200), .ZN(U_cr_n9) );
  AOI21_X1 U_cr_U13 ( .B1(cr_t_ref[11]), .B2(U_cr_n169), .A(U_cr_n8), .ZN(
        U_cr_n456) );
  NAND4_X1 U_cr_U12 ( .A1(U_cr_n5), .A2(U_cr_n6), .A3(U_cr_n7), .A4(U_cr_n378), 
        .ZN(U_cr_n8) );
  AOI22_X1 U_cr_U11 ( .A1(n[24]), .A2(U_cr_n407), .B1(U_cr_sctlr_default_11), 
        .B2(U_cr_n422), .ZN(U_cr_n7) );
  AOI22_X1 U_cr_U10 ( .A1(U_cr_n171), .A2(cr_t_init[11]), .B1(U_cr_n430), .B2(
        cr_t_rp[2]), .ZN(U_cr_n6) );
  AOI22_X1 U_cr_U9 ( .A1(U_cr_n424), .A2(U_cr_n560), .B1(cr_exn_mode_value[11]), .B2(U_cr_n423), .ZN(U_cr_n5) );
  AOI222_X1 U_cr_U8 ( .A1(U_addrdec_n40), .A2(hiu_wr_data[2]), .B1(
        hiu_wr_data[26]), .B2(U_cr_n168), .C1(hiu_wr_data[10]), .C2(U_cr_n319), 
        .ZN(U_cr_n518) );
  AOI211_X1 U_cr_U7 ( .C1(U_cr_n169), .C2(cr_t_ref[8]), .A(U_cr_n392), .B(
        U_cr_n4), .ZN(U_cr_n493) );
  NAND3_X1 U_cr_U6 ( .A1(U_cr_n1), .A2(U_cr_n2), .A3(U_cr_n3), .ZN(U_cr_n4) );
  AOI222_X1 U_cr_U5 ( .A1(U_cr_n430), .A2(cr_t_rcd[2]), .B1(U_cr_n423), .B2(
        cr_exn_mode_value[8]), .C1(U_cr_n407), .C2(cr_row_addr_width[3]), .ZN(
        U_cr_n3) );
  AOI22_X1 U_cr_U4 ( .A1(U_cr_n422), .A2(s_read_pipe[2]), .B1(U_cr_n525), .B2(
        U_cr_n553), .ZN(U_cr_n2) );
  AOI22_X1 U_cr_U3 ( .A1(U_cr_n171), .A2(cr_t_init[8]), .B1(U_cr_n424), .B2(
        U_cr_n562), .ZN(U_cr_n1) );
  DFFR_X2 U_cr_smskr0_reg_8_ ( .D(U_cr_n94), .CK(hclk), .RN(hresetn), .Q(
        U_cr_n553), .QN(U_cr_n154) );
  DFFR_X2 U_cr_smskr0_reg_10_ ( .D(U_cr_n92), .CK(hclk), .RN(hresetn), .Q(
        U_cr_n551), .QN(U_cr_n153) );
  DFFR_X2 U_cr_cr_cs_reg_2_ ( .D(U_cr_n96), .CK(hclk), .RN(hresetn), .Q(
        U_cr_cr_cs_2_), .QN(U_cr_n24) );
  DFFR_X2 U_cr_cr_cs_reg_0_ ( .D(U_cr_n99), .CK(hclk), .RN(hresetn), .Q(
        U_cr_cr_cs_0_), .QN(U_cr_n16) );
  DFFR_X2 U_cr_cr_cs_reg_1_ ( .D(U_cr_n98), .CK(hclk), .RN(hresetn), .Q(
        U_cr_cr_cs_1_), .QN(U_cr_n23) );
  DFFR_X2 U_cr_open_banks_o_reg_4_ ( .D(U_cr_N574), .CK(hclk), .RN(hresetn), 
        .Q(cr_num_open_banks[4]) );
  DFFR_X2 U_cr_sctlr_reg_11_ ( .D(ctl_sd_in_sf_mode), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_sctlr_default_11) );
  DFFR_X2 U_cr_open_banks_o_reg_3_ ( .D(U_cr_N573), .CK(hclk), .RN(hresetn), 
        .Q(cr_num_open_banks[3]), .QN(n92) );
  DFFR_X2 U_cr_cas_latency_o_reg_2_ ( .D(U_cr_N577), .CK(hclk), .RN(hresetn), 
        .Q(s_cas_latency[2]), .QN(n91) );
  DFFR_X2 U_cr_open_banks_o_reg_2_ ( .D(U_cr_N572), .CK(hclk), .RN(hresetn), 
        .Q(cr_num_open_banks[2]) );
  DFFR_X2 U_cr_s_sda_d1_reg ( .D(U_cr_s_sda_d), .CK(hclk), .RN(hresetn), .Q(
        U_cr_s_sda_d1) );
  DFFR_X2 U_cr_cas_latency_o_reg_0_ ( .D(U_cr_n20), .CK(hclk), .RN(hresetn), 
        .Q(s_cas_latency[0]), .QN(n90) );
  DFFR_X2 U_cr_syflash_opcode_reg_10_ ( .D(U_cr_n90), .CK(hclk), .RN(hresetn), 
        .QN(U_cr_n37) );
  DFFS_X2 U_cr_srefr_reg_1_ ( .D(U_cr_n286), .CK(hclk), .SN(hresetn), .QN(
        cr_t_ref[1]) );
  DFFS_X2 U_cr_srefr_reg_0_ ( .D(U_cr_n285), .CK(hclk), .SN(hresetn), .Q(n87), 
        .QN(cr_t_ref[0]) );
  DFFR_X1 U_cr_srefr_reg_16_ ( .D(U_cr_N648), .CK(hclk), .RN(hresetn), .Q(
        gpo[0]), .QN(U_cr_n47) );
  DFFR_X1 U_cr_srefr_reg_17_ ( .D(U_cr_N649), .CK(hclk), .RN(hresetn), .Q(
        gpo[1]), .QN(U_cr_n29) );
  DFFR_X1 U_cr_srefr_reg_18_ ( .D(U_cr_N650), .CK(hclk), .RN(hresetn), .Q(
        gpo[2]), .QN(U_cr_n48) );
  DFFR_X1 U_cr_srefr_reg_19_ ( .D(U_cr_N651), .CK(hclk), .RN(hresetn), .Q(
        gpo[3]), .QN(U_cr_n49) );
  DFFR_X1 U_cr_srefr_reg_20_ ( .D(U_cr_N652), .CK(hclk), .RN(hresetn), .Q(
        gpo[4]), .QN(U_cr_n50) );
  DFFR_X1 U_cr_srefr_reg_21_ ( .D(U_cr_N653), .CK(hclk), .RN(hresetn), .Q(
        gpo[5]), .QN(U_cr_n19) );
  DFFR_X1 U_cr_srefr_reg_22_ ( .D(U_cr_N654), .CK(hclk), .RN(hresetn), .Q(
        gpo[6]), .QN(U_cr_n46) );
  DFFR_X1 U_cr_srefr_reg_23_ ( .D(U_cr_N655), .CK(hclk), .RN(hresetn), .Q(
        gpo[7]), .QN(U_cr_n51) );
  DFFR_X1 U_cr_sctlr_reg_18_ ( .D(U_cr_N567), .CK(hclk), .RN(hresetn), .Q(
        cr_exn_mode_reg_update) );
  DFFR_X1 U_cr_sctlr_reg_17_ ( .D(U_cr_N566), .CK(hclk), .RN(hresetn), .Q(
        cr_s_ready_valid) );
  DFFR_X1 U_cr_sctlr_reg_16_ ( .D(U_cr_N565), .CK(hclk), .RN(hresetn), .Q(
        U_cr_sctlr_16_) );
  DFFR_X1 U_cr_sctlr_reg_19_ ( .D(U_cr_n73), .CK(hclk), .RN(hresetn), .Q(
        U_cr_n572) );
  DFFS_X2 U_cr_stmg1r_reg_16_ ( .D(U_cr_n74), .CK(hclk), .SN(hresetn), .Q(
        cr_num_init_ref[0]), .QN(U_cr_n115) );
  DFFS_X2 U_cr_stmg1r_reg_17_ ( .D(U_cr_n75), .CK(hclk), .SN(hresetn), .Q(
        cr_num_init_ref[1]), .QN(U_cr_n117) );
  DFFS_X2 U_cr_stmg1r_reg_18_ ( .D(U_cr_n76), .CK(hclk), .SN(hresetn), .Q(
        cr_num_init_ref[2]), .QN(U_cr_n116) );
  DFFR_X1 U_cr_stmg1r_reg_19_ ( .D(U_cr_n77), .CK(hclk), .RN(hresetn), .Q(
        cr_num_init_ref[3]), .QN(U_cr_n109) );
  DFFR_X1 U_cr_stmg1r_reg_20_ ( .D(U_cr_n78), .CK(hclk), .RN(hresetn), .Q(
        cr_t_wtr[0]), .QN(U_cr_n53) );
  DFFR_X1 U_cr_stmg1r_reg_21_ ( .D(U_cr_n79), .CK(hclk), .RN(hresetn), .Q(
        cr_t_wtr[1]), .QN(U_cr_n60) );
  DFFS_X2 U_cr_stmg0r_reg_24_ ( .D(U_cr_N413), .CK(hclk), .SN(hresetn), .Q(
        cr_t_rc[2]), .QN(n96) );
  DFFR_X1 U_cr_stmg0r_reg_25_ ( .D(U_cr_N414), .CK(hclk), .RN(hresetn), .Q(
        cr_t_rc[3]) );
  DFFR_X1 U_cr_stmg0r_reg_26_ ( .D(U_cr_N415), .CK(hclk), .RN(hresetn), .Q(
        U_cr_stmg0r_26) );
  DFFR_X1 U_cr_stmg0r_reg_27_ ( .D(U_cr_N416), .CK(hclk), .RN(hresetn), .Q(
        cr_t_xsr[4]) );
  DFFR_X1 U_cr_stmg0r_reg_28_ ( .D(U_cr_N417), .CK(hclk), .RN(hresetn), .Q(
        cr_t_xsr[5]) );
  DFFR_X1 U_cr_stmg0r_reg_29_ ( .D(U_cr_N418), .CK(hclk), .RN(hresetn), .Q(
        cr_t_xsr[6]) );
  DFFR_X1 U_cr_stmg0r_reg_30_ ( .D(U_cr_N419), .CK(hclk), .RN(hresetn), .Q(
        cr_t_xsr[7]) );
  DFFR_X1 U_cr_stmg0r_reg_31_ ( .D(U_cr_N420), .CK(hclk), .RN(hresetn), .Q(
        cr_t_xsr[8]) );
  DFFS_X2 U_cr_stmg0r_reg_16_ ( .D(U_cr_N405), .CK(hclk), .SN(hresetn), .Q(
        cr_t_rcar[2]), .QN(U_cr_n104) );
  DFFR_X1 U_cr_stmg0r_reg_17_ ( .D(U_cr_N406), .CK(hclk), .RN(hresetn), .Q(
        cr_t_rcar[3]), .QN(U_cr_n72) );
  DFFR_X1 U_cr_stmg0r_reg_18_ ( .D(U_cr_N407), .CK(hclk), .RN(hresetn), .Q(
        cr_t_xsr[0]), .QN(U_cr_n108) );
  DFFS_X2 U_cr_stmg0r_reg_19_ ( .D(U_cr_N408), .CK(hclk), .SN(hresetn), .Q(
        cr_t_xsr[1]), .QN(U_cr_n32) );
  DFFR_X1 U_cr_stmg0r_reg_20_ ( .D(U_cr_N409), .CK(hclk), .RN(hresetn), .Q(
        cr_t_xsr[2]), .QN(U_cr_n33) );
  DFFS_X2 U_cr_stmg0r_reg_21_ ( .D(U_cr_N410), .CK(hclk), .SN(hresetn), .Q(
        cr_t_xsr[3]), .QN(U_cr_n34) );
  DFFR_X1 U_cr_stmg0r_reg_22_ ( .D(U_cr_N411), .CK(hclk), .RN(hresetn), .QN(
        U_cr_n64) );
  DFFS_X2 U_cr_stmg0r_reg_23_ ( .D(U_cr_N412), .CK(hclk), .SN(hresetn), .Q(
        cr_t_rc[1]), .QN(U_cr_n106) );
  DFFR_X1 U_cr_sconr_reg_16_ ( .D(U_cr_N311), .CK(hclk), .RN(hresetn), .Q(
        s_sa[1]), .QN(U_cr_n28) );
  DFFR_X1 U_cr_sconr_reg_17_ ( .D(U_cr_N312), .CK(hclk), .RN(hresetn), .Q(
        s_sa[2]), .QN(U_cr_n31) );
  DFFS_X2 U_cr_sconr_reg_18_ ( .D(U_cr_N313), .CK(hclk), .SN(hresetn), .Q(
        s_scl), .QN(U_cr_n30) );
  DFFS_X2 U_cr_sconr_reg_19_ ( .D(U_cr_N314), .CK(hclk), .SN(hresetn), .Q(
        s_sda_out), .QN(U_cr_n62) );
  DFFS_X2 U_cr_sconr_reg_20_ ( .D(U_cr_N315), .CK(hclk), .SN(hresetn), .Q(
        s_sda_oe_n), .QN(U_cr_n57) );
  DFFR_X1 U_cr_exn_mode_reg_reg_7_ ( .D(U_cr_N695), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[7]), .QN(U_cr_n100) );
  DFFR_X1 U_cr_exn_mode_reg_reg_6_ ( .D(U_cr_N694), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[6]), .QN(U_cr_n125) );
  DFFR_X1 U_cr_exn_mode_reg_reg_5_ ( .D(U_cr_N693), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[5]), .QN(U_cr_n124) );
  DFFR_X1 U_cr_exn_mode_reg_reg_4_ ( .D(U_cr_N692), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[4]), .QN(U_cr_n26) );
  DFFR_X1 U_cr_exn_mode_reg_reg_3_ ( .D(U_cr_N691), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[3]), .QN(U_cr_n97) );
  DFFR_X1 U_cr_exn_mode_reg_reg_2_ ( .D(U_cr_N690), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[2]) );
  DFFR_X1 U_cr_exn_mode_reg_reg_1_ ( .D(U_cr_N689), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[1]) );
  DFFR_X1 U_cr_exn_mode_reg_reg_0_ ( .D(U_cr_N688), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[0]) );
  DFFR_X1 U_cr_smskr0_reg_7_ ( .D(U_cr_n80), .CK(hclk), .RN(hresetn), .Q(
        cr_block_size1[7]), .QN(U_cr_n167) );
  DFFR_X1 U_cr_smskr0_reg_6_ ( .D(U_cr_n81), .CK(hclk), .RN(hresetn), .Q(
        cr_block_size1[6]), .QN(U_cr_n119) );
  DFFR_X1 U_cr_smskr0_reg_5_ ( .D(U_cr_n82), .CK(hclk), .RN(hresetn), .Q(
        cr_block_size1[5]), .QN(U_cr_n110) );
  DFFR_X1 U_cr_smskr0_reg_4_ ( .D(U_cr_n83), .CK(hclk), .RN(hresetn), .Q(
        U_cr_n554), .QN(U_cr_n152) );
  DFFS_X2 U_cr_smskr0_reg_3_ ( .D(U_cr_n84), .CK(hclk), .SN(hresetn), .Q(
        U_cr_n555), .QN(U_cr_n165) );
  DFFS_X2 U_cr_smskr0_reg_2_ ( .D(U_cr_n85), .CK(hclk), .SN(hresetn), .Q(
        U_cr_n556) );
  DFFR_X1 U_cr_smskr0_reg_1_ ( .D(U_cr_n86), .CK(hclk), .RN(hresetn), .Q(
        U_cr_n557) );
  DFFS_X2 U_cr_smskr0_reg_0_ ( .D(U_cr_n87), .CK(hclk), .SN(hresetn), .Q(
        U_cr_n558) );
  DFFR_X1 U_cr_srefr_reg_7_ ( .D(U_cr_N639), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[7]), .QN(U_cr_n113) );
  DFFR_X1 U_cr_srefr_reg_6_ ( .D(U_cr_N638), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[6]), .QN(U_cr_n121) );
  DFFR_X1 U_cr_srefr_reg_5_ ( .D(U_cr_N637), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[5]), .QN(U_cr_n112) );
  DFFS_X2 U_cr_srefr_reg_4_ ( .D(U_cr_N636), .CK(hclk), .SN(hresetn), .Q(
        cr_t_ref[4]), .QN(U_cr_n130) );
  DFFR_X1 U_cr_srefr_reg_3_ ( .D(U_cr_N635), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[3]), .QN(U_cr_n69) );
  DFFR_X1 U_cr_srefr_reg_2_ ( .D(U_cr_N634), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[2]) );
  DFFS_X2 U_cr_sctlr_reg_7_ ( .D(U_cr_N557), .CK(hclk), .SN(hresetn), .Q(
        s_read_pipe[1]), .QN(U_cr_n59) );
  DFFR_X1 U_cr_sctlr_reg_6_ ( .D(U_cr_N556), .CK(hclk), .RN(hresetn), .Q(
        s_read_pipe[0]), .QN(U_cr_n40) );
  DFFR_X1 U_cr_sctlr_reg_5_ ( .D(U_cr_N555), .CK(hclk), .RN(hresetn), .Q(
        cr_ref_all_after_sr), .QN(U_cr_n132) );
  DFFR_X1 U_cr_sctlr_reg_4_ ( .D(U_cr_N554), .CK(hclk), .RN(hresetn), .Q(
        cr_ref_all_before_sr), .QN(U_cr_n139) );
  DFFS_X2 U_cr_sctlr_reg_3_ ( .D(U_cr_N553), .CK(hclk), .SN(hresetn), .Q(
        cr_delayed_precharge), .QN(U_cr_n58) );
  DFFR_X1 U_cr_sctlr_reg_2_ ( .D(U_cr_N552), .CK(hclk), .RN(hresetn), .Q(
        cr_do_power_down) );
  DFFR_X1 U_cr_sctlr_reg_1_ ( .D(U_cr_N551), .CK(hclk), .RN(hresetn), .Q(
        cr_do_self_ref_rp), .QN(U_cr_n39) );
  DFFS_X2 U_cr_sctlr_reg_0_ ( .D(U_cr_N550), .CK(hclk), .SN(hresetn), .Q(
        cr_do_initialize), .QN(U_cr_n56) );
  DFFR_X1 U_cr_stmg1r_reg_7_ ( .D(U_cr_N471), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[7]), .QN(U_cr_n142) );
  DFFR_X1 U_cr_stmg1r_reg_6_ ( .D(U_cr_N470), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[6]), .QN(U_cr_n135) );
  DFFR_X1 U_cr_stmg1r_reg_5_ ( .D(U_cr_N469), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[5]), .QN(U_cr_n141) );
  DFFR_X1 U_cr_stmg1r_reg_4_ ( .D(U_cr_N468), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[4]), .QN(U_cr_n134) );
  DFFS_X2 U_cr_stmg1r_reg_3_ ( .D(U_cr_N467), .CK(hclk), .SN(hresetn), .Q(
        cr_t_init[3]), .QN(U_cr_n150) );
  DFFR_X1 U_cr_stmg1r_reg_2_ ( .D(U_cr_N466), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[2]) );
  DFFR_X1 U_cr_stmg1r_reg_1_ ( .D(U_cr_N465), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[1]) );
  DFFR_X1 U_cr_stmg1r_reg_0_ ( .D(U_cr_N464), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[0]) );
  DFFR_X1 U_cr_stmg0r_reg_7_ ( .D(U_cr_N396), .CK(hclk), .RN(hresetn), .Q(
        cr_t_rcd[1]), .QN(U_cr_n133) );
  DFFS_X2 U_cr_stmg0r_reg_6_ ( .D(U_cr_N395), .CK(hclk), .SN(hresetn), .Q(
        cr_t_rcd[0]), .QN(U_cr_n149) );
  DFFR_X1 U_cr_stmg0r_reg_5_ ( .D(U_cr_N394), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ras_min[3]), .QN(U_cr_n54) );
  DFFS_X2 U_cr_stmg0r_reg_4_ ( .D(U_cr_N393), .CK(hclk), .SN(hresetn), .Q(
        cr_t_ras_min[2]), .QN(U_cr_n128) );
  DFFR_X1 U_cr_stmg0r_reg_3_ ( .D(U_cr_N392), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ras_min[1]), .QN(U_cr_n120) );
  DFFR_X1 U_cr_stmg0r_reg_2_ ( .D(U_cr_N391), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ras_min[0]), .QN(n95) );
  DFFS_X2 U_cr_cas_latency_o_reg_1_ ( .D(U_cr_N576), .CK(hclk), .SN(hresetn), 
        .Q(s_cas_latency[1]), .QN(n93) );
  DFFR_X1 U_cr_stmg0r_reg_1_ ( .D(U_cr_N390), .CK(hclk), .RN(hresetn), .Q(
        U_cr_stmg0r_1_), .QN(U_cr_n43) );
  DFFS_X2 U_cr_stmg0r_reg_0_ ( .D(U_cr_N389), .CK(hclk), .SN(hresetn), .Q(
        U_cr_stmg0r_0_), .QN(U_cr_n20) );
  DFFS_X2 U_cr_sconr_reg_7_ ( .D(U_cr_N302), .CK(hclk), .SN(hresetn), .Q(
        cr_row_addr_width[2]), .QN(U_cr_n55) );
  DFFR_X1 U_cr_sconr_reg_6_ ( .D(U_cr_N301), .CK(hclk), .RN(hresetn), .Q(
        cr_row_addr_width[1]), .QN(U_cr_n42) );
  DFFR_X1 U_cr_sconr_reg_5_ ( .D(U_cr_N300), .CK(hclk), .RN(hresetn), .Q(
        cr_row_addr_width[0]), .QN(U_cr_n21) );
  DFFR_X1 U_cr_sconr_reg_4_ ( .D(U_cr_N299), .CK(hclk), .RN(hresetn), .Q(
        cr_bank_addr_width[1]), .QN(U_cr_n66) );
  DFFS_X2 U_cr_sconr_reg_3_ ( .D(U_cr_N298), .CK(hclk), .SN(hresetn), .Q(
        cr_bank_addr_width[0]), .QN(U_cr_n36) );
  DFFR_X1 U_cr_syflash_opcode_reg_7_ ( .D(U_cr_N740), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n563), .QN(U_cr_n159) );
  DFFR_X1 U_cr_syflash_opcode_reg_6_ ( .D(U_cr_N739), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n564), .QN(U_cr_n158) );
  DFFR_X1 U_cr_syflash_opcode_reg_5_ ( .D(U_cr_N738), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n565), .QN(U_cr_n157) );
  DFFR_X1 U_cr_syflash_opcode_reg_4_ ( .D(U_cr_N737), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n566), .QN(U_cr_n164) );
  DFFR_X1 U_cr_syflash_opcode_reg_3_ ( .D(U_cr_N736), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n567), .QN(U_cr_n156) );
  DFFR_X1 U_cr_syflash_opcode_reg_2_ ( .D(U_cr_N735), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n568) );
  DFFR_X1 U_cr_syflash_opcode_reg_1_ ( .D(U_cr_N734), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n569) );
  DFFR_X1 U_cr_syflash_opcode_reg_0_ ( .D(U_cr_N733), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n570) );
  DFFR_X1 U_cr_syflash_opcode_reg_8_ ( .D(U_cr_n88), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n562), .QN(U_cr_n161) );
  DFFR_X1 U_cr_syflash_opcode_reg_9_ ( .D(U_cr_n89), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n561), .QN(U_cr_n162) );
  DFFR_X1 U_cr_syflash_opcode_reg_11_ ( .D(U_cr_n91), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n560), .QN(U_cr_n163) );
  DFFR_X1 U_cr_syflash_opcode_reg_12_ ( .D(U_cr_N745), .CK(hclk), .RN(hresetn), 
        .Q(U_cr_n571), .QN(U_cr_n160) );
  DFFR_X1 U_cr_exn_mode_reg_reg_12_ ( .D(U_cr_N700), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[12]), .QN(U_cr_n103) );
  DFFR_X1 U_cr_exn_mode_reg_reg_11_ ( .D(U_cr_N699), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[11]), .QN(U_cr_n102) );
  DFFR_X1 U_cr_exn_mode_reg_reg_10_ ( .D(U_cr_N698), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[10]), .QN(U_cr_n71) );
  DFFR_X1 U_cr_exn_mode_reg_reg_9_ ( .D(U_cr_N697), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[9]), .QN(U_cr_n101) );
  DFFR_X1 U_cr_exn_mode_reg_reg_8_ ( .D(U_cr_N696), .CK(hclk), .RN(hresetn), 
        .Q(cr_exn_mode_value[8]), .QN(U_cr_n126) );
  DFFS_X2 U_cr_smskr0_reg_9_ ( .D(U_cr_n93), .CK(hclk), .SN(hresetn), .Q(
        U_cr_n552), .QN(U_cr_n166) );
  DFFR_X1 U_cr_srefr_reg_15_ ( .D(U_cr_N647), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[15]), .QN(U_cr_n114) );
  DFFR_X1 U_cr_srefr_reg_14_ ( .D(U_cr_N646), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[14]), .QN(U_cr_n123) );
  DFFR_X1 U_cr_srefr_reg_13_ ( .D(U_cr_N645), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[13]), .QN(U_cr_n68) );
  DFFR_X1 U_cr_srefr_reg_12_ ( .D(U_cr_N644), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[12]), .QN(U_cr_n122) );
  DFFR_X1 U_cr_srefr_reg_11_ ( .D(U_cr_N643), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[11]), .QN(U_cr_n111) );
  DFFS_X2 U_cr_srefr_reg_10_ ( .D(U_cr_N642), .CK(hclk), .SN(hresetn), .Q(
        cr_t_ref[10]), .QN(U_cr_n129) );
  DFFR_X1 U_cr_srefr_reg_9_ ( .D(U_cr_N641), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[9]), .QN(U_cr_n105) );
  DFFR_X1 U_cr_srefr_reg_8_ ( .D(U_cr_N640), .CK(hclk), .RN(hresetn), .Q(
        cr_t_ref[8]), .QN(U_cr_n118) );
  DFFR_X1 U_cr_sctlr_reg_15_ ( .D(U_cr_N564), .CK(hclk), .RN(hresetn), .Q(
        U_cr_sctlr_15_), .QN(U_cr_n44) );
  DFFR_X1 U_cr_sctlr_reg_14_ ( .D(U_cr_N563), .CK(hclk), .RN(hresetn), .Q(
        U_cr_sctlr_14_), .QN(U_cr_n35) );
  DFFS_X2 U_cr_sctlr_reg_13_ ( .D(U_cr_N562), .CK(hclk), .SN(hresetn), .Q(
        U_cr_sctlr_13_), .QN(U_cr_n27) );
  DFFS_X2 U_cr_sctlr_reg_12_ ( .D(U_cr_N561), .CK(hclk), .SN(hresetn), .Q(
        U_cr_sctlr_12_), .QN(U_cr_n18) );
  DFFR_X1 U_cr_sctlr_reg_10_ ( .D(U_cr_N560), .CK(hclk), .RN(hresetn), .Q(
        U_cr_n559), .QN(U_cr_n155) );
  DFFR_X1 U_cr_sctlr_reg_9_ ( .D(U_cr_N559), .CK(hclk), .RN(hresetn), .Q(
        cr_mode_reg_update), .QN(U_cr_n61) );
  DFFR_X1 U_cr_sctlr_reg_8_ ( .D(U_cr_N558), .CK(hclk), .RN(hresetn), .Q(
        s_read_pipe[2]), .QN(U_cr_n41) );
  DFFR_X1 U_cr_stmg1r_reg_15_ ( .D(U_cr_N479), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[15]), .QN(U_cr_n146) );
  DFFR_X1 U_cr_stmg1r_reg_14_ ( .D(U_cr_N478), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[14]), .QN(U_cr_n138) );
  DFFR_X1 U_cr_stmg1r_reg_13_ ( .D(U_cr_N477), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[13]), .QN(U_cr_n145) );
  DFFR_X1 U_cr_stmg1r_reg_12_ ( .D(U_cr_N476), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[12]), .QN(U_cr_n131) );
  DFFR_X1 U_cr_stmg1r_reg_11_ ( .D(U_cr_N475), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[11]), .QN(U_cr_n144) );
  DFFR_X1 U_cr_stmg1r_reg_10_ ( .D(U_cr_N474), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[10]), .QN(U_cr_n137) );
  DFFR_X1 U_cr_stmg1r_reg_9_ ( .D(U_cr_N473), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[9]), .QN(U_cr_n143) );
  DFFR_X1 U_cr_stmg1r_reg_8_ ( .D(U_cr_N472), .CK(hclk), .RN(hresetn), .Q(
        cr_t_init[8]), .QN(U_cr_n136) );
  DFFS_X2 U_cr_stmg0r_reg_15_ ( .D(U_cr_N404), .CK(hclk), .SN(hresetn), .Q(
        cr_t_rcar[1]), .QN(U_cr_n151) );
  DFFS_X2 U_cr_stmg0r_reg_14_ ( .D(U_cr_N403), .CK(hclk), .SN(hresetn), .Q(
        cr_t_rcar[0]), .QN(U_cr_n127) );
  DFFR_X1 U_cr_stmg0r_reg_13_ ( .D(U_cr_N402), .CK(hclk), .RN(hresetn), .Q(
        cr_t_wr[1]), .QN(U_cr_n67) );
  DFFS_X2 U_cr_stmg0r_reg_12_ ( .D(U_cr_N401), .CK(hclk), .SN(hresetn), .Q(
        cr_t_wr[0]), .QN(U_cr_n107) );
  DFFR_X1 U_cr_stmg0r_reg_11_ ( .D(U_cr_N400), .CK(hclk), .RN(hresetn), .Q(
        cr_t_rp[2]), .QN(U_cr_n148) );
  DFFS_X2 U_cr_stmg0r_reg_10_ ( .D(U_cr_N399), .CK(hclk), .SN(hresetn), .Q(
        cr_t_rp[1]), .QN(U_cr_n147) );
  DFFR_X1 U_cr_stmg0r_reg_9_ ( .D(U_cr_N398), .CK(hclk), .RN(hresetn), .Q(
        cr_t_rp[0]), .QN(U_cr_n45) );
  DFFR_X1 U_cr_stmg0r_reg_8_ ( .D(U_cr_N397), .CK(hclk), .RN(hresetn), .Q(
        cr_t_rcd[2]), .QN(U_cr_n140) );
  DFFR_X1 U_cr_sconr_reg_15_ ( .D(U_cr_N310), .CK(hclk), .RN(hresetn), .Q(
        s_sa[0]), .QN(U_cr_n52) );
  DFFS_X2 U_cr_sdram_data_width_reg_0_ ( .D(U_cr_n95), .CK(hclk), .SN(hresetn), 
        .Q(n27), .QN(U_cr_n17) );
  DFFS_X2 U_cr_sconr_reg_13_ ( .D(U_cr_N308), .CK(hclk), .SN(hresetn), .Q(
        cr_s_data_width_early_0_), .QN(n85) );
  DFFS_X2 U_cr_sconr_reg_12_ ( .D(U_cr_N307), .CK(hclk), .SN(hresetn), .Q(
        n[23]), .QN(U_cr_n65) );
  DFFR_X1 U_cr_sconr_reg_11_ ( .D(U_cr_N306), .CK(hclk), .RN(hresetn), .Q(
        n[24]), .QN(U_cr_n38) );
  DFFS_X2 U_cr_sconr_reg_10_ ( .D(U_cr_N305), .CK(hclk), .SN(hresetn), .Q(
        n[25]), .QN(U_cr_n22) );
  DFFS_X2 U_cr_sconr_reg_9_ ( .D(U_cr_N304), .CK(hclk), .SN(hresetn), .Q(n[26]), .QN(U_cr_n63) );
  DFFS_X2 U_cr_sconr_reg_8_ ( .D(U_cr_N303), .CK(hclk), .SN(hresetn), .Q(
        cr_row_addr_width[3]), .QN(U_cr_n70) );
  DFFR_X1 U_cr_s_sda_d_reg ( .D(s_sda_in), .CK(hclk), .RN(hresetn), .Q(
        U_cr_s_sda_d) );
  DFFR_X1 U_cr_srefr_reg_24_ ( .D(gpi[0]), .CK(hclk), .RN(hresetn), .Q(
        U_cr_srefr[24]) );
  DFFR_X1 U_cr_srefr_reg_25_ ( .D(gpi[1]), .CK(hclk), .RN(hresetn), .Q(
        U_cr_srefr[25]) );
  DFFR_X1 U_cr_srefr_reg_26_ ( .D(gpi[2]), .CK(hclk), .RN(hresetn), .Q(
        U_cr_srefr[26]) );
  DFFR_X1 U_cr_srefr_reg_27_ ( .D(gpi[3]), .CK(hclk), .RN(hresetn), .Q(
        U_cr_srefr[27]) );
  DFFR_X1 U_cr_srefr_reg_28_ ( .D(gpi[4]), .CK(hclk), .RN(hresetn), .Q(
        U_cr_srefr[28]) );
  DFFR_X1 U_cr_srefr_reg_29_ ( .D(gpi[5]), .CK(hclk), .RN(hresetn), .Q(
        U_cr_srefr[29]) );
  DFFR_X1 U_cr_srefr_reg_30_ ( .D(gpi[6]), .CK(hclk), .RN(hresetn), .Q(
        U_cr_srefr[30]) );
  DFFR_X1 U_cr_srefr_reg_31_ ( .D(gpi[7]), .CK(hclk), .RN(hresetn), .Q(
        U_cr_srefr[31]) );
  DFFS_X2 U_cr_open_banks_o_reg_0_ ( .D(U_cr_n18), .CK(hclk), .SN(hresetn), 
        .Q(cr_num_open_banks[0]) );
  DFFS_X2 U_cr_open_banks_o_reg_1_ ( .D(U_cr_N571), .CK(hclk), .SN(hresetn), 
        .Q(cr_num_open_banks[1]) );
  NAND2_X2 U_addrdec_U359 ( .A1(U_addrdec_n16), .A2(U_addrdec_n21), .ZN(
        U_addrdec_n113) );
  NAND2_X2 U_addrdec_U358 ( .A1(U_addrdec_bcawp_2_), .A2(U_addrdec_bcawp_1_), 
        .ZN(U_addrdec_n105) );
  NAND2_X2 U_addrdec_U357 ( .A1(U_addrdec_n101), .A2(U_addrdec_bcawp_3_), .ZN(
        U_addrdec_n114) );
  MUX2_X2 U_addrdec_U356 ( .A(U_addrdec_n79), .B(debug_ad_col_addr_13_), .S(
        n[25]), .Z(U_addrdec_n84) );
  AND2_X4 U_addrdec_U355 ( .A1(U_addrdec_n253), .A2(
        U_addrdec_row_addr_mask[13]), .ZN(debug_ad_row_addr[13]) );
  OAI211_X2 U_addrdec_U354 ( .C1(n[23]), .C2(U_addrdec_n80), .A(U_addrdec_n78), 
        .B(U_addrdec_bank_addr_mask_1_), .ZN(U_addrdec_n94) );
  NOR2_X2 U_addrdec_U353 ( .A1(U_addrdec_n80), .A2(n[26]), .ZN(U_addrdec_n86)
         );
  AND2_X4 U_addrdec_U352 ( .A1(U_addrdec_n278), .A2(
        U_addrdec_row_addr_mask[15]), .ZN(debug_ad_row_addr[15]) );
  NAND2_X2 U_addrdec_U351 ( .A1(U_addrdec_n44), .A2(U_addrdec_n43), .ZN(
        debug_ad_col_addr_8_) );
  AND2_X4 U_addrdec_U350 ( .A1(hiu_addr[12]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n32) );
  NOR2_X2 U_addrdec_U349 ( .A1(U_addrdec_n117), .A2(U_addrdec_n113), .ZN(
        U_addrdec_n28) );
  AND2_X4 U_addrdec_U348 ( .A1(hiu_addr[13]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n27) );
  NOR2_X2 U_addrdec_U347 ( .A1(U_addrdec_n117), .A2(U_addrdec_n105), .ZN(
        U_addrdec_n26) );
  OR2_X4 U_addrdec_U346 ( .A1(U_addrdec_n114), .A2(U_addrdec_n105), .ZN(
        U_addrdec_n24) );
  OR2_X4 U_addrdec_U345 ( .A1(U_addrdec_n114), .A2(U_addrdec_n113), .ZN(
        U_addrdec_n23) );
  OR2_X4 U_addrdec_U344 ( .A1(U_addrdec_n117), .A2(U_addrdec_n115), .ZN(
        U_addrdec_n22) );
  NOR3_X2 U_addrdec_U343 ( .A1(U_addrdec_n106), .A2(U_addrdec_n105), .A3(
        U_addrdec_bcawp_3_), .ZN(U_addrdec_n18) );
  AND2_X4 U_addrdec_U342 ( .A1(U_addrdec_n104), .A2(U_addrdec_n103), .ZN(
        U_addrdec_n13) );
  NOR2_X2 U_addrdec_U341 ( .A1(U_addrdec_n114), .A2(U_addrdec_n115), .ZN(
        U_addrdec_n272) );
  NOR3_X2 U_addrdec_U340 ( .A1(U_addrdec_n67), .A2(n[23]), .A3(U_cr_n63), .ZN(
        U_addrdec_n74) );
  NOR2_X2 U_addrdec_U339 ( .A1(U_cr_n38), .A2(n[25]), .ZN(U_addrdec_n81) );
  NOR2_X2 U_addrdec_U338 ( .A1(U_addrdec_n91), .A2(U_addrdec_n90), .ZN(
        U_addrdec_n92) );
  AOI21_X2 U_addrdec_U337 ( .B1(U_addrdec_n59), .B2(n[26]), .A(U_addrdec_n57), 
        .ZN(U_addrdec_n73) );
  AOI22_X2 U_addrdec_U336 ( .A1(U_addrdec_n74), .A2(debug_ad_col_addr_8_), 
        .B1(debug_ad_col_addr_15_), .B2(U_addrdec_n75), .ZN(U_addrdec_n70) );
  AND2_X4 U_addrdec_U335 ( .A1(U_addrdec_n263), .A2(
        U_addrdec_row_addr_mask[14]), .ZN(debug_ad_row_addr[14]) );
  MUX2_X2 U_addrdec_U334 ( .A(ad_cr_data_mask[1]), .B(ad_cr_data_mask[3]), .S(
        U_addrdec_n304), .Z(ad_data_mask[1]) );
  MUX2_X2 U_addrdec_U333 ( .A(ad_cr_data_mask[0]), .B(ad_cr_data_mask[2]), .S(
        U_addrdec_n304), .Z(ad_data_mask[0]) );
  AOI22_X1 U_addrdec_U332 ( .A1(U_addrdec_n220), .A2(hiu_addr[8]), .B1(
        hiu_addr[7]), .B2(U_addrdec_n39), .ZN(U_addrdec_n100) );
  XNOR2_X2 U_addrdec_U331 ( .A(cr_bank_addr_width[1]), .B(U_addrdec_n286), 
        .ZN(U_addrdec_N108) );
  NAND2_X2 U_addrdec_U329 ( .A1(U_addrdec_n15), .A2(U_addrdec_bcawp_0_), .ZN(
        U_addrdec_n106) );
  NAND2_X2 U_addrdec_U328 ( .A1(U_addrdec_n16), .A2(U_addrdec_bcawp_1_), .ZN(
        U_addrdec_n115) );
  INV_X4 U_addrdec_U325 ( .A(U_addrdec_n102), .ZN(U_addrdec_n180) );
  NAND3_X2 U_addrdec_U324 ( .A1(U_addrdec_n20), .A2(U_addrdec_n15), .A3(
        U_addrdec_bcawp_3_), .ZN(U_addrdec_n117) );
  NAND2_X2 U_addrdec_U323 ( .A1(U_addrdec_n21), .A2(U_addrdec_bcawp_2_), .ZN(
        U_addrdec_n116) );
  NOR2_X2 U_addrdec_U322 ( .A1(U_addrdec_n117), .A2(U_addrdec_n116), .ZN(
        U_addrdec_n17) );
  INV_X4 U_addrdec_U321 ( .A(U_addrdec_n17), .ZN(U_addrdec_n161) );
  OAI22_X2 U_addrdec_U320 ( .A1(U_addrdec_n180), .A2(U_addrdec_n161), .B1(
        U_addrdec_n13), .B2(U_addrdec_n130), .ZN(U_addrdec_n136) );
  NAND2_X2 U_addrdec_U319 ( .A1(hiu_addr[20]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n107) );
  NAND2_X2 U_addrdec_U318 ( .A1(U_addrdec_n108), .A2(U_addrdec_n107), .ZN(
        U_addrdec_n181) );
  INV_X4 U_addrdec_U317 ( .A(U_addrdec_n24), .ZN(U_addrdec_n35) );
  AOI22_X2 U_addrdec_U316 ( .A1(U_addrdec_n26), .A2(U_addrdec_n34), .B1(
        U_addrdec_n181), .B2(U_addrdec_n35), .ZN(U_addrdec_n134) );
  NAND2_X2 U_addrdec_U315 ( .A1(hiu_addr[22]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n132) );
  NAND2_X2 U_addrdec_U314 ( .A1(hiu_addr[21]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n131) );
  NAND2_X2 U_addrdec_U313 ( .A1(U_addrdec_n132), .A2(U_addrdec_n131), .ZN(
        U_addrdec_n232) );
  NAND2_X2 U_addrdec_U312 ( .A1(hiu_addr[20]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n122) );
  NAND2_X2 U_addrdec_U311 ( .A1(hiu_addr[21]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n121) );
  INV_X4 U_addrdec_U310 ( .A(U_addrdec_n25), .ZN(U_addrdec_n36) );
  AOI22_X2 U_addrdec_U309 ( .A1(U_addrdec_n30), .A2(U_addrdec_n232), .B1(
        U_addrdec_n219), .B2(U_addrdec_n36), .ZN(U_addrdec_n133) );
  NAND2_X2 U_addrdec_U308 ( .A1(U_addrdec_n134), .A2(U_addrdec_n133), .ZN(
        U_addrdec_n135) );
  AOI211_X2 U_addrdec_U307 ( .C1(U_addrdec_n272), .C2(debug_ad_col_addr_15_), 
        .A(U_addrdec_n136), .B(U_addrdec_n135), .ZN(U_addrdec_n139) );
  INV_X4 U_addrdec_U306 ( .A(debug_ad_col_addr_12_), .ZN(
        debug_ad_col_addr_12__BAR_BAR) );
  NAND2_X2 U_addrdec_U305 ( .A1(hiu_addr[12]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n54) );
  AOI22_X2 U_addrdec_U304 ( .A1(debug_ad_col_addr_12__BAR_BAR), .A2(
        U_addrdec_n28), .B1(debug_ad_col_addr_11_), .B2(U_addrdec_n18), .ZN(
        U_addrdec_n138) );
  INV_X4 U_addrdec_U303 ( .A(U_addrdec_n23), .ZN(U_addrdec_n37) );
  INV_X4 U_addrdec_U299 ( .A(U_addrdec_n22), .ZN(U_addrdec_n38) );
  AOI22_X2 U_addrdec_U298 ( .A1(debug_ad_col_addr_13__BAR_BAR), .A2(
        U_addrdec_n37), .B1(debug_ad_col_addr_14_), .B2(U_addrdec_n38), .ZN(
        U_addrdec_n137) );
  NAND3_X2 U_addrdec_U297 ( .A1(U_addrdec_n139), .A2(U_addrdec_n138), .A3(
        U_addrdec_n137), .ZN(debug_ad_row_addr[2]) );
  INV_X4 U_addrdec_U296 ( .A(hiu_mem_req), .ZN(U_addrdec_n310) );
  OAI22_X2 U_addrdec_U295 ( .A1(U_addrdec_n180), .A2(U_addrdec_n130), .B1(
        U_addrdec_n13), .B2(U_addrdec_n256), .ZN(U_addrdec_n126) );
  AOI22_X2 U_addrdec_U294 ( .A1(U_addrdec_n35), .A2(U_addrdec_n34), .B1(
        U_addrdec_n219), .B2(U_addrdec_n30), .ZN(U_addrdec_n124) );
  AOI22_X2 U_addrdec_U293 ( .A1(U_addrdec_n28), .A2(debug_ad_col_addr_11_), 
        .B1(U_addrdec_n181), .B2(U_addrdec_n36), .ZN(U_addrdec_n123) );
  NAND2_X2 U_addrdec_U292 ( .A1(U_addrdec_n124), .A2(U_addrdec_n123), .ZN(
        U_addrdec_n125) );
  AOI211_X2 U_addrdec_U291 ( .C1(U_addrdec_n17), .C2(debug_ad_col_addr_15_), 
        .A(U_addrdec_n126), .B(U_addrdec_n125), .ZN(U_addrdec_n129) );
  AOI22_X2 U_addrdec_U288 ( .A1(debug_ad_col_addr_12__BAR_BAR), .A2(
        U_addrdec_n37), .B1(debug_ad_col_addr_10_), .B2(U_addrdec_n18), .ZN(
        U_addrdec_n128) );
  AOI22_X2 U_addrdec_U287 ( .A1(debug_ad_col_addr_13__BAR_BAR), .A2(
        U_addrdec_n38), .B1(debug_ad_col_addr_14_), .B2(U_addrdec_n272), .ZN(
        U_addrdec_n127) );
  NAND3_X2 U_addrdec_U286 ( .A1(U_addrdec_n129), .A2(U_addrdec_n128), .A3(
        U_addrdec_n127), .ZN(debug_ad_row_addr[1]) );
  INV_X4 U_addrdec_U285 ( .A(debug_ad_col_addr_11_), .ZN(U_addrdec_n79) );
  NAND2_X2 U_addrdec_U282 ( .A1(n[24]), .A2(n[25]), .ZN(U_addrdec_n67) );
  NAND2_X2 U_addrdec_U280 ( .A1(debug_ad_col_addr_9_), .A2(U_addrdec_n74), 
        .ZN(U_addrdec_n77) );
  NAND2_X2 U_addrdec_U276 ( .A1(U_addrdec_n102), .A2(U_addrdec_n75), .ZN(
        U_addrdec_n76) );
  NAND2_X2 U_addrdec_U275 ( .A1(U_addrdec_n77), .A2(U_addrdec_n76), .ZN(
        U_addrdec_n80) );
  NOR2_X2 U_addrdec_U274 ( .A1(U_addrdec_n80), .A2(U_cr_n63), .ZN(
        U_addrdec_n83) );
  NAND2_X2 U_addrdec_U273 ( .A1(debug_ad_col_addr_15_), .A2(U_addrdec_n81), 
        .ZN(U_addrdec_n82) );
  INV_X4 U_addrdec_U272 ( .A(U_addrdec_n85), .ZN(U_addrdec_n93) );
  NAND2_X2 U_addrdec_U271 ( .A1(debug_ad_col_addr_14_), .A2(U_addrdec_n81), 
        .ZN(U_addrdec_n88) );
  NAND3_X2 U_addrdec_U270 ( .A1(U_addrdec_n86), .A2(n[24]), .A3(U_addrdec_n88), 
        .ZN(U_addrdec_n78) );
  NAND2_X2 U_addrdec_U269 ( .A1(debug_ad_col_addr_10_), .A2(U_cr_n22), .ZN(
        U_addrdec_n87) );
  OAI211_X2 U_addrdec_U268 ( .C1(debug_ad_col_addr_12_), .C2(U_cr_n22), .A(
        U_addrdec_n88), .B(U_addrdec_n87), .ZN(U_addrdec_n90) );
  NOR3_X2 U_addrdec_U267 ( .A1(U_addrdec_n93), .A2(U_addrdec_n94), .A3(
        U_addrdec_n92), .ZN(n44) );
  NOR3_X2 U_addrdec_U266 ( .A1(debug_ad_col_addr_13_), .A2(n[26]), .A3(
        U_addrdec_n56), .ZN(U_addrdec_n57) );
  NOR3_X2 U_addrdec_U265 ( .A1(debug_ad_col_addr_12__BAR_BAR), .A2(U_cr_n63), 
        .A3(U_cr_n22), .ZN(U_addrdec_n60) );
  NOR3_X2 U_addrdec_U264 ( .A1(U_addrdec_n60), .A2(n[24]), .A3(U_cr_n65), .ZN(
        U_addrdec_n66) );
  NAND3_X2 U_addrdec_U263 ( .A1(U_addrdec_n79), .A2(n[25]), .A3(U_cr_n63), 
        .ZN(U_addrdec_n65) );
  NAND3_X2 U_addrdec_U262 ( .A1(U_addrdec_n61), .A2(U_cr_n63), .A3(U_cr_n22), 
        .ZN(U_addrdec_n64) );
  NAND3_X2 U_addrdec_U261 ( .A1(U_addrdec_n62), .A2(n[26]), .A3(U_cr_n22), 
        .ZN(U_addrdec_n63) );
  NAND4_X2 U_addrdec_U260 ( .A1(U_addrdec_n66), .A2(U_addrdec_n65), .A3(
        U_addrdec_n64), .A4(U_addrdec_n63), .ZN(U_addrdec_n71) );
  NAND2_X2 U_addrdec_U259 ( .A1(hiu_addr[9]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n44) );
  NAND2_X2 U_addrdec_U258 ( .A1(hiu_addr[8]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n43) );
  NAND2_X2 U_addrdec_U257 ( .A1(hiu_addr[23]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n141) );
  NAND2_X2 U_addrdec_U256 ( .A1(hiu_addr[22]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n140) );
  NAND2_X2 U_addrdec_U255 ( .A1(U_addrdec_n141), .A2(U_addrdec_n140), .ZN(
        U_addrdec_n242) );
  AOI22_X2 U_addrdec_U254 ( .A1(U_addrdec_n18), .A2(U_addrdec_n219), .B1(
        U_addrdec_n242), .B2(U_addrdec_n37), .ZN(U_addrdec_n226) );
  NAND2_X2 U_addrdec_U253 ( .A1(hiu_addr[24]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n156) );
  NAND2_X2 U_addrdec_U252 ( .A1(hiu_addr[23]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n155) );
  NAND2_X2 U_addrdec_U251 ( .A1(U_addrdec_n156), .A2(U_addrdec_n155), .ZN(
        U_addrdec_n254) );
  NAND2_X2 U_addrdec_U250 ( .A1(hiu_addr[25]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n167) );
  NAND2_X2 U_addrdec_U249 ( .A1(hiu_addr[24]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n166) );
  NAND2_X2 U_addrdec_U248 ( .A1(U_addrdec_n167), .A2(U_addrdec_n166), .ZN(
        U_addrdec_n264) );
  AOI22_X2 U_addrdec_U247 ( .A1(U_addrdec_n38), .A2(U_addrdec_n254), .B1(
        U_addrdec_n264), .B2(U_addrdec_n272), .ZN(U_addrdec_n225) );
  NAND2_X2 U_addrdec_U246 ( .A1(U_addrdec_n222), .A2(U_addrdec_n221), .ZN(
        U_addrdec_n270) );
  AOI22_X2 U_addrdec_U245 ( .A1(U_addrdec_n232), .A2(U_addrdec_n28), .B1(
        U_addrdec_n270), .B2(U_addrdec_n30), .ZN(U_addrdec_n224) );
  NAND4_X2 U_addrdec_U244 ( .A1(U_addrdec_n226), .A2(U_addrdec_n225), .A3(
        U_addrdec_n224), .A4(U_addrdec_n223), .ZN(U_addrdec_n230) );
  NAND2_X2 U_addrdec_U243 ( .A1(hiu_addr[25]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n176) );
  NAND2_X2 U_addrdec_U242 ( .A1(U_addrdec_n176), .A2(U_addrdec_n175), .ZN(
        U_addrdec_n265) );
  NAND2_X2 U_addrdec_U241 ( .A1(U_addrdec_n196), .A2(U_addrdec_n195), .ZN(
        U_addrdec_n267) );
  AOI22_X2 U_addrdec_U240 ( .A1(U_addrdec_n17), .A2(U_addrdec_n265), .B1(
        U_addrdec_n267), .B2(U_addrdec_n26), .ZN(U_addrdec_n228) );
  NAND2_X2 U_addrdec_U239 ( .A1(U_addrdec_n206), .A2(U_addrdec_n205), .ZN(
        U_addrdec_n273) );
  NAND2_X2 U_addrdec_U238 ( .A1(U_addrdec_n187), .A2(U_addrdec_n186), .ZN(
        U_addrdec_n266) );
  AOI22_X2 U_addrdec_U237 ( .A1(U_addrdec_n35), .A2(U_addrdec_n273), .B1(
        U_addrdec_n266), .B2(U_addrdec_n269), .ZN(U_addrdec_n227) );
  NAND2_X2 U_addrdec_U236 ( .A1(U_addrdec_n228), .A2(U_addrdec_n227), .ZN(
        U_addrdec_n229) );
  OAI21_X2 U_addrdec_U235 ( .B1(U_addrdec_n230), .B2(U_addrdec_n229), .A(
        U_addrdec_row_addr_mask[11]), .ZN(U_addrdec_n231) );
  INV_X4 U_addrdec_U234 ( .A(U_addrdec_n231), .ZN(debug_ad_row_addr[11]) );
  INV_X4 U_addrdec_U233 ( .A(U_addrdec_n18), .ZN(U_addrdec_n245) );
  INV_X4 U_addrdec_U232 ( .A(U_addrdec_n181), .ZN(U_addrdec_n210) );
  INV_X4 U_addrdec_U231 ( .A(U_addrdec_n28), .ZN(U_addrdec_n243) );
  OAI22_X2 U_addrdec_U230 ( .A1(U_addrdec_n200), .A2(U_addrdec_n245), .B1(
        U_addrdec_n210), .B2(U_addrdec_n243), .ZN(U_addrdec_n204) );
  AOI22_X2 U_addrdec_U229 ( .A1(U_addrdec_n37), .A2(U_addrdec_n219), .B1(
        U_addrdec_n242), .B2(U_addrdec_n272), .ZN(U_addrdec_n202) );
  AOI22_X2 U_addrdec_U228 ( .A1(U_addrdec_n38), .A2(U_addrdec_n232), .B1(
        U_addrdec_n254), .B2(U_addrdec_n17), .ZN(U_addrdec_n201) );
  NAND2_X2 U_addrdec_U227 ( .A1(U_addrdec_n202), .A2(U_addrdec_n201), .ZN(
        U_addrdec_n203) );
  AOI211_X2 U_addrdec_U226 ( .C1(U_addrdec_n36), .C2(U_addrdec_n267), .A(
        U_addrdec_n204), .B(U_addrdec_n203), .ZN(U_addrdec_n209) );
  AOI22_X2 U_addrdec_U225 ( .A1(U_addrdec_n26), .A2(U_addrdec_n265), .B1(
        U_addrdec_n264), .B2(U_addrdec_n269), .ZN(U_addrdec_n208) );
  AOI22_X2 U_addrdec_U224 ( .A1(U_addrdec_n30), .A2(U_addrdec_n273), .B1(
        U_addrdec_n266), .B2(U_addrdec_n35), .ZN(U_addrdec_n207) );
  NAND3_X2 U_addrdec_U223 ( .A1(U_addrdec_n209), .A2(U_addrdec_n208), .A3(
        U_addrdec_n207), .ZN(debug_ad_row_addr[9]) );
  OAI22_X2 U_addrdec_U222 ( .A1(U_addrdec_n180), .A2(U_addrdec_n23), .B1(
        U_addrdec_n210), .B2(U_addrdec_n161), .ZN(U_addrdec_n165) );
  AOI22_X2 U_addrdec_U221 ( .A1(U_addrdec_n26), .A2(U_addrdec_n232), .B1(
        U_addrdec_n219), .B2(U_addrdec_n269), .ZN(U_addrdec_n163) );
  OAI211_X2 U_addrdec_U220 ( .C1(U_addrdec_n13), .C2(U_addrdec_n22), .A(
        U_addrdec_n163), .B(U_addrdec_n162), .ZN(U_addrdec_n164) );
  AOI22_X2 U_addrdec_U219 ( .A1(U_addrdec_n35), .A2(U_addrdec_n242), .B1(
        U_addrdec_n264), .B2(U_addrdec_n30), .ZN(U_addrdec_n169) );
  AOI22_X2 U_addrdec_U218 ( .A1(U_addrdec_n28), .A2(debug_ad_col_addr_15_), 
        .B1(U_addrdec_n254), .B2(U_addrdec_n36), .ZN(U_addrdec_n168) );
  NAND3_X2 U_addrdec_U217 ( .A1(U_addrdec_n170), .A2(U_addrdec_n169), .A3(
        U_addrdec_n168), .ZN(debug_ad_row_addr[5]) );
  AOI22_X2 U_addrdec_U216 ( .A1(U_addrdec_n28), .A2(U_addrdec_n265), .B1(
        U_addrdec_n264), .B2(U_addrdec_n18), .ZN(U_addrdec_n277) );
  AOI22_X2 U_addrdec_U215 ( .A1(U_addrdec_n38), .A2(U_addrdec_n267), .B1(
        U_addrdec_n266), .B2(U_addrdec_n37), .ZN(U_addrdec_n276) );
  NAND2_X2 U_addrdec_U214 ( .A1(hiu_addr[31]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n255) );
  AOI22_X2 U_addrdec_U213 ( .A1(U_addrdec_n270), .A2(U_addrdec_n269), .B1(
        U_addrdec_n268), .B2(U_addrdec_n26), .ZN(U_addrdec_n275) );
  AOI22_X2 U_addrdec_U212 ( .A1(U_addrdec_n273), .A2(U_addrdec_n272), .B1(
        U_addrdec_n271), .B2(U_addrdec_n17), .ZN(U_addrdec_n274) );
  NAND4_X2 U_addrdec_U211 ( .A1(U_addrdec_n277), .A2(U_addrdec_n276), .A3(
        U_addrdec_n275), .A4(U_addrdec_n274), .ZN(U_addrdec_n278) );
  NOR2_X2 U_addrdec_U210 ( .A1(U_addrdec_n255), .A2(U_addrdec_n25), .ZN(
        U_addrdec_n248) );
  OAI22_X2 U_addrdec_U209 ( .A1(U_addrdec_n246), .A2(U_addrdec_n245), .B1(
        U_addrdec_n244), .B2(U_addrdec_n243), .ZN(U_addrdec_n247) );
  AOI211_X2 U_addrdec_U208 ( .C1(U_addrdec_n35), .C2(U_addrdec_n270), .A(
        U_addrdec_n248), .B(U_addrdec_n247), .ZN(U_addrdec_n252) );
  AOI22_X2 U_addrdec_U207 ( .A1(U_addrdec_n272), .A2(U_addrdec_n266), .B1(
        U_addrdec_n264), .B2(U_addrdec_n37), .ZN(U_addrdec_n251) );
  AOI22_X2 U_addrdec_U206 ( .A1(U_addrdec_n38), .A2(U_addrdec_n265), .B1(
        U_addrdec_n273), .B2(U_addrdec_n269), .ZN(U_addrdec_n250) );
  AOI22_X2 U_addrdec_U205 ( .A1(U_addrdec_n267), .A2(U_addrdec_n17), .B1(
        U_addrdec_n271), .B2(U_addrdec_n26), .ZN(U_addrdec_n249) );
  NAND4_X2 U_addrdec_U204 ( .A1(U_addrdec_n252), .A2(U_addrdec_n251), .A3(
        U_addrdec_n250), .A4(U_addrdec_n249), .ZN(U_addrdec_n253) );
  OAI22_X2 U_addrdec_U203 ( .A1(U_addrdec_n180), .A2(U_addrdec_n245), .B1(
        U_addrdec_n13), .B2(U_addrdec_n243), .ZN(U_addrdec_n185) );
  AOI22_X2 U_addrdec_U202 ( .A1(U_addrdec_n38), .A2(U_addrdec_n181), .B1(
        U_addrdec_n219), .B2(U_addrdec_n272), .ZN(U_addrdec_n183) );
  AOI22_X2 U_addrdec_U201 ( .A1(U_addrdec_n17), .A2(U_addrdec_n232), .B1(
        U_addrdec_n34), .B2(U_addrdec_n37), .ZN(U_addrdec_n182) );
  NAND2_X2 U_addrdec_U200 ( .A1(U_addrdec_n183), .A2(U_addrdec_n182), .ZN(
        U_addrdec_n184) );
  AOI211_X2 U_addrdec_U199 ( .C1(U_addrdec_n36), .C2(U_addrdec_n265), .A(
        U_addrdec_n185), .B(U_addrdec_n184), .ZN(U_addrdec_n190) );
  AOI22_X2 U_addrdec_U198 ( .A1(U_addrdec_n26), .A2(U_addrdec_n254), .B1(
        U_addrdec_n242), .B2(U_addrdec_n269), .ZN(U_addrdec_n189) );
  AOI22_X2 U_addrdec_U197 ( .A1(U_addrdec_n30), .A2(U_addrdec_n266), .B1(
        U_addrdec_n264), .B2(U_addrdec_n35), .ZN(U_addrdec_n188) );
  NAND3_X2 U_addrdec_U196 ( .A1(U_addrdec_n190), .A2(U_addrdec_n189), .A3(
        U_addrdec_n188), .ZN(debug_ad_row_addr[7]) );
  AOI22_X2 U_addrdec_U195 ( .A1(U_addrdec_n28), .A2(U_addrdec_n242), .B1(
        U_addrdec_n232), .B2(U_addrdec_n18), .ZN(U_addrdec_n236) );
  AOI22_X2 U_addrdec_U194 ( .A1(U_addrdec_n37), .A2(U_addrdec_n254), .B1(
        U_addrdec_n265), .B2(U_addrdec_n272), .ZN(U_addrdec_n235) );
  AOI22_X2 U_addrdec_U193 ( .A1(U_addrdec_n270), .A2(U_addrdec_n36), .B1(
        U_addrdec_n268), .B2(U_addrdec_n30), .ZN(U_addrdec_n234) );
  NAND4_X2 U_addrdec_U192 ( .A1(U_addrdec_n236), .A2(U_addrdec_n235), .A3(
        U_addrdec_n234), .A4(U_addrdec_n233), .ZN(U_addrdec_n240) );
  AOI22_X2 U_addrdec_U191 ( .A1(U_addrdec_n17), .A2(U_addrdec_n266), .B1(
        U_addrdec_n264), .B2(U_addrdec_n38), .ZN(U_addrdec_n238) );
  AOI22_X2 U_addrdec_U190 ( .A1(U_addrdec_n26), .A2(U_addrdec_n273), .B1(
        U_addrdec_n267), .B2(U_addrdec_n269), .ZN(U_addrdec_n237) );
  NAND2_X2 U_addrdec_U189 ( .A1(U_addrdec_n238), .A2(U_addrdec_n237), .ZN(
        U_addrdec_n239) );
  OAI21_X2 U_addrdec_U188 ( .B1(U_addrdec_n240), .B2(U_addrdec_n239), .A(
        U_addrdec_row_addr_mask[12]), .ZN(U_addrdec_n241) );
  INV_X4 U_addrdec_U187 ( .A(U_addrdec_n241), .ZN(debug_ad_row_addr[12]) );
  OAI22_X2 U_addrdec_U186 ( .A1(U_addrdec_n180), .A2(U_addrdec_n150), .B1(
        U_addrdec_n13), .B2(U_addrdec_n161), .ZN(U_addrdec_n145) );
  AOI22_X2 U_addrdec_U185 ( .A1(U_addrdec_n26), .A2(U_addrdec_n181), .B1(
        U_addrdec_n34), .B2(U_addrdec_n269), .ZN(U_addrdec_n143) );
  AOI22_X2 U_addrdec_U184 ( .A1(U_addrdec_n35), .A2(U_addrdec_n219), .B1(
        U_addrdec_n242), .B2(U_addrdec_n30), .ZN(U_addrdec_n142) );
  NAND2_X2 U_addrdec_U183 ( .A1(U_addrdec_n143), .A2(U_addrdec_n142), .ZN(
        U_addrdec_n144) );
  AOI211_X2 U_addrdec_U182 ( .C1(U_addrdec_n38), .C2(debug_ad_col_addr_15_), 
        .A(U_addrdec_n145), .B(U_addrdec_n144), .ZN(U_addrdec_n149) );
  AOI22_X2 U_addrdec_U181 ( .A1(debug_ad_col_addr_13__BAR_BAR), .A2(
        U_addrdec_n28), .B1(U_addrdec_n232), .B2(U_addrdec_n36), .ZN(
        U_addrdec_n148) );
  AOI22_X2 U_addrdec_U180 ( .A1(debug_ad_col_addr_12__BAR_BAR), .A2(
        U_addrdec_n18), .B1(debug_ad_col_addr_14_), .B2(U_addrdec_n37), .ZN(
        U_addrdec_n147) );
  NAND3_X2 U_addrdec_U179 ( .A1(U_addrdec_n149), .A2(U_addrdec_n148), .A3(
        U_addrdec_n147), .ZN(debug_ad_row_addr[3]) );
  OAI22_X2 U_addrdec_U178 ( .A1(U_addrdec_n180), .A2(U_addrdec_n243), .B1(
        U_addrdec_n13), .B2(U_addrdec_n23), .ZN(U_addrdec_n174) );
  AOI22_X2 U_addrdec_U177 ( .A1(U_addrdec_n38), .A2(U_addrdec_n34), .B1(
        U_addrdec_n181), .B2(U_addrdec_n272), .ZN(U_addrdec_n172) );
  AOI22_X2 U_addrdec_U176 ( .A1(U_addrdec_n17), .A2(U_addrdec_n219), .B1(
        U_addrdec_n242), .B2(U_addrdec_n26), .ZN(U_addrdec_n171) );
  NAND2_X2 U_addrdec_U175 ( .A1(U_addrdec_n172), .A2(U_addrdec_n171), .ZN(
        U_addrdec_n173) );
  AOI211_X2 U_addrdec_U174 ( .C1(U_addrdec_n18), .C2(debug_ad_col_addr_15_), 
        .A(U_addrdec_n174), .B(U_addrdec_n173), .ZN(U_addrdec_n179) );
  AOI22_X2 U_addrdec_U173 ( .A1(U_addrdec_n269), .A2(U_addrdec_n232), .B1(
        U_addrdec_n254), .B2(U_addrdec_n35), .ZN(U_addrdec_n178) );
  AOI22_X2 U_addrdec_U172 ( .A1(U_addrdec_n30), .A2(U_addrdec_n265), .B1(
        U_addrdec_n264), .B2(U_addrdec_n36), .ZN(U_addrdec_n177) );
  NAND3_X2 U_addrdec_U171 ( .A1(U_addrdec_n179), .A2(U_addrdec_n178), .A3(
        U_addrdec_n177), .ZN(debug_ad_row_addr[6]) );
  OAI22_X2 U_addrdec_U170 ( .A1(U_addrdec_n210), .A2(U_addrdec_n23), .B1(
        U_addrdec_n13), .B2(U_addrdec_n245), .ZN(U_addrdec_n194) );
  AOI22_X2 U_addrdec_U169 ( .A1(U_addrdec_n28), .A2(U_addrdec_n34), .B1(
        U_addrdec_n232), .B2(U_addrdec_n272), .ZN(U_addrdec_n192) );
  AOI22_X2 U_addrdec_U168 ( .A1(U_addrdec_n38), .A2(U_addrdec_n219), .B1(
        U_addrdec_n242), .B2(U_addrdec_n17), .ZN(U_addrdec_n191) );
  NAND2_X2 U_addrdec_U167 ( .A1(U_addrdec_n192), .A2(U_addrdec_n191), .ZN(
        U_addrdec_n193) );
  AOI211_X2 U_addrdec_U166 ( .C1(U_addrdec_n36), .C2(U_addrdec_n266), .A(
        U_addrdec_n194), .B(U_addrdec_n193), .ZN(U_addrdec_n199) );
  AOI22_X2 U_addrdec_U165 ( .A1(U_addrdec_n269), .A2(U_addrdec_n254), .B1(
        U_addrdec_n264), .B2(U_addrdec_n26), .ZN(U_addrdec_n198) );
  AOI22_X2 U_addrdec_U164 ( .A1(U_addrdec_n35), .A2(U_addrdec_n265), .B1(
        U_addrdec_n267), .B2(U_addrdec_n30), .ZN(U_addrdec_n197) );
  NAND3_X2 U_addrdec_U163 ( .A1(U_addrdec_n199), .A2(U_addrdec_n198), .A3(
        U_addrdec_n197), .ZN(debug_ad_row_addr[8]) );
  OAI22_X2 U_addrdec_U162 ( .A1(U_addrdec_n180), .A2(U_addrdec_n22), .B1(
        U_addrdec_n13), .B2(U_addrdec_n150), .ZN(U_addrdec_n154) );
  AOI22_X2 U_addrdec_U161 ( .A1(U_addrdec_n26), .A2(U_addrdec_n219), .B1(
        U_addrdec_n181), .B2(U_addrdec_n269), .ZN(U_addrdec_n152) );
  AOI22_X2 U_addrdec_U160 ( .A1(U_addrdec_n17), .A2(U_addrdec_n34), .B1(
        U_addrdec_n232), .B2(U_addrdec_n35), .ZN(U_addrdec_n151) );
  NAND2_X2 U_addrdec_U159 ( .A1(U_addrdec_n152), .A2(U_addrdec_n151), .ZN(
        U_addrdec_n153) );
  AOI211_X2 U_addrdec_U158 ( .C1(U_addrdec_n37), .C2(debug_ad_col_addr_15_), 
        .A(U_addrdec_n154), .B(U_addrdec_n153), .ZN(U_addrdec_n160) );
  AOI22_X2 U_addrdec_U157 ( .A1(U_addrdec_n30), .A2(U_addrdec_n254), .B1(
        U_addrdec_n242), .B2(U_addrdec_n36), .ZN(U_addrdec_n159) );
  AOI22_X2 U_addrdec_U156 ( .A1(debug_ad_col_addr_13__BAR_BAR), .A2(
        U_addrdec_n18), .B1(debug_ad_col_addr_14_), .B2(U_addrdec_n28), .ZN(
        U_addrdec_n158) );
  NAND3_X2 U_addrdec_U155 ( .A1(U_addrdec_n160), .A2(U_addrdec_n159), .A3(
        U_addrdec_n158), .ZN(debug_ad_row_addr[4]) );
  OAI22_X2 U_addrdec_U154 ( .A1(U_addrdec_n180), .A2(U_addrdec_n256), .B1(
        U_addrdec_n13), .B2(U_addrdec_n24), .ZN(U_addrdec_n112) );
  AOI22_X2 U_addrdec_U153 ( .A1(U_addrdec_n30), .A2(U_addrdec_n181), .B1(
        U_addrdec_n34), .B2(U_addrdec_n36), .ZN(U_addrdec_n109) );
  NAND2_X2 U_addrdec_U152 ( .A1(U_addrdec_n110), .A2(U_addrdec_n109), .ZN(
        U_addrdec_n111) );
  AOI211_X2 U_addrdec_U151 ( .C1(U_addrdec_n272), .C2(
        debug_ad_col_addr_13__BAR_BAR), .A(U_addrdec_n112), .B(U_addrdec_n111), 
        .ZN(U_addrdec_n120) );
  AOI22_X2 U_addrdec_U150 ( .A1(U_addrdec_n37), .A2(debug_ad_col_addr_11_), 
        .B1(debug_ad_col_addr_15_), .B2(U_addrdec_n269), .ZN(U_addrdec_n119)
         );
  AOI22_X2 U_addrdec_U149 ( .A1(debug_ad_col_addr_12__BAR_BAR), .A2(
        U_addrdec_n38), .B1(debug_ad_col_addr_14_), .B2(U_addrdec_n17), .ZN(
        U_addrdec_n118) );
  NAND3_X2 U_addrdec_U148 ( .A1(U_addrdec_n120), .A2(U_addrdec_n119), .A3(
        U_addrdec_n118), .ZN(debug_ad_row_addr[0]) );
  INV_X4 U_addrdec_U147 ( .A(U_addrdec_n219), .ZN(U_addrdec_n211) );
  OAI22_X2 U_addrdec_U146 ( .A1(U_addrdec_n211), .A2(U_addrdec_n243), .B1(
        U_addrdec_n210), .B2(U_addrdec_n245), .ZN(U_addrdec_n215) );
  AOI22_X2 U_addrdec_U145 ( .A1(U_addrdec_n272), .A2(U_addrdec_n254), .B1(
        U_addrdec_n232), .B2(U_addrdec_n37), .ZN(U_addrdec_n213) );
  AOI22_X2 U_addrdec_U144 ( .A1(U_addrdec_n38), .A2(U_addrdec_n242), .B1(
        U_addrdec_n264), .B2(U_addrdec_n17), .ZN(U_addrdec_n212) );
  NAND2_X2 U_addrdec_U143 ( .A1(U_addrdec_n213), .A2(U_addrdec_n212), .ZN(
        U_addrdec_n214) );
  AOI211_X2 U_addrdec_U142 ( .C1(U_addrdec_n36), .C2(U_addrdec_n273), .A(
        U_addrdec_n215), .B(U_addrdec_n214), .ZN(U_addrdec_n218) );
  AOI22_X2 U_addrdec_U141 ( .A1(U_addrdec_n269), .A2(U_addrdec_n265), .B1(
        U_addrdec_n266), .B2(U_addrdec_n26), .ZN(U_addrdec_n217) );
  AOI22_X2 U_addrdec_U140 ( .A1(U_addrdec_n267), .A2(U_addrdec_n35), .B1(
        U_addrdec_n271), .B2(U_addrdec_n30), .ZN(U_addrdec_n216) );
  NAND3_X2 U_addrdec_U139 ( .A1(U_addrdec_n218), .A2(U_addrdec_n217), .A3(
        U_addrdec_n216), .ZN(debug_ad_row_addr[10]) );
  AOI22_X2 U_addrdec_U138 ( .A1(U_addrdec_n18), .A2(U_addrdec_n254), .B1(
        U_addrdec_n264), .B2(U_addrdec_n28), .ZN(U_addrdec_n262) );
  OAI22_X2 U_addrdec_U137 ( .A1(U_addrdec_n257), .A2(U_addrdec_n256), .B1(
        U_addrdec_n255), .B2(U_addrdec_n24), .ZN(U_addrdec_n258) );
  AOI21_X2 U_addrdec_U136 ( .B1(U_addrdec_n269), .B2(U_addrdec_n271), .A(
        U_addrdec_n258), .ZN(U_addrdec_n261) );
  AOI22_X2 U_addrdec_U135 ( .A1(U_addrdec_n38), .A2(U_addrdec_n266), .B1(
        U_addrdec_n265), .B2(U_addrdec_n37), .ZN(U_addrdec_n260) );
  AOI22_X2 U_addrdec_U134 ( .A1(U_addrdec_n17), .A2(U_addrdec_n273), .B1(
        U_addrdec_n267), .B2(U_addrdec_n272), .ZN(U_addrdec_n259) );
  NAND4_X2 U_addrdec_U133 ( .A1(U_addrdec_n262), .A2(U_addrdec_n261), .A3(
        U_addrdec_n260), .A4(U_addrdec_n259), .ZN(U_addrdec_n263) );
  NOR3_X2 U_addrdec_U132 ( .A1(U_addrdec_flash_select_0_), .A2(
        U_addrdec_rom_select_0_), .A3(U_addrdec_sram_select_0_), .ZN(
        U_addrdec_n311) );
  NOR3_X2 U_addrdec_U131 ( .A1(U_addrdec_n311), .A2(ad_sdram_type_0_), .A3(
        U_addrdec_n310), .ZN(ad_static_mem_req) );
  AOI22_X2 U_addrdec_U130 ( .A1(hiu_haddr[0]), .A2(hiu_hsize[0]), .B1(
        hiu_haddr[1]), .B2(U_addrdec_n293), .ZN(U_addrdec_n295) );
  NOR2_X2 U_addrdec_U129 ( .A1(hiu_haddr[0]), .A2(hiu_hsize[0]), .ZN(
        U_addrdec_n300) );
  AOI22_X2 U_addrdec_U128 ( .A1(big_endian), .A2(U_addrdec_n295), .B1(
        U_addrdec_n296), .B2(U_addrdec_n40), .ZN(U_addrdec_n294) );
  NAND2_X2 U_addrdec_U127 ( .A1(hiu_haddr[1]), .A2(hiu_haddr[0]), .ZN(
        U_addrdec_n297) );
  AOI21_X2 U_addrdec_U126 ( .B1(U_addrdec_n294), .B2(U_addrdec_n297), .A(
        U_addrdec_n301), .ZN(ad_cr_data_mask[1]) );
  AOI22_X2 U_addrdec_U125 ( .A1(big_endian), .A2(hiu_haddr[1]), .B1(
        U_addrdec_n291), .B2(U_addrdec_n40), .ZN(U_addrdec_n299) );
  AOI221_X2 U_addrdec_U124 ( .B1(hiu_haddr[0]), .B2(big_endian), .C1(
        U_addrdec_n300), .C2(U_addrdec_n40), .A(U_addrdec_n303), .ZN(
        U_addrdec_n302) );
  NOR2_X2 U_addrdec_U123 ( .A1(U_addrdec_n302), .A2(U_addrdec_n301), .ZN(
        ad_cr_data_mask[3]) );
  AOI221_X2 U_addrdec_U122 ( .B1(U_addrdec_n300), .B2(big_endian), .C1(
        hiu_haddr[0]), .C2(U_addrdec_n40), .A(U_addrdec_n299), .ZN(
        U_addrdec_n292) );
  NOR2_X2 U_addrdec_U121 ( .A1(U_addrdec_n292), .A2(U_addrdec_n301), .ZN(
        ad_cr_data_mask[0]) );
  AOI22_X2 U_addrdec_U120 ( .A1(big_endian), .A2(U_addrdec_n296), .B1(
        U_addrdec_n295), .B2(U_addrdec_n40), .ZN(U_addrdec_n298) );
  AOI21_X2 U_addrdec_U119 ( .B1(U_addrdec_n298), .B2(U_addrdec_n297), .A(
        U_addrdec_n301), .ZN(ad_cr_data_mask[2]) );
  INV_X4 U_addrdec_U118 ( .A(U_addrdec_n96), .ZN(debug_ad_col_addr_1_) );
  INV_X4 U_addrdec_U117 ( .A(U_addrdec_n97), .ZN(debug_ad_col_addr_4_) );
  INV_X4 U_addrdec_U116 ( .A(U_addrdec_n99), .ZN(debug_ad_col_addr_6_) );
  INV_X4 U_addrdec_U115 ( .A(U_addrdec_n98), .ZN(debug_ad_col_addr_5_) );
  INV_X4 U_addrdec_U114 ( .A(U_addrdec_n100), .ZN(debug_ad_col_addr_7_) );
  NAND2_X2 U_addrdec_U113 ( .A1(U_addrdec_n282), .A2(U_addrdec_n281), .ZN(
        U_addrdec_n283) );
  NAND2_X2 U_addrdec_U112 ( .A1(U_addrdec_n281), .A2(U_addrdec_n280), .ZN(
        U_addrdec_n286) );
  OAI221_X2 U_addrdec_U111 ( .B1(cr_row_addr_width[2]), .B2(
        cr_row_addr_width[1]), .C1(U_addrdec_n290), .C2(U_cr_n21), .A(
        cr_row_addr_width[3]), .ZN(U_addrdec_N133) );
  NOR3_X2 U_addrdec_U110 ( .A1(cr_block_size1[7]), .A2(cr_block_size1[5]), 
        .A3(cr_block_size1[6]), .ZN(U_addrdec_n347) );
  NAND2_X2 U_addrdec_U109 ( .A1(cr_block_size1[5]), .A2(U_cr_n167), .ZN(
        U_addrdec_n309) );
  NOR2_X2 U_addrdec_U108 ( .A1(cr_block_size1[6]), .A2(U_addrdec_n309), .ZN(
        U_addrdec_n348) );
  NOR3_X2 U_addrdec_U107 ( .A1(cr_block_size1[7]), .A2(cr_block_size1[5]), 
        .A3(U_cr_n119), .ZN(U_addrdec_n346) );
  NOR2_X2 U_addrdec_U106 ( .A1(U_addrdec_n309), .A2(U_cr_n119), .ZN(
        U_addrdec_n345) );
  NOR2_X2 U_addrdec_U105 ( .A1(U_addrdec_n114), .A2(U_addrdec_n116), .ZN(
        U_addrdec_n269) );
  NAND2_X4 U_addrdec_U104 ( .A1(U_addrdec_n54), .A2(U_addrdec_n53), .ZN(
        debug_ad_col_addr_11_) );
  NOR2_X1 U_addrdec_U103 ( .A1(U_addrdec_n39), .A2(U_addrdec_n95), .ZN(
        debug_ad_col_addr_0_) );
  NOR2_X1 U_addrdec_U102 ( .A1(n27), .A2(U_addrdec_n303), .ZN(U_addrdec_n304)
         );
  NAND2_X2 U_addrdec_U101 ( .A1(hiu_addr[11]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n53) );
  NAND2_X1 U_addrdec_U100 ( .A1(n27), .A2(U_addrdec_n306), .ZN(ad_data_mask[3]) );
  NAND2_X1 U_addrdec_U99 ( .A1(n27), .A2(U_addrdec_n305), .ZN(ad_data_mask[2])
         );
  AOI22_X2 U_addrdec_U98 ( .A1(U_addrdec_n28), .A2(debug_ad_col_addr_10_), 
        .B1(debug_ad_col_addr_9_), .B2(U_addrdec_n18), .ZN(U_addrdec_n110) );
  INV_X1 U_addrdec_U97 ( .A(debug_ad_col_addr_13_), .ZN(
        debug_ad_col_addr_13__BAR_BAR) );
  AOI211_X4 U_addrdec_U90 ( .C1(U_addrdec_n18), .C2(debug_ad_col_addr_14_), 
        .A(U_addrdec_n165), .B(U_addrdec_n164), .ZN(U_addrdec_n170) );
  NAND2_X1 U_addrdec_U89 ( .A1(n[26]), .A2(cr_bank_addr_width[0]), .ZN(
        U_addrdec_n42) );
  OR2_X2 U_addrdec_U87 ( .A1(cr_bank_addr_width[1]), .A2(cr_bank_addr_width[0]), .ZN(U_addrdec_N119) );
  NAND2_X1 U_addrdec_U84 ( .A1(cr_row_addr_width[2]), .A2(cr_row_addr_width[3]), .ZN(U_addrdec_n287) );
  NAND2_X1 U_addrdec_U81 ( .A1(cr_row_addr_width[2]), .A2(cr_row_addr_width[1]), .ZN(U_addrdec_n290) );
  NAND3_X1 U_addrdec_U79 ( .A1(cr_row_addr_width[1]), .A2(cr_row_addr_width[3]), .A3(U_cr_n55), .ZN(U_addrdec_N130) );
  NAND2_X1 U_addrdec_U77 ( .A1(U_addrdec_n42), .A2(U_cr_n22), .ZN(
        U_addrdec_n280) );
  INV_X2 U_addrdec_U76 ( .A(U_addrdec_n106), .ZN(U_addrdec_n101) );
  OAI21_X1 U_addrdec_U75 ( .B1(cr_row_addr_width[1]), .B2(U_addrdec_n287), .A(
        U_addrdec_N130), .ZN(U_addrdec_n58) );
  OR2_X2 U_addrdec_U74 ( .A1(U_addrdec_N130), .A2(cr_row_addr_width[0]), .ZN(
        U_addrdec_N129) );
  NAND2_X1 U_addrdec_U73 ( .A1(U_addrdec_n41), .A2(n[25]), .ZN(U_addrdec_n281)
         );
  INV_X1 U_addrdec_U72 ( .A(U_addrdec_n81), .ZN(U_addrdec_n56) );
  NAND2_X1 U_addrdec_U71 ( .A1(hiu_addr[28]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n205) );
  NAND2_X1 U_addrdec_U70 ( .A1(hiu_addr[29]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n206) );
  NAND2_X1 U_addrdec_U69 ( .A1(hiu_addr[28]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n196) );
  OAI21_X1 U_addrdec_U68 ( .B1(U_cr_n21), .B2(U_cr_n55), .A(U_addrdec_n58), 
        .ZN(U_addrdec_N131) );
  INV_X2 U_addrdec_U67 ( .A(hiu_addr[1]), .ZN(U_addrdec_n95) );
  NAND2_X1 U_addrdec_U66 ( .A1(U_addrdec_n283), .A2(n[24]), .ZN(U_addrdec_n285) );
  INV_X1 U_addrdec_U65 ( .A(hiu_haddr[0]), .ZN(U_addrdec_n293) );
  NAND2_X1 U_addrdec_U64 ( .A1(hiu_addr[18]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n104) );
  NAND2_X1 U_addrdec_U63 ( .A1(hiu_addr[17]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n103) );
  NAND2_X1 U_addrdec_U62 ( .A1(hiu_addr[19]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n108) );
  INV_X2 U_addrdec_U59 ( .A(U_addrdec_n255), .ZN(U_addrdec_n268) );
  INV_X2 U_addrdec_U58 ( .A(U_addrdec_n272), .ZN(U_addrdec_n150) );
  INV_X2 U_addrdec_U57 ( .A(U_addrdec_n269), .ZN(U_addrdec_n130) );
  INV_X2 U_addrdec_U56 ( .A(U_addrdec_n254), .ZN(U_addrdec_n244) );
  INV_X2 U_addrdec_U55 ( .A(U_addrdec_n242), .ZN(U_addrdec_n246) );
  NAND2_X1 U_addrdec_U54 ( .A1(U_addrdec_n271), .A2(U_addrdec_n35), .ZN(
        U_addrdec_n233) );
  NAND2_X1 U_addrdec_U53 ( .A1(U_addrdec_n271), .A2(U_addrdec_n36), .ZN(
        U_addrdec_n223) );
  NOR2_X2 U_addrdec_U49 ( .A1(U_addrdec_n32), .A2(U_addrdec_n27), .ZN(
        debug_ad_col_addr_12_) );
  INV_X2 U_addrdec_U48 ( .A(U_addrdec_n270), .ZN(U_addrdec_n257) );
  OR2_X2 U_addrdec_U47 ( .A1(hiu_haddr[1]), .A2(U_addrdec_n300), .ZN(
        U_addrdec_n296) );
  OAI21_X1 U_addrdec_U46 ( .B1(n[24]), .B2(U_addrdec_n283), .A(U_addrdec_n285), 
        .ZN(U_addrdec_n284) );
  XOR2_X1 U_addrdec_U45 ( .A(U_addrdec_n285), .B(U_cr_n65), .Z(U_addrdec_N110)
         );
  NOR2_X1 U_addrdec_U44 ( .A1(U_addrdec_n285), .A2(U_cr_n65), .ZN(
        U_addrdec_N111) );
  INV_X2 U_addrdec_U43 ( .A(debug_ad_col_addr_10_), .ZN(U_addrdec_n62) );
  INV_X2 U_addrdec_U42 ( .A(debug_ad_col_addr_9_), .ZN(U_addrdec_n61) );
  INV_X2 U_addrdec_U41 ( .A(U_addrdec_n34), .ZN(U_addrdec_n200) );
  NAND2_X1 U_addrdec_U40 ( .A1(U_addrdec_n34), .A2(U_addrdec_n272), .ZN(
        U_addrdec_n162) );
  INV_X2 U_addrdec_U39 ( .A(U_addrdec_n299), .ZN(U_addrdec_n303) );
  INV_X2 U_addrdec_U38 ( .A(U_addrdec_n284), .ZN(U_addrdec_N109) );
  INV_X1 U_addrdec_U37 ( .A(U_addrdec_n88), .ZN(U_addrdec_n59) );
  NOR2_X2 U_addrdec_U36 ( .A1(ad_sdram_chip_select_0_), .A2(U_addrdec_n310), 
        .ZN(sdram_req_i) );
  INV_X1 U_addrdec_U35 ( .A(ad_cr_data_mask[2]), .ZN(U_addrdec_n305) );
  INV_X1 U_addrdec_U34 ( .A(ad_cr_data_mask[3]), .ZN(U_addrdec_n306) );
  INV_X2 U_addrdec_U33 ( .A(U_addrdec_n86), .ZN(U_addrdec_n91) );
  INV_X1 U_addrdec_U32 ( .A(U_addrdec_n42), .ZN(U_addrdec_n41) );
  NAND2_X2 U_addrdec_U31 ( .A1(U_addrdec_n280), .A2(cr_bank_addr_width[1]), 
        .ZN(U_addrdec_n282) );
  INV_X2 U_addrdec_U30 ( .A(U_addrdec_n26), .ZN(U_addrdec_n256) );
  NAND2_X1 U_addrdec_U29 ( .A1(hiu_addr[31]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n221) );
  NAND2_X1 U_addrdec_U28 ( .A1(hiu_addr[30]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n222) );
  NAND2_X1 U_addrdec_U27 ( .A1(hiu_addr[26]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n175) );
  NAND2_X1 U_addrdec_U26 ( .A1(hiu_addr[27]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n195) );
  NAND2_X1 U_addrdec_U25 ( .A1(hiu_addr[27]), .A2(U_addrdec_n220), .ZN(
        U_addrdec_n187) );
  NAND2_X1 U_addrdec_U24 ( .A1(hiu_addr[26]), .A2(U_addrdec_n39), .ZN(
        U_addrdec_n186) );
  INV_X2 U_addrdec_U23 ( .A(hiu_haddr[1]), .ZN(U_addrdec_n291) );
  XNOR2_X1 U_addrdec_U21 ( .A(U_cr_n63), .B(cr_bank_addr_width[0]), .ZN(
        U_addrdec_N107) );
  INV_X1 U_addrdec_U20 ( .A(U_addrdec_n11), .ZN(U_addrdec_n271) );
  AOI22_X1 U_addrdec_U19 ( .A1(U_addrdec_n220), .A2(hiu_addr[30]), .B1(
        U_addrdec_n39), .B2(hiu_addr[29]), .ZN(U_addrdec_n11) );
  INV_X1 U_addrdec_U18 ( .A(U_addrdec_n10), .ZN(U_addrdec_n34) );
  AOI22_X1 U_addrdec_U17 ( .A1(U_addrdec_n39), .A2(hiu_addr[18]), .B1(
        U_addrdec_n220), .B2(hiu_addr[19]), .ZN(U_addrdec_n10) );
  INV_X1 U_addrdec_U16 ( .A(U_addrdec_n9), .ZN(debug_ad_col_addr_3_) );
  AOI22_X1 U_addrdec_U15 ( .A1(hiu_addr[4]), .A2(U_addrdec_n220), .B1(
        hiu_addr[3]), .B2(U_addrdec_n39), .ZN(U_addrdec_n9) );
  AOI22_X2 U_addrdec_U14 ( .A1(U_addrdec_bcawp_3_), .A2(U_addrdec_n15), .B1(
        U_addrdec_n5), .B2(U_addrdec_n7), .ZN(U_addrdec_n30) );
  AOI22_X2 U_addrdec_U13 ( .A1(U_addrdec_n15), .A2(U_addrdec_n20), .B1(
        U_addrdec_bcawp_0_), .B2(U_addrdec_n21), .ZN(U_addrdec_n7) );
  AOI221_X2 U_addrdec_U12 ( .B1(U_addrdec_bcawp_3_), .B2(U_addrdec_bcawp_4_), 
        .C1(U_addrdec_bcawp_2_), .C2(U_addrdec_bcawp_4_), .A(U_addrdec_n4), 
        .ZN(U_addrdec_n5) );
  INV_X4 U_addrdec_U11 ( .A(U_addrdec_n115), .ZN(U_addrdec_n4) );
  NAND4_X1 U_addrdec_U10 ( .A1(U_addrdec_n14), .A2(U_addrdec_bcawp_4_), .A3(
        U_addrdec_n20), .A4(U_addrdec_n3), .ZN(U_addrdec_n25) );
  INV_X1 U_addrdec_U9 ( .A(U_addrdec_n113), .ZN(U_addrdec_n3) );
  OR2_X1 U_addrdec_U8 ( .A1(hiu_hsize[2]), .A2(hiu_hsize[1]), .ZN(
        U_addrdec_n301) );
  INV_X1 U_addrdec_U7 ( .A(U_addrdec_n2), .ZN(debug_ad_col_addr_2_) );
  AOI22_X1 U_addrdec_U6 ( .A1(hiu_addr[2]), .A2(U_addrdec_n39), .B1(
        hiu_addr[3]), .B2(U_addrdec_n220), .ZN(U_addrdec_n2) );
  INV_X1 U_addrdec_U5 ( .A(U_addrdec_n1), .ZN(U_addrdec_n102) );
  AOI22_X2 U_addrdec_U4 ( .A1(U_addrdec_n220), .A2(hiu_addr[17]), .B1(
        U_addrdec_n39), .B2(hiu_addr[16]), .ZN(U_addrdec_n1) );
  NAND2_X2 U_addrdec_U3 ( .A1(U_addrdec_n122), .A2(U_addrdec_n121), .ZN(
        U_addrdec_n219) );
  DFFR_X2 U_addrdec_bcawp_reg_3_ ( .D(U_addrdec_N110), .CK(hclk), .RN(hresetn), 
        .Q(U_addrdec_bcawp_3_), .QN(U_addrdec_n14) );
  DFFR_X2 U_addrdec_bcawp_reg_2_ ( .D(U_addrdec_N109), .CK(hclk), .RN(hresetn), 
        .Q(U_addrdec_bcawp_2_), .QN(U_addrdec_n16) );
  DFFR_X2 U_addrdec_bcawp_reg_1_ ( .D(U_addrdec_N108), .CK(hclk), .RN(hresetn), 
        .Q(U_addrdec_bcawp_1_), .QN(U_addrdec_n21) );
  DFFR_X2 U_addrdec_bcawp_reg_4_ ( .D(U_addrdec_N111), .CK(hclk), .RN(hresetn), 
        .Q(U_addrdec_bcawp_4_), .QN(U_addrdec_n15) );
  DFFR_X2 U_addrdec_bcawp_reg_0_ ( .D(U_addrdec_N107), .CK(hclk), .RN(hresetn), 
        .Q(U_addrdec_bcawp_0_), .QN(U_addrdec_n20) );
  DFFR_X2 U_addrdec_sdram_select_reg_0_ ( .D(U_addrdec_n347), .CK(hclk), .RN(
        hresetn), .Q(ad_sdram_type_0_), .QN(ad_sdram_chip_select_0_) );
  DFFR_X2 U_addrdec_s_data_width_prog_buf_reg_0_ ( .D(n27), .CK(hclk), .RN(
        hresetn), .Q(U_addrdec_n220), .QN(U_addrdec_n39) );
  DFFR_X2 U_addrdec_sram_select_reg_0_ ( .D(U_addrdec_n348), .CK(hclk), .RN(
        hresetn), .Q(U_addrdec_sram_select_0_) );
  DFFR_X2 U_addrdec_rom_select_reg_0_ ( .D(U_addrdec_n345), .CK(hclk), .RN(
        hresetn), .Q(U_addrdec_rom_select_0_) );
  DFFR_X2 U_addrdec_flash_select_reg_0_ ( .D(U_addrdec_n346), .CK(hclk), .RN(
        hresetn), .Q(U_addrdec_flash_select_0_) );
  DFFS_X2 U_addrdec_row_addr_mask_hi_reg_0_ ( .D(U_addrdec_N129), .CK(hclk), 
        .SN(hresetn), .Q(U_addrdec_row_addr_mask[11]) );
  DFFS_X2 U_addrdec_row_addr_mask_hi_reg_1_ ( .D(U_addrdec_N130), .CK(hclk), 
        .SN(hresetn), .Q(U_addrdec_row_addr_mask[12]) );
  DFFS_X2 U_addrdec_row_addr_mask_hi_reg_2_ ( .D(U_addrdec_N131), .CK(hclk), 
        .SN(hresetn), .Q(U_addrdec_row_addr_mask[13]) );
  DFFR_X1 U_addrdec_row_addr_mask_hi_reg_3_ ( .D(U_addrdec_n58), .CK(hclk), 
        .RN(hresetn), .QN(U_addrdec_row_addr_mask[14]) );
  DFFS_X2 U_addrdec_row_addr_mask_hi_reg_4_ ( .D(U_addrdec_N133), .CK(hclk), 
        .SN(hresetn), .Q(U_addrdec_row_addr_mask[15]) );
  DFFS_X2 U_addrdec_bank_addr_mask_reg_1_ ( .D(U_addrdec_N119), .CK(hclk), 
        .SN(hresetn), .Q(U_addrdec_bank_addr_mask_1_) );
  OAI221_X2 U_refctl_U142 ( .B1(U_refctl_current_state_1_), .B2(
        U_refctl_current_state_0_), .C1(U_refctl_current_state_1_), .C2(
        U_refctl_n97), .A(ctl_auto_ref_en), .ZN(U_refctl_n112) );
  NOR2_X2 U_refctl_U141 ( .A1(U_refctl_n112), .A2(U_refctl_count_0_), .ZN(
        U_refctl_count_next_0_) );
  NOR2_X2 U_refctl_U140 ( .A1(U_refctl_N27), .A2(U_refctl_n91), .ZN(
        U_refctl_n119) );
  OAI22_X2 U_refctl_U139 ( .A1(U_refctl_N29), .A2(U_refctl_n81), .B1(
        U_refctl_N28), .B2(U_refctl_n86), .ZN(U_refctl_n120) );
  AOI22_X2 U_refctl_U138 ( .A1(U_refctl_N22), .A2(U_refctl_n87), .B1(
        U_refctl_N23), .B2(U_refctl_n78), .ZN(U_refctl_n115) );
  AOI211_X2 U_refctl_U137 ( .C1(U_refctl_n121), .C2(U_refctl_count_12_), .A(
        U_refctl_n120), .B(U_refctl_n119), .ZN(U_refctl_n122) );
  INV_X4 U_refctl_U136 ( .A(U_refctl_n124), .ZN(U_refctl_n127) );
  AOI221_X2 U_refctl_U135 ( .B1(U_refctl_current_state_1_), .B2(U_refctl_n127), 
        .C1(U_refctl_n92), .C2(U_refctl_n126), .A(n94), .ZN(
        U_refctl_ref_req_next) );
  NAND4_X2 U_refctl_U134 ( .A1(U_refctl_count_3_), .A2(U_refctl_count_2_), 
        .A3(U_refctl_count_1_), .A4(U_refctl_count_0_), .ZN(U_refctl_n106) );
  NOR2_X2 U_refctl_U133 ( .A1(U_refctl_n84), .A2(U_refctl_n106), .ZN(
        U_refctl_n105) );
  INV_X4 U_refctl_U132 ( .A(U_refctl_n105), .ZN(U_refctl_n107) );
  NOR2_X2 U_refctl_U131 ( .A1(U_refctl_n85), .A2(U_refctl_n107), .ZN(
        U_refctl_n108) );
  NAND2_X2 U_refctl_U130 ( .A1(U_refctl_count_6_), .A2(U_refctl_n108), .ZN(
        U_refctl_n109) );
  NOR2_X2 U_refctl_U129 ( .A1(U_refctl_n89), .A2(U_refctl_n109), .ZN(
        U_refctl_n110) );
  NAND2_X2 U_refctl_U128 ( .A1(U_refctl_count_8_), .A2(U_refctl_n110), .ZN(
        U_refctl_n113) );
  NOR2_X2 U_refctl_U127 ( .A1(U_refctl_n78), .A2(U_refctl_n113), .ZN(
        U_refctl_n111) );
  NAND2_X2 U_refctl_U126 ( .A1(U_refctl_count_10_), .A2(U_refctl_n111), .ZN(
        U_refctl_n98) );
  NOR2_X2 U_refctl_U125 ( .A1(U_refctl_n80), .A2(U_refctl_n98), .ZN(
        U_refctl_n99) );
  NAND2_X2 U_refctl_U124 ( .A1(U_refctl_count_12_), .A2(U_refctl_n99), .ZN(
        U_refctl_n100) );
  NOR2_X2 U_refctl_U123 ( .A1(U_refctl_n91), .A2(U_refctl_n100), .ZN(
        U_refctl_n101) );
  AOI211_X2 U_refctl_U122 ( .C1(U_refctl_n91), .C2(U_refctl_n100), .A(
        U_refctl_n112), .B(U_refctl_n101), .ZN(U_refctl_count_next_13_) );
  AOI211_X2 U_refctl_U121 ( .C1(U_refctl_n78), .C2(U_refctl_n113), .A(
        U_refctl_n112), .B(U_refctl_n111), .ZN(U_refctl_count_next_9_) );
  AOI211_X2 U_refctl_U120 ( .C1(U_refctl_n84), .C2(U_refctl_n106), .A(
        U_refctl_n112), .B(U_refctl_n105), .ZN(U_refctl_count_next_4_) );
  AOI211_X2 U_refctl_U119 ( .C1(U_refctl_n80), .C2(U_refctl_n98), .A(
        U_refctl_n112), .B(U_refctl_n99), .ZN(U_refctl_count_next_11_) );
  AOI211_X2 U_refctl_U118 ( .C1(U_refctl_n89), .C2(U_refctl_n109), .A(
        U_refctl_n112), .B(U_refctl_n110), .ZN(U_refctl_count_next_7_) );
  AOI211_X2 U_refctl_U117 ( .C1(U_refctl_n85), .C2(U_refctl_n107), .A(
        U_refctl_n112), .B(U_refctl_n108), .ZN(U_refctl_count_next_5_) );
  INV_X4 U_refctl_U116 ( .A(U_refctl_n101), .ZN(U_refctl_n102) );
  NOR2_X2 U_refctl_U115 ( .A1(U_refctl_n86), .A2(U_refctl_n102), .ZN(
        U_refctl_n104) );
  AOI211_X2 U_refctl_U114 ( .C1(U_refctl_n86), .C2(U_refctl_n102), .A(
        U_refctl_n112), .B(U_refctl_n104), .ZN(U_refctl_count_next_14_) );
  AOI21_X2 U_refctl_U113 ( .B1(U_refctl_current_state_1_), .B2(U_refctl_n124), 
        .A(U_refctl_n123), .ZN(U_refctl_next_state_0_) );
  AOI221_X2 U_refctl_U112 ( .B1(U_refctl_count_1_), .B2(U_refctl_count_0_), 
        .C1(U_refctl_n73), .C2(U_refctl_n83), .A(U_refctl_n112), .ZN(
        U_refctl_count_next_1_) );
  AOI221_X2 U_refctl_U111 ( .B1(U_refctl_count_15_), .B2(U_refctl_n104), .C1(
        U_refctl_n81), .C2(U_refctl_n103), .A(U_refctl_n112), .ZN(
        U_refctl_count_next_15_) );
  NOR4_X2 U_refctl_U110 ( .A1(U_refctl_N30), .A2(U_refctl_n66), .A3(
        U_refctl_n65), .A4(U_refctl_n64), .ZN(U_refctl_N31) );
  NAND4_X2 U_refctl_U109 ( .A1(U_refctl_n63), .A2(U_refctl_n62), .A3(
        U_refctl_n61), .A4(U_refctl_n60), .ZN(U_refctl_n64) );
  NOR4_X2 U_refctl_U108 ( .A1(U_refctl_n59), .A2(U_refctl_n58), .A3(
        U_refctl_n57), .A4(U_refctl_n56), .ZN(U_refctl_n63) );
  NAND4_X2 U_refctl_U107 ( .A1(U_refctl_n55), .A2(U_refctl_n54), .A3(
        U_refctl_n53), .A4(U_refctl_n52), .ZN(U_refctl_n56) );
  NOR4_X2 U_refctl_U106 ( .A1(U_refctl_n51), .A2(U_refctl_n50), .A3(
        U_refctl_n49), .A4(U_refctl_n48), .ZN(U_refctl_n55) );
  OAI221_X2 U_refctl_U105 ( .B1(U_refctl_count_1_), .B2(U_refctl_n47), .C1(
        cr_t_ref[0]), .C2(U_refctl_count_0_), .A(U_refctl_n46), .ZN(
        U_refctl_n48) );
  AOI22_X2 U_refctl_U104 ( .A1(U_refctl_count_1_), .A2(U_refctl_n47), .B1(
        cr_t_ref[0]), .B2(U_refctl_count_0_), .ZN(U_refctl_n46) );
  NOR3_X2 U_refctl_U103 ( .A1(cr_t_ref[2]), .A2(cr_t_ref[1]), .A3(cr_t_ref[0]), 
        .ZN(U_refctl_n33) );
  NOR2_X2 U_refctl_U102 ( .A1(cr_t_ref[1]), .A2(cr_t_ref[0]), .ZN(U_refctl_n32) );
  NOR2_X2 U_refctl_U101 ( .A1(cr_t_ref[15]), .A2(U_refctl_n45), .ZN(
        U_refctl_N30) );
  NAND2_X2 U_refctl_U100 ( .A1(U_refctl_n44), .A2(U_cr_n123), .ZN(U_refctl_n45) );
  NOR2_X2 U_refctl_U98 ( .A1(cr_t_ref[13]), .A2(U_refctl_n43), .ZN(
        U_refctl_n44) );
  NAND2_X2 U_refctl_U97 ( .A1(U_refctl_n42), .A2(U_cr_n122), .ZN(U_refctl_n43)
         );
  NOR2_X2 U_refctl_U95 ( .A1(cr_t_ref[11]), .A2(U_refctl_n41), .ZN(
        U_refctl_n42) );
  NAND2_X2 U_refctl_U94 ( .A1(U_refctl_n40), .A2(U_cr_n129), .ZN(U_refctl_n41)
         );
  NOR2_X2 U_refctl_U92 ( .A1(cr_t_ref[9]), .A2(U_refctl_n39), .ZN(U_refctl_n40) );
  NAND2_X2 U_refctl_U91 ( .A1(U_refctl_n38), .A2(U_cr_n118), .ZN(U_refctl_n39)
         );
  NOR2_X2 U_refctl_U89 ( .A1(cr_t_ref[7]), .A2(U_refctl_n37), .ZN(U_refctl_n38) );
  NAND2_X2 U_refctl_U88 ( .A1(U_refctl_n36), .A2(U_cr_n121), .ZN(U_refctl_n37)
         );
  NOR2_X2 U_refctl_U86 ( .A1(cr_t_ref[5]), .A2(U_refctl_n35), .ZN(U_refctl_n36) );
  NAND2_X2 U_refctl_U85 ( .A1(U_refctl_n34), .A2(U_cr_n130), .ZN(U_refctl_n35)
         );
  NOR4_X2 U_refctl_U83 ( .A1(cr_t_ref[3]), .A2(cr_t_ref[2]), .A3(cr_t_ref[1]), 
        .A4(cr_t_ref[0]), .ZN(U_refctl_n34) );
  XNOR2_X2 U_refctl_U82 ( .A(U_refctl_count_12_), .B(U_refctl_N26), .ZN(
        U_refctl_n61) );
  XNOR2_X2 U_refctl_U81 ( .A(U_refctl_n42), .B(U_cr_n122), .ZN(U_refctl_N26)
         );
  XNOR2_X2 U_refctl_U80 ( .A(U_refctl_count_11_), .B(U_refctl_N25), .ZN(
        U_refctl_n62) );
  XNOR2_X2 U_refctl_U79 ( .A(cr_t_ref[11]), .B(U_refctl_n41), .ZN(U_refctl_N25) );
  XNOR2_X2 U_refctl_U78 ( .A(U_refctl_count_7_), .B(U_refctl_N21), .ZN(
        U_refctl_n52) );
  XNOR2_X2 U_refctl_U77 ( .A(cr_t_ref[7]), .B(U_refctl_n37), .ZN(U_refctl_N21)
         );
  XNOR2_X2 U_refctl_U76 ( .A(U_refctl_count_5_), .B(U_refctl_N19), .ZN(
        U_refctl_n53) );
  XNOR2_X2 U_refctl_U75 ( .A(cr_t_ref[5]), .B(U_refctl_n35), .ZN(U_refctl_N19)
         );
  XNOR2_X2 U_refctl_U74 ( .A(U_refctl_n36), .B(U_cr_n121), .ZN(U_refctl_N20)
         );
  XOR2_X2 U_refctl_U73 ( .A(cr_t_ref[1]), .B(cr_t_ref[0]), .Z(U_refctl_n47) );
  XOR2_X2 U_refctl_U72 ( .A(cr_t_ref[3]), .B(U_refctl_n33), .Z(U_refctl_N17)
         );
  XOR2_X2 U_refctl_U71 ( .A(cr_t_ref[2]), .B(U_refctl_n32), .Z(U_refctl_N16)
         );
  XOR2_X2 U_refctl_U70 ( .A(U_refctl_count_4_), .B(U_refctl_N18), .Z(
        U_refctl_n51) );
  XNOR2_X2 U_refctl_U69 ( .A(U_refctl_n34), .B(U_cr_n130), .ZN(U_refctl_N18)
         );
  XOR2_X2 U_refctl_U68 ( .A(U_refctl_count_9_), .B(U_refctl_N23), .Z(
        U_refctl_n57) );
  XNOR2_X2 U_refctl_U67 ( .A(cr_t_ref[9]), .B(U_refctl_n39), .ZN(U_refctl_N23)
         );
  XOR2_X2 U_refctl_U66 ( .A(U_refctl_count_10_), .B(U_refctl_N24), .Z(
        U_refctl_n58) );
  XNOR2_X2 U_refctl_U65 ( .A(U_refctl_n40), .B(U_cr_n129), .ZN(U_refctl_N24)
         );
  XOR2_X2 U_refctl_U64 ( .A(U_refctl_count_8_), .B(U_refctl_N22), .Z(
        U_refctl_n59) );
  XNOR2_X2 U_refctl_U63 ( .A(U_refctl_n38), .B(U_cr_n118), .ZN(U_refctl_N22)
         );
  XOR2_X2 U_refctl_U62 ( .A(U_refctl_count_14_), .B(U_refctl_N28), .Z(
        U_refctl_n65) );
  XNOR2_X2 U_refctl_U61 ( .A(U_refctl_n44), .B(U_cr_n123), .ZN(U_refctl_N28)
         );
  XOR2_X2 U_refctl_U60 ( .A(U_refctl_count_15_), .B(U_refctl_N29), .Z(
        U_refctl_n66) );
  XNOR2_X2 U_refctl_U59 ( .A(cr_t_ref[15]), .B(U_refctl_n45), .ZN(U_refctl_N29) );
  XNOR2_X2 U_refctl_U58 ( .A(U_refctl_count_13_), .B(U_refctl_N27), .ZN(
        U_refctl_n60) );
  XNOR2_X2 U_refctl_U57 ( .A(cr_t_ref[13]), .B(U_refctl_n43), .ZN(U_refctl_N27) );
  XOR2_X1 U_refctl_U55 ( .A(U_refctl_count_2_), .B(U_refctl_N16), .Z(
        U_refctl_n50) );
  XOR2_X1 U_refctl_U54 ( .A(U_refctl_count_3_), .B(U_refctl_N17), .Z(
        U_refctl_n49) );
  XNOR2_X1 U_refctl_U53 ( .A(U_refctl_count_6_), .B(U_refctl_N20), .ZN(
        U_refctl_n54) );
  INV_X2 U_refctl_U52 ( .A(U_refctl_N21), .ZN(U_refctl_n118) );
  OAI21_X1 U_refctl_U51 ( .B1(U_refctl_n108), .B2(U_refctl_count_6_), .A(
        U_refctl_n109), .ZN(U_refctl_n95) );
  OAI21_X1 U_refctl_U50 ( .B1(U_refctl_n110), .B2(U_refctl_count_8_), .A(
        U_refctl_n113), .ZN(U_refctl_n96) );
  OAI211_X1 U_refctl_U49 ( .C1(U_refctl_N25), .C2(U_refctl_n80), .A(
        U_refctl_N24), .B(U_refctl_n90), .ZN(U_refctl_n114) );
  OAI21_X1 U_refctl_U48 ( .B1(U_refctl_n111), .B2(U_refctl_count_10_), .A(
        U_refctl_n98), .ZN(U_refctl_n93) );
  INV_X1 U_refctl_U47 ( .A(U_refctl_N26), .ZN(U_refctl_n121) );
  OAI21_X1 U_refctl_U46 ( .B1(U_refctl_n99), .B2(U_refctl_count_12_), .A(
        U_refctl_n100), .ZN(U_refctl_n94) );
  INV_X2 U_refctl_U45 ( .A(U_refctl_n104), .ZN(U_refctl_n103) );
  NAND2_X1 U_refctl_U44 ( .A1(U_refctl_current_state_0_), .A2(U_refctl_N31), 
        .ZN(U_refctl_n126) );
  INV_X2 U_refctl_U43 ( .A(U_refctl_N31), .ZN(U_refctl_n97) );
  OAI21_X1 U_refctl_U42 ( .B1(U_refctl_n126), .B2(U_refctl_current_state_1_), 
        .A(ctl_auto_ref_en), .ZN(U_refctl_n123) );
  NOR2_X1 U_refctl_U41 ( .A1(U_refctl_n112), .A2(U_refctl_n96), .ZN(
        U_refctl_n76) );
  NOR2_X1 U_refctl_U40 ( .A1(U_refctl_n112), .A2(U_refctl_n95), .ZN(
        U_refctl_n75) );
  NOR2_X1 U_refctl_U39 ( .A1(U_refctl_n112), .A2(U_refctl_n93), .ZN(
        U_refctl_n79) );
  NOR2_X1 U_refctl_U38 ( .A1(U_refctl_n112), .A2(U_refctl_n94), .ZN(
        U_refctl_n82) );
  AOI22_X1 U_refctl_U37 ( .A1(U_refctl_n28), .A2(U_refctl_count_3_), .B1(
        U_refctl_n74), .B2(U_refctl_n30), .ZN(U_refctl_count_next_3_) );
  NAND4_X1 U_refctl_U36 ( .A1(U_refctl_count_0_), .A2(U_refctl_count_2_), .A3(
        U_refctl_count_1_), .A4(U_refctl_n29), .ZN(U_refctl_n30) );
  INV_X1 U_refctl_U35 ( .A(U_refctl_n112), .ZN(U_refctl_n29) );
  NOR2_X1 U_refctl_U34 ( .A1(U_refctl_count_next_0_), .A2(U_refctl_n27), .ZN(
        U_refctl_n28) );
  AOI21_X1 U_refctl_U33 ( .B1(U_refctl_count_1_), .B2(U_refctl_count_2_), .A(
        U_refctl_n112), .ZN(U_refctl_n27) );
  OAI222_X1 U_refctl_U32 ( .A1(U_refctl_n78), .A2(U_refctl_N23), .B1(
        U_refctl_N24), .B2(U_refctl_n90), .C1(U_refctl_N25), .C2(U_refctl_n80), 
        .ZN(U_refctl_n116) );
  AOI221_X1 U_refctl_U30 ( .B1(U_refctl_n23), .B2(U_refctl_n25), .C1(
        U_refctl_n77), .C2(U_refctl_n25), .A(U_refctl_n112), .ZN(
        U_refctl_count_next_2_) );
  NAND3_X1 U_refctl_U29 ( .A1(U_refctl_count_0_), .A2(U_refctl_count_1_), .A3(
        U_refctl_n77), .ZN(U_refctl_n25) );
  NOR2_X1 U_refctl_U27 ( .A1(U_refctl_n83), .A2(U_refctl_n73), .ZN(
        U_refctl_n23) );
  OAI221_X1 U_refctl_U26 ( .B1(U_refctl_N20), .B2(U_refctl_n21), .C1(
        U_refctl_n88), .C2(U_refctl_n22), .A(U_refctl_n11), .ZN(U_refctl_n117)
         );
  AND2_X1 U_refctl_U25 ( .A1(U_refctl_N20), .A2(U_refctl_n21), .ZN(
        U_refctl_n22) );
  AOI222_X1 U_refctl_U24 ( .A1(U_refctl_count_5_), .A2(U_refctl_n19), .B1(
        U_refctl_count_5_), .B2(U_refctl_n20), .C1(U_refctl_n19), .C2(
        U_refctl_n20), .ZN(U_refctl_n21) );
  INV_X1 U_refctl_U23 ( .A(U_refctl_N19), .ZN(U_refctl_n20) );
  AOI21_X1 U_refctl_U22 ( .B1(U_refctl_n84), .B2(U_refctl_N18), .A(
        U_refctl_n18), .ZN(U_refctl_n19) );
  AOI221_X1 U_refctl_U21 ( .B1(U_refctl_n14), .B2(U_refctl_n15), .C1(
        U_refctl_n16), .C2(U_refctl_n15), .A(U_refctl_n17), .ZN(U_refctl_n18)
         );
  OAI22_X1 U_refctl_U20 ( .A1(U_refctl_N17), .A2(U_refctl_n74), .B1(
        U_refctl_N18), .B2(U_refctl_n84), .ZN(U_refctl_n17) );
  OAI22_X1 U_refctl_U19 ( .A1(U_refctl_N16), .A2(U_refctl_n77), .B1(
        U_refctl_n73), .B2(U_refctl_n12), .ZN(U_refctl_n16) );
  AOI22_X1 U_refctl_U18 ( .A1(U_refctl_N17), .A2(U_refctl_n74), .B1(
        U_refctl_N16), .B2(U_refctl_n77), .ZN(U_refctl_n15) );
  AOI22_X1 U_refctl_U17 ( .A1(U_refctl_n73), .A2(U_refctl_n12), .B1(
        U_refctl_n83), .B2(n87), .ZN(U_refctl_n14) );
  INV_X1 U_refctl_U15 ( .A(U_refctl_n47), .ZN(U_refctl_n12) );
  NAND2_X1 U_refctl_U14 ( .A1(U_refctl_n118), .A2(U_refctl_count_7_), .ZN(
        U_refctl_n11) );
  OAI221_X1 U_refctl_U13 ( .B1(U_refctl_n5), .B2(U_refctl_n122), .C1(
        U_refctl_n5), .C2(U_refctl_n10), .A(ctl_ref_ack), .ZN(U_refctl_n124)
         );
  OAI21_X1 U_refctl_U12 ( .B1(U_refctl_n116), .B2(U_refctl_n7), .A(U_refctl_n9), .ZN(U_refctl_n10) );
  AOI21_X1 U_refctl_U11 ( .B1(U_refctl_N25), .B2(U_refctl_n80), .A(U_refctl_n8), .ZN(U_refctl_n9) );
  OAI21_X1 U_refctl_U10 ( .B1(U_refctl_n116), .B2(U_refctl_n115), .A(
        U_refctl_n114), .ZN(U_refctl_n8) );
  OAI21_X1 U_refctl_U9 ( .B1(U_refctl_N22), .B2(U_refctl_n87), .A(U_refctl_n6), 
        .ZN(U_refctl_n7) );
  OAI21_X1 U_refctl_U8 ( .B1(U_refctl_count_7_), .B2(U_refctl_n118), .A(
        U_refctl_n117), .ZN(U_refctl_n6) );
  OAI211_X1 U_refctl_U7 ( .C1(U_refctl_n120), .C2(U_refctl_n2), .A(U_refctl_n3), .B(U_refctl_n4), .ZN(U_refctl_n5) );
  OAI211_X1 U_refctl_U6 ( .C1(U_refctl_N29), .C2(U_refctl_n81), .A(
        U_refctl_N28), .B(U_refctl_n86), .ZN(U_refctl_n4) );
  AOI21_X1 U_refctl_U5 ( .B1(U_refctl_n81), .B2(U_refctl_N29), .A(U_refctl_N30), .ZN(U_refctl_n3) );
  AOI22_X1 U_refctl_U4 ( .A1(U_refctl_N27), .A2(U_refctl_n91), .B1(
        U_refctl_N26), .B2(U_refctl_n1), .ZN(U_refctl_n2) );
  NOR2_X1 U_refctl_U3 ( .A1(U_refctl_count_12_), .A2(U_refctl_n119), .ZN(
        U_refctl_n1) );
  DFFR_X1 U_refctl_count_reg_0_ ( .D(U_refctl_count_next_0_), .CK(hclk), .RN(
        hresetn), .Q(U_refctl_count_0_), .QN(U_refctl_n83) );
  DFFR_X1 U_refctl_count_reg_10_ ( .D(U_refctl_n79), .CK(hclk), .RN(hresetn), 
        .Q(U_refctl_count_10_), .QN(U_refctl_n90) );
  DFFR_X1 U_refctl_count_reg_11_ ( .D(U_refctl_count_next_11_), .CK(hclk), 
        .RN(hresetn), .Q(U_refctl_count_11_), .QN(U_refctl_n80) );
  DFFR_X1 U_refctl_count_reg_12_ ( .D(U_refctl_n82), .CK(hclk), .RN(hresetn), 
        .Q(U_refctl_count_12_) );
  DFFR_X1 U_refctl_count_reg_13_ ( .D(U_refctl_count_next_13_), .CK(hclk), 
        .RN(hresetn), .Q(U_refctl_count_13_), .QN(U_refctl_n91) );
  DFFR_X1 U_refctl_count_reg_14_ ( .D(U_refctl_count_next_14_), .CK(hclk), 
        .RN(hresetn), .Q(U_refctl_count_14_), .QN(U_refctl_n86) );
  DFFR_X1 U_refctl_count_reg_15_ ( .D(U_refctl_count_next_15_), .CK(hclk), 
        .RN(hresetn), .Q(U_refctl_count_15_), .QN(U_refctl_n81) );
  DFFR_X1 U_refctl_count_reg_1_ ( .D(U_refctl_count_next_1_), .CK(hclk), .RN(
        hresetn), .Q(U_refctl_count_1_), .QN(U_refctl_n73) );
  DFFR_X1 U_refctl_count_reg_2_ ( .D(U_refctl_count_next_2_), .CK(hclk), .RN(
        hresetn), .Q(U_refctl_count_2_), .QN(U_refctl_n77) );
  DFFR_X1 U_refctl_count_reg_3_ ( .D(U_refctl_count_next_3_), .CK(hclk), .RN(
        hresetn), .Q(U_refctl_count_3_), .QN(U_refctl_n74) );
  DFFR_X1 U_refctl_count_reg_4_ ( .D(U_refctl_count_next_4_), .CK(hclk), .RN(
        hresetn), .Q(U_refctl_count_4_), .QN(U_refctl_n84) );
  DFFR_X1 U_refctl_count_reg_5_ ( .D(U_refctl_count_next_5_), .CK(hclk), .RN(
        hresetn), .Q(U_refctl_count_5_), .QN(U_refctl_n85) );
  DFFR_X1 U_refctl_count_reg_6_ ( .D(U_refctl_n75), .CK(hclk), .RN(hresetn), 
        .Q(U_refctl_count_6_), .QN(U_refctl_n88) );
  DFFR_X1 U_refctl_count_reg_7_ ( .D(U_refctl_count_next_7_), .CK(hclk), .RN(
        hresetn), .Q(U_refctl_count_7_), .QN(U_refctl_n89) );
  DFFR_X1 U_refctl_count_reg_8_ ( .D(U_refctl_n76), .CK(hclk), .RN(hresetn), 
        .Q(U_refctl_count_8_), .QN(U_refctl_n87) );
  DFFR_X1 U_refctl_count_reg_9_ ( .D(U_refctl_count_next_9_), .CK(hclk), .RN(
        hresetn), .Q(U_refctl_count_9_), .QN(U_refctl_n78) );
  DFFR_X1 U_refctl_current_state_reg_1_ ( .D(U_refctl_ref_req_next), .CK(hclk), 
        .RN(hresetn), .Q(U_refctl_current_state_1_), .QN(U_refctl_n92) );
  DFFR_X1 U_refctl_ref_req_reg ( .D(U_refctl_ref_req_next), .CK(hclk), .RN(
        hresetn), .Q(debug_ref_req), .QN(n84) );
  DFFR_X1 U_refctl_current_state_reg_0_ ( .D(U_refctl_next_state_0_), .CK(hclk), .RN(hresetn), .Q(U_refctl_current_state_0_) );
  AND3_X4 U_dmc_U76 ( .A1(U_dmc_n63), .A2(U_dmc_n8), .A3(U_dmc_n19), .ZN(
        U_dmc_n52) );
  AND2_X4 U_dmc_U75 ( .A1(U_dmc_n62), .A2(U_dmc_n6), .ZN(U_dmc_n8) );
  NOR2_X2 U_dmc_U73 ( .A1(U_dmc_n70), .A2(U_dmc_n33), .ZN(U_dmc_n39) );
  AND4_X4 U_dmc_U72 ( .A1(U_dmc_terminate), .A2(hiu_wrapped_burst), .A3(
        U_dmc_n62), .A4(U_dmc_n63), .ZN(U_dmc_n12) );
  NOR3_X2 U_dmc_U69 ( .A1(U_dmc_data_cnt_4_), .A2(U_dmc_data_cnt_5_), .A3(
        U_dmc_n58), .ZN(U_dmc_n18) );
  NAND2_X2 U_dmc_U68 ( .A1(U_dmc_n63), .A2(U_dmc_n18), .ZN(U_dmc_n20) );
  NAND2_X2 U_dmc_U67 ( .A1(U_dmc_n20), .A2(U_dmc_n6), .ZN(U_dmc_n59) );
  NAND2_X2 U_dmc_U66 ( .A1(U_dmc_n4), .A2(U_dmc_dmc_cs_1_), .ZN(U_dmc_n15) );
  NOR2_X2 U_dmc_U65 ( .A1(U_dmc_n15), .A2(U_dmc_dmc_cs_2_), .ZN(U_dmc_n53) );
  INV_X4 U_dmc_U64 ( .A(U_dmc_n53), .ZN(U_dmc_n27) );
  NAND2_X2 U_dmc_U63 ( .A1(U_dmc_dmc_cs_1_), .A2(U_dmc_dmc_cs_0_), .ZN(
        U_dmc_n10) );
  NOR2_X2 U_dmc_U62 ( .A1(U_dmc_n10), .A2(U_dmc_dmc_cs_2_), .ZN(U_dmc_n55) );
  AOI211_X2 U_dmc_U61 ( .C1(U_dmc_n25), .C2(U_dmc_n24), .A(U_dmc_n23), .B(
        hiu_terminate), .ZN(U_dmc_n30) );
  NAND2_X2 U_dmc_U60 ( .A1(U_dmc_n7), .A2(U_dmc_dmc_cs_0_), .ZN(U_dmc_n11) );
  NOR2_X2 U_dmc_U59 ( .A1(U_dmc_n11), .A2(U_dmc_dmc_cs_2_), .ZN(U_dmc_n54) );
  OAI211_X2 U_dmc_U58 ( .C1(U_dmc_n32), .C2(U_dmc_n27), .A(U_dmc_n30), .B(
        U_dmc_n26), .ZN(U_dmc_N23) );
  INV_X4 U_dmc_U57 ( .A(U_dmc_n54), .ZN(U_dmc_n31) );
  OAI211_X2 U_dmc_U56 ( .C1(U_dmc_n32), .C2(U_dmc_n31), .A(U_dmc_n30), .B(
        U_dmc_n29), .ZN(U_dmc_N24) );
  NAND2_X2 U_dmc_U55 ( .A1(U_dmc_n4), .A2(U_dmc_n7), .ZN(U_dmc_n61) );
  NAND2_X2 U_dmc_U54 ( .A1(U_dmc_n31), .A2(U_dmc_n27), .ZN(U_dmc_n62) );
  AOI22_X2 U_dmc_U53 ( .A1(U_dmc_terminate), .A2(U_dmc_n55), .B1(U_dmc_n62), 
        .B2(U_dmc_n59), .ZN(U_dmc_n60) );
  AOI21_X2 U_dmc_U51 ( .B1(N28), .B2(U_dmc_n25), .A(U_dmc_n21), .ZN(U_dmc_n70)
         );
  NAND2_X2 U_dmc_U50 ( .A1(U_dmc_n35), .A2(U_dmc_n34), .ZN(U_dmc_n48) );
  NOR2_X2 U_dmc_U49 ( .A1(U_dmc_n51), .A2(U_dmc_n48), .ZN(U_dmc_n47) );
  NAND2_X2 U_dmc_U47 ( .A1(U_dmc_n47), .A2(U_dmc_n45), .ZN(U_dmc_n46) );
  NOR2_X2 U_dmc_U45 ( .A1(U_dmc_n46), .A2(U_dmc_n43), .ZN(U_dmc_n42) );
  NAND2_X2 U_dmc_U44 ( .A1(U_dmc_n42), .A2(U_dmc_n40), .ZN(U_dmc_n41) );
  NOR2_X2 U_dmc_U43 ( .A1(U_dmc_n39), .A2(U_dmc_n52), .ZN(U_dmc_n50) );
  AOI21_X2 U_dmc_U42 ( .B1(U_dmc_n43), .B2(U_dmc_n46), .A(U_dmc_n42), .ZN(
        U_dmc_n44) );
  NOR2_X2 U_dmc_U41 ( .A1(U_dmc_n44), .A2(U_dmc_n50), .ZN(
        U_dmc_data_cnt_nxt[3]) );
  AOI21_X2 U_dmc_U40 ( .B1(U_dmc_n51), .B2(U_dmc_n48), .A(U_dmc_n47), .ZN(
        U_dmc_n49) );
  NOR2_X2 U_dmc_U39 ( .A1(U_dmc_n49), .A2(U_dmc_n50), .ZN(
        U_dmc_data_cnt_nxt[1]) );
  NAND3_X2 U_dmc_U38 ( .A1(U_dmc_n8), .A2(hiu_wrapped_burst), .A3(U_dmc_n64), 
        .ZN(U_dmc_n69) );
  AOI21_X2 U_dmc_U37 ( .B1(U_dmc_n54), .B2(U_dmc_n66), .A(U_dmc_n52), .ZN(
        U_dmc_n67) );
  AOI21_X1 U_dmc_U36 ( .B1(hiu_rw), .B2(U_dmc_n28), .A(U_dmc_n54), .ZN(
        U_dmc_n26) );
  INV_X1 U_dmc_U35 ( .A(U_dmc_n18), .ZN(U_dmc_n19) );
  AOI22_X2 U_dmc_U34 ( .A1(U_dmc_n39), .A2(hiu_burst_size[4]), .B1(
        U_dmc_data_cnt_4_), .B2(U_dmc_n52), .ZN(U_dmc_n40) );
  INV_X1 U_dmc_U33 ( .A(U_dmc_n20), .ZN(U_dmc_n64) );
  OAI211_X1 U_dmc_U32 ( .C1(U_dmc_n70), .C2(hiu_rw), .A(U_dmc_n65), .B(
        U_dmc_n69), .ZN(U_dmc_n13) );
  INV_X1 U_dmc_U31 ( .A(U_dmc_n59), .ZN(U_dmc_n32) );
  INV_X1 U_dmc_U30 ( .A(U_dmc_n63), .ZN(U_dmc_n33) );
  NOR3_X1 U_dmc_U29 ( .A1(U_dmc_dmc_cs_2_), .A2(U_dmc_dmc_cs_1_), .A3(
        U_dmc_dmc_cs_0_), .ZN(U_dmc_n25) );
  OR4_X2 U_dmc_U28 ( .A1(U_dmc_data_cnt_1_), .A2(U_dmc_data_cnt_2_), .A3(
        U_dmc_data_cnt_0_), .A4(U_dmc_data_cnt_3_), .ZN(U_dmc_n58) );
  INV_X1 U_dmc_U27 ( .A(U_dmc_n55), .ZN(U_dmc_n22) );
  NOR2_X1 U_dmc_U26 ( .A1(U_dmc_n22), .A2(U_dmc_terminate), .ZN(U_dmc_n21) );
  OAI21_X1 U_dmc_U25 ( .B1(U_dmc_n22), .B2(U_dmc_n6), .A(U_dmc_n5), .ZN(
        U_dmc_n23) );
  AOI21_X1 U_dmc_U24 ( .B1(U_dsdc_n1438), .B2(U_dmc_n28), .A(U_dmc_n53), .ZN(
        U_dmc_n29) );
  AOI22_X1 U_dmc_U22 ( .A1(U_dmc_dmc_cs_1_), .A2(U_dmc_n52), .B1(U_dmc_n53), 
        .B2(U_dmc_n66), .ZN(U_dmc_n65) );
  NAND2_X1 U_dmc_U21 ( .A1(U_dmc_n52), .A2(U_dmc_data_cnt_1_), .ZN(U_dmc_n34)
         );
  OR2_X1 U_dmc_U18 ( .A1(U_dmc_n4), .A2(U_dmc_n67), .ZN(U_dmc_n68) );
  INV_X2 U_dmc_U17 ( .A(N28), .ZN(U_dmc_n24) );
  NAND2_X1 U_dmc_U15 ( .A1(U_dmc_n39), .A2(hiu_burst_size[1]), .ZN(U_dmc_n35)
         );
  NOR2_X1 U_dmc_U14 ( .A1(U_dmc_n51), .A2(U_dmc_n50), .ZN(
        U_dmc_data_cnt_nxt[0]) );
  OR2_X1 U_dmc_U13 ( .A1(U_dmc_n25), .A2(U_dmc_n55), .ZN(U_dmc_n28) );
  INV_X4 U_dmc_U12 ( .A(hiu_burst_size[4]), .ZN(U_dmc_n16) );
  NOR2_X1 U_dmc_U11 ( .A1(U_dmc_terminate), .A2(U_dmc_n63), .ZN(U_dmc_n66) );
  OAI211_X1 U_dmc_U10 ( .C1(U_dmc_n70), .C2(U_dsdc_n1438), .A(U_dmc_n69), .B(
        U_dmc_n68), .ZN(U_dmc_n14) );
  AOI221_X1 U_dmc_U9 ( .B1(U_dmc_n47), .B2(U_dmc_n46), .C1(U_dmc_n45), .C2(
        U_dmc_n46), .A(U_dmc_n50), .ZN(U_dmc_data_cnt_nxt[2]) );
  AOI221_X1 U_dmc_U8 ( .B1(U_dmc_n42), .B2(U_dmc_n41), .C1(U_dmc_n40), .C2(
        U_dmc_n41), .A(U_dmc_n50), .ZN(U_dmc_data_cnt_nxt[4]) );
  AOI211_X1 U_dmc_U7 ( .C1(U_dmc_n41), .C2(U_dmc_n2), .A(U_dmc_n50), .B(
        U_dmc_n3), .ZN(U_dmc_data_cnt_nxt[5]) );
  NOR2_X1 U_dmc_U6 ( .A1(U_dmc_n41), .A2(U_dmc_n2), .ZN(U_dmc_n3) );
  AOI22_X1 U_dmc_U5 ( .A1(U_dmc_n52), .A2(U_dmc_data_cnt_5_), .B1(
        hiu_burst_size[5]), .B2(U_dmc_n39), .ZN(U_dmc_n2) );
  INV_X1 U_dmc_U4 ( .A(U_dmc_n1), .ZN(U_dmc_n51) );
  AOI22_X1 U_dmc_U3 ( .A1(hiu_burst_size[0]), .A2(U_dmc_n39), .B1(
        U_dmc_data_cnt_0_), .B2(U_dmc_n52), .ZN(U_dmc_n1) );
  DFFR_X2 U_dmc_terminate_reg ( .D(hiu_terminate), .CK(hclk), .RN(hresetn), 
        .Q(U_dmc_terminate), .QN(U_dmc_n6) );
  DFFR_X2 U_dmc_dmc_cs_reg_0_ ( .D(U_dmc_n14), .CK(hclk), .RN(hresetn), .Q(
        U_dmc_dmc_cs_0_), .QN(U_dmc_n4) );
  DFFR_X2 U_dmc_dmc_cs_reg_1_ ( .D(U_dmc_n13), .CK(hclk), .RN(hresetn), .Q(
        U_dmc_dmc_cs_1_), .QN(U_dmc_n7) );
  DFFR_X2 U_dmc_dmc_cs_reg_2_ ( .D(U_dmc_n12), .CK(hclk), .RN(hresetn), .Q(
        U_dmc_dmc_cs_2_), .QN(U_dmc_n5) );
  DFFS_X2 U_dmc_miu_pop_n_reg ( .D(U_dmc_N23), .CK(hclk), .SN(hresetn), .Q(
        dmc_pop_n) );
  DFFS_X2 U_dmc_miu_push_n_reg ( .D(U_dmc_N24), .CK(hclk), .SN(hresetn), .Q(
        dmc_push_n) );
  DFFR_X1 U_dmc_data_cnt_reg_5_ ( .D(U_dmc_data_cnt_nxt[5]), .CK(hclk), .RN(
        hresetn), .Q(U_dmc_data_cnt_5_) );
  DFFR_X1 U_dmc_data_cnt_reg_4_ ( .D(U_dmc_data_cnt_nxt[4]), .CK(hclk), .RN(
        hresetn), .Q(U_dmc_data_cnt_4_) );
  DFFR_X1 U_dmc_data_cnt_reg_3_ ( .D(U_dmc_data_cnt_nxt[3]), .CK(hclk), .RN(
        hresetn), .Q(U_dmc_data_cnt_3_) );
  DFFR_X1 U_dmc_data_cnt_reg_2_ ( .D(U_dmc_data_cnt_nxt[2]), .CK(hclk), .RN(
        hresetn), .Q(U_dmc_data_cnt_2_) );
  DFFR_X1 U_dmc_data_cnt_reg_1_ ( .D(U_dmc_data_cnt_nxt[1]), .CK(hclk), .RN(
        hresetn), .Q(U_dmc_data_cnt_1_) );
  DFFR_X1 U_dmc_data_cnt_reg_0_ ( .D(U_dmc_data_cnt_nxt[0]), .CK(hclk), .RN(
        hresetn), .Q(U_dmc_data_cnt_0_) );
  NAND2_X2 U_dsdc_U_minmax1_dwbb_U40 ( .A1(U_dsdc_U_minmax1_dwbb_n26), .A2(
        U_dsdc_U_minmax1_dwbb_n2), .ZN(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_1_) );
  NAND4_X2 U_dsdc_U_minmax1_dwbb_U39 ( .A1(U_dsdc_U_minmax1_dwbb_n22), .A2(
        U_dsdc_U_minmax1_dwbb_n21), .A3(U_dsdc_U_minmax1_dwbb_n20), .A4(
        U_dsdc_U_minmax1_dwbb_n19), .ZN(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_0_) );
  MUX2_X2 U_dsdc_U_minmax1_dwbb_U37 ( .A(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_), .B(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_), .S(
        U_dsdc_oldest_bank_1_), .Z(U_dsdc_oldest_bank_0_) );
  OR2_X1 U_dsdc_U_minmax1_dwbb_U32 ( .A1(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_), .A2(
        U_dsdc_bm_bank_age_0__0_), .ZN(U_dsdc_U_minmax1_dwbb_n21) );
  NAND2_X1 U_dsdc_U_minmax1_dwbb_U31 ( .A1(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_), .A2(U_dsdc_n352), 
        .ZN(U_dsdc_U_minmax1_dwbb_n20) );
  NAND2_X1 U_dsdc_U_minmax1_dwbb_U30 ( .A1(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_), .A2(
        U_dsdc_bm_bank_age_3__0_), .ZN(U_dsdc_U_minmax1_dwbb_n19) );
  NAND2_X1 U_dsdc_U_minmax1_dwbb_U29 ( .A1(U_dsdc_U_minmax1_dwbb_n24), .A2(
        U_dsdc_bm_bank_age_2__0_), .ZN(U_dsdc_U_minmax1_dwbb_n22) );
  AND2_X2 U_dsdc_U_minmax1_dwbb_U28 ( .A1(U_dsdc_U_minmax1_dwbb_n33), .A2(
        U_dsdc_U_minmax1_dwbb_n31), .ZN(U_dsdc_U_minmax1_dwbb_n32) );
  OR2_X2 U_dsdc_U_minmax1_dwbb_U27 ( .A1(U_dsdc_U_minmax1_dwbb_n33), .A2(
        U_dsdc_U_minmax1_dwbb_n31), .ZN(U_dsdc_U_minmax1_dwbb_n34) );
  INV_X2 U_dsdc_U_minmax1_dwbb_U26 ( .A(U_dsdc_U_minmax1_dwbb_n30), .ZN(
        U_dsdc_U_minmax1_dwbb_n26) );
  AND2_X2 U_dsdc_U_minmax1_dwbb_U25 ( .A1(U_dsdc_U_minmax1_dwbb_n30), .A2(
        U_dsdc_U_minmax1_dwbb_n29), .ZN(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_PI_1_) );
  INV_X1 U_dsdc_U_minmax1_dwbb_U22 ( .A(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_), .ZN(
        U_dsdc_U_minmax1_dwbb_n24) );
  OAI21_X1 U_dsdc_U_minmax1_dwbb_U21 ( .B1(U_dsdc_bm_bank_age_2__2_), .B2(
        U_dsdc_n303), .A(U_dsdc_U_minmax1_dwbb_n15), .ZN(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_) );
  OAI211_X1 U_dsdc_U_minmax1_dwbb_U20 ( .C1(U_dsdc_bm_bank_age_3__2_), .C2(
        U_dsdc_n336), .A(U_dsdc_U_minmax1_dwbb_n12), .B(
        U_dsdc_U_minmax1_dwbb_n11), .ZN(U_dsdc_U_minmax1_dwbb_n15) );
  NAND2_X1 U_dsdc_U_minmax1_dwbb_U17 ( .A1(U_dsdc_bm_bank_age_2__1_), .A2(
        U_dsdc_n302), .ZN(U_dsdc_U_minmax1_dwbb_n12) );
  OAI211_X1 U_dsdc_U_minmax1_dwbb_U16 ( .C1(U_dsdc_bm_bank_age_2__1_), .C2(
        U_dsdc_n302), .A(U_dsdc_n304), .B(U_dsdc_bm_bank_age_2__0_), .ZN(
        U_dsdc_U_minmax1_dwbb_n11) );
  AOI22_X1 U_dsdc_U_minmax1_dwbb_U15 ( .A1(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_), .A2(
        U_dsdc_bm_bank_age_3__2_), .B1(U_dsdc_bm_bank_age_2__2_), .B2(
        U_dsdc_U_minmax1_dwbb_n24), .ZN(U_dsdc_U_minmax1_dwbb_n33) );
  OAI21_X1 U_dsdc_U_minmax1_dwbb_U13 ( .B1(U_dsdc_bm_bank_age_0__2_), .B2(
        U_dsdc_n337), .A(U_dsdc_U_minmax1_dwbb_n9), .ZN(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_) );
  OAI211_X1 U_dsdc_U_minmax1_dwbb_U12 ( .C1(U_dsdc_bm_bank_age_1__2_), .C2(
        U_dsdc_n334), .A(U_dsdc_U_minmax1_dwbb_n6), .B(
        U_dsdc_U_minmax1_dwbb_n5), .ZN(U_dsdc_U_minmax1_dwbb_n9) );
  NAND2_X1 U_dsdc_U_minmax1_dwbb_U9 ( .A1(U_dsdc_bm_bank_age_0__1_), .A2(
        U_dsdc_n335), .ZN(U_dsdc_U_minmax1_dwbb_n6) );
  OAI211_X1 U_dsdc_U_minmax1_dwbb_U8 ( .C1(U_dsdc_bm_bank_age_0__1_), .C2(
        U_dsdc_n335), .A(U_dsdc_n352), .B(U_dsdc_bm_bank_age_0__0_), .ZN(
        U_dsdc_U_minmax1_dwbb_n5) );
  AOI22_X2 U_dsdc_U_minmax1_dwbb_U7 ( .A1(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_), .A2(
        U_dsdc_bm_bank_age_1__1_), .B1(U_dsdc_bm_bank_age_0__1_), .B2(
        U_dsdc_U_minmax1_dwbb_n4), .ZN(U_dsdc_U_minmax1_dwbb_n30) );
  INV_X4 U_dsdc_U_minmax1_dwbb_U6 ( .A(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_), .ZN(
        U_dsdc_U_minmax1_dwbb_n4) );
  INV_X1 U_dsdc_U_minmax1_dwbb_U4 ( .A(U_dsdc_U_minmax1_dwbb_n2), .ZN(
        U_dsdc_U_minmax1_dwbb_n29) );
  AOI22_X1 U_dsdc_U_minmax1_dwbb_U3 ( .A1(U_dsdc_bm_bank_age_2__1_), .A2(
        U_dsdc_U_minmax1_dwbb_n24), .B1(U_dsdc_bm_bank_age_3__1_), .B2(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_1_prefix_GT_8_), .ZN(
        U_dsdc_U_minmax1_dwbb_n2) );
  OAI21_X2 U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_UGT1_1_0_0 ( .B1(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_PI_1_), .B2(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_0_), .A(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_GI_1_), .ZN(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_GT_4_) );
  AOI21_X2 U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_UGT0_2_0_0 ( .B1(
        U_dsdc_U_minmax1_dwbb_n34), .B2(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_1_0_prefix_GT_4_), .A(
        U_dsdc_U_minmax1_dwbb_n32), .ZN(U_dsdc_oldest_bank_1_) );
  OAI33_X1 U17 ( .A1(U_dsdc_n165), .A2(U_dsdc_n903), .A3(U_dsdc_n934), .B1(
        U_dsdc_n740), .B2(U_dsdc_n739), .B3(U_dsdc_n741), .ZN(n45) );
  INV_X4 U22 ( .A(n45), .ZN(U_dsdc_n744) );
  AOI22_X1 U23 ( .A1(hiu_burst_size[2]), .A2(U_dmc_n39), .B1(U_dmc_data_cnt_2_), .B2(U_dmc_n52), .ZN(U_dmc_n45) );
  OAI22_X1 U28 ( .A1(U_dsdc_n1424), .A2(U_dsdc_n1628), .B1(U_dsdc_n1426), .B2(
        U_dsdc_n1421), .ZN(n46) );
  NOR3_X1 U46 ( .A1(U_dsdc_n1872), .A2(U_dsdc_n967), .A3(n46), .ZN(n47) );
  INV_X1 U47 ( .A(U_dsdc_n1591), .ZN(n48) );
  NAND3_X1 U57 ( .A1(U_dsdc_n705), .A2(n47), .A3(n48), .ZN(U_dsdc_n1383) );
  AOI22_X2 U58 ( .A1(U_addrdec_n39), .A2(hiu_addr[13]), .B1(U_addrdec_n220), 
        .B2(hiu_addr[14]), .ZN(debug_ad_col_addr_13_) );
  NOR4_X1 U59 ( .A1(hiu_burst_size[2]), .A2(hiu_burst_size[3]), .A3(
        hiu_burst_size[0]), .A4(hiu_burst_size[1]), .ZN(n49) );
  INV_X1 U60 ( .A(hiu_burst_size[5]), .ZN(n50) );
  NAND3_X1 U61 ( .A1(U_dmc_n16), .A2(n49), .A3(n50), .ZN(U_dmc_n63) );
  NOR4_X2 U62 ( .A1(U_dsdc_r_burst_size_4_), .A2(U_dsdc_r_burst_size_3_), .A3(
        U_dsdc_r_burst_size_5_), .A4(U_dsdc_r_burst_size_0_), .ZN(n51) );
  NAND2_X1 U63 ( .A1(U_dsdc_n687), .A2(n51), .ZN(U_dsdc_n1312) );
  NAND2_X1 U64 ( .A1(U_dsdc_n1284), .A2(hiu_rw), .ZN(n52) );
  NOR3_X1 U65 ( .A1(n52), .A2(U_dsdc_n1286), .A3(U_dsdc_n1053), .ZN(
        U_dsdc_n1124) );
  AOI22_X2 U66 ( .A1(U_addrdec_n220), .A2(hiu_addr[10]), .B1(U_addrdec_n39), 
        .B2(hiu_addr[9]), .ZN(n53) );
  INV_X4 U67 ( .A(n53), .ZN(debug_ad_col_addr_9_) );
  AOI22_X2 U68 ( .A1(U_addrdec_n220), .A2(hiu_addr[15]), .B1(U_addrdec_n39), 
        .B2(hiu_addr[14]), .ZN(n54) );
  INV_X4 U69 ( .A(n54), .ZN(debug_ad_col_addr_14_) );
  AOI22_X2 U70 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__0_), .B1(
        U_dsdc_bm_row_addr_0__0_), .B2(U_dsdc_n998), .ZN(U_dsdc_n558) );
  AOI22_X1 U71 ( .A1(hiu_burst_size[3]), .A2(U_dmc_n39), .B1(U_dmc_data_cnt_3_), .B2(U_dmc_n52), .ZN(n55) );
  INV_X1 U72 ( .A(n55), .ZN(U_dmc_n43) );
  AND2_X1 U73 ( .A1(U_dsdc_n1254), .A2(U_dsdc_n1253), .ZN(n56) );
  OAI221_X1 U74 ( .B1(n56), .B2(U_dsdc_n1546), .C1(n56), .C2(U_dsdc_n2013), 
        .A(U_dsdc_n1409), .ZN(U_dsdc_n1270) );
  AOI211_X1 U75 ( .C1(U_dsdc_n1876), .C2(U_dsdc_n1416), .A(U_dsdc_n1412), .B(
        U_dsdc_n1872), .ZN(n57) );
  OAI211_X1 U76 ( .C1(U_dsdc_n1414), .C2(U_dsdc_n2071), .A(U_dsdc_n705), .B(
        n57), .ZN(n58) );
  OAI21_X1 U77 ( .B1(U_dsdc_n991), .B2(U_dsdc_n856), .A(U_dsdc_n2072), .ZN(n59) );
  AOI211_X1 U78 ( .C1(U_dsdc_n721), .C2(U_dsdc_n708), .A(n58), .B(n59), .ZN(
        U_dsdc_n183) );
  AOI22_X2 U79 ( .A1(U_addrdec_n220), .A2(hiu_addr[11]), .B1(U_addrdec_n39), 
        .B2(hiu_addr[10]), .ZN(n60) );
  INV_X4 U80 ( .A(n60), .ZN(debug_ad_col_addr_10_) );
  AOI222_X2 U81 ( .A1(U_dsdc_n604), .A2(U_dsdc_bm_row_addr_1__3_), .B1(
        U_dsdc_n978), .B2(U_dsdc_bm_row_addr_3__3_), .C1(U_dsdc_n159), .C2(
        U_dsdc_bm_row_addr_2__3_), .ZN(n61) );
  INV_X1 U82 ( .A(n61), .ZN(U_dsdc_n798) );
  AOI22_X1 U83 ( .A1(U_dsdc_U_minmax1_dwbb_n4), .A2(U_dsdc_bm_bank_age_0__2_), 
        .B1(U_dsdc_bm_bank_age_1__2_), .B2(
        U_dsdc_U_minmax1_dwbb_U1_minmax2_0_0_prefix_GT_8_), .ZN(n62) );
  INV_X1 U84 ( .A(n62), .ZN(U_dsdc_U_minmax1_dwbb_n31) );
  OAI21_X2 U85 ( .B1(U_dsdc_n1945), .B2(U_dsdc_n1836), .A(U_dsdc_n1837), .ZN(
        n63) );
  AOI222_X1 U86 ( .A1(U_dsdc_n1953), .A2(U_dsdc_bm_bank_age_2__3_), .B1(
        U_dsdc_n1953), .B2(n63), .C1(U_dsdc_bm_bank_age_2__3_), .C2(n63), .ZN(
        n64) );
  AOI222_X2 U87 ( .A1(U_dsdc_n1954), .A2(U_dsdc_n350), .B1(U_dsdc_n1954), .B2(
        n64), .C1(U_dsdc_n350), .C2(n64), .ZN(U_dsdc_n1849) );
  AOI22_X2 U88 ( .A1(U_addrdec_n220), .A2(hiu_addr[16]), .B1(U_addrdec_n39), 
        .B2(hiu_addr[15]), .ZN(n65) );
  INV_X4 U89 ( .A(n65), .ZN(debug_ad_col_addr_15_) );
  NAND3_X1 U90 ( .A1(U_dsdc_n1393), .A2(U_dsdc_cas_latency_cnt_0_), .A3(
        U_dsdc_cas_latency_cnt_1_), .ZN(n66) );
  INV_X1 U91 ( .A(U_dsdc_n1393), .ZN(n67) );
  NAND2_X1 U92 ( .A1(U_dsdc_cas_latency_1_), .A2(n67), .ZN(n68) );
  OAI211_X1 U93 ( .C1(U_dsdc_n1090), .C2(U_dsdc_n1087), .A(n66), .B(n68), .ZN(
        U_dsdc_N4127) );
  OAI33_X1 U94 ( .A1(U_dsdc_n815), .A2(U_dsdc_bm_row_addr_0__1_), .A3(
        U_dsdc_n814), .B1(U_addrdec_n231), .B2(U_dsdc_n812), .B3(
        U_dsdc_bm_row_addr_0__11_), .ZN(n69) );
  INV_X1 U95 ( .A(n69), .ZN(U_dsdc_n536) );
  OAI211_X1 U96 ( .C1(U_dsdc_n602), .C2(U_dsdc_n816), .A(U_dsdc_n488), .B(
        U_dsdc_n51), .ZN(n70) );
  INV_X1 U97 ( .A(n70), .ZN(U_dsdc_n499) );
  NAND2_X1 U98 ( .A1(U_dsdc_r_cas_latency_3_), .A2(U_dsdc_n753), .ZN(n71) );
  XNOR2_X1 U99 ( .A(n71), .B(U_dsdc_DP_OP_1642_126_2028_n85), .ZN(
        U_dsdc_DP_OP_1642_126_2028_n19) );
  INV_X1 U100 ( .A(U_cr_n65), .ZN(n72) );
  AOI21_X1 U101 ( .B1(U_addrdec_n67), .B2(n72), .A(U_addrdec_n74), .ZN(
        U_addrdec_n75) );
  OAI21_X1 U102 ( .B1(U_dsdc_bm_bank_age_0__1_), .B2(U_dsdc_n1948), .A(
        U_dsdc_n1947), .ZN(n73) );
  OAI21_X1 U103 ( .B1(U_dsdc_n1951), .B2(U_dsdc_n334), .A(n73), .ZN(n74) );
  AOI222_X1 U104 ( .A1(U_dsdc_bm_bank_age_0__3_), .A2(U_dsdc_n1953), .B1(
        U_dsdc_bm_bank_age_0__3_), .B2(n74), .C1(U_dsdc_n1953), .C2(n74), .ZN(
        n75) );
  AOI222_X1 U105 ( .A1(U_dsdc_n1954), .A2(U_dsdc_n434), .B1(U_dsdc_n1954), 
        .B2(n75), .C1(U_dsdc_n434), .C2(n75), .ZN(U_dsdc_n2080) );
  OR2_X1 U106 ( .A1(U_dsdc_n1805), .A2(U_dsdc_n1359), .ZN(n76) );
  NAND4_X1 U107 ( .A1(U_dsdc_n1342), .A2(U_dsdc_n1978), .A3(U_dsdc_n1368), 
        .A4(n76), .ZN(n89) );
  NAND3_X1 U108 ( .A1(U_dsdc_n1393), .A2(U_dsdc_n1087), .A3(
        U_dsdc_cas_latency_cnt_2_), .ZN(n77) );
  INV_X1 U109 ( .A(U_dsdc_n1393), .ZN(n78) );
  NAND2_X1 U110 ( .A1(U_dsdc_cas_latency_2_), .A2(n78), .ZN(n79) );
  OAI211_X1 U111 ( .C1(U_dsdc_n1094), .C2(U_dsdc_n1090), .A(n77), .B(n79), 
        .ZN(U_dsdc_N4128) );
  OAI21_X1 U112 ( .B1(U_dmc_n5), .B2(U_dmc_n61), .A(U_dmc_n60), .ZN(n80) );
  NOR2_X1 U113 ( .A1(ctl_burst_done), .A2(n80), .ZN(n81) );
  OAI211_X1 U114 ( .C1(U_cr_n503), .C2(U_cr_n502), .A(U_cr_n197), .B(n81), 
        .ZN(miu_burst_done) );
  OAI21_X4 U115 ( .B1(U_dsdc_n1024), .B2(U_dsdc_n1023), .A(
        U_dsdc_bm_num_open_bank_4_), .ZN(U_dsdc_n1025) );
  AOI21_X4 U116 ( .B1(U_dsdc_n159), .B2(U_dsdc_bm_row_addr_2__0_), .A(
        U_dsdc_n560), .ZN(U_dsdc_n561) );
  OAI211_X4 U117 ( .C1(U_addrdec_n73), .C2(U_cr_n65), .A(U_addrdec_n71), .B(
        U_addrdec_n70), .ZN(debug_ad_bank_addr[0]) );
  NAND2_X1 U118 ( .A1(U_dsdc_n981), .A2(U_dsdc_n979), .ZN(U_dsdc_n913) );
  NAND2_X1 U119 ( .A1(debug_ad_bank_addr[1]), .A2(debug_ad_bank_addr[0]), .ZN(
        U_dsdc_n987) );
  AOI22_X1 U120 ( .A1(U_addrdec_n220), .A2(hiu_addr[2]), .B1(hiu_addr[1]), 
        .B2(U_addrdec_n39), .ZN(U_addrdec_n96) );
  AOI22_X1 U121 ( .A1(U_addrdec_n220), .A2(hiu_addr[5]), .B1(hiu_addr[4]), 
        .B2(U_addrdec_n39), .ZN(U_addrdec_n97) );
  AOI22_X1 U122 ( .A1(U_addrdec_n220), .A2(hiu_addr[7]), .B1(hiu_addr[6]), 
        .B2(U_addrdec_n39), .ZN(U_addrdec_n99) );
  AOI22_X1 U123 ( .A1(U_addrdec_n220), .A2(hiu_addr[6]), .B1(hiu_addr[5]), 
        .B2(U_addrdec_n39), .ZN(U_addrdec_n98) );
  NOR2_X2 U124 ( .A1(U_dsdc_n537), .A2(U_dsdc_n333), .ZN(U_dsdc_n538) );
  OAI211_X2 U125 ( .C1(n[24]), .C2(U_addrdec_n84), .A(U_addrdec_n83), .B(
        U_addrdec_n82), .ZN(U_addrdec_n85) );
  INV_X16 U126 ( .A(n14), .ZN(debug_ad_bank_addr[1]) );
  INV_X16 U127 ( .A(n18), .ZN(n16) );
  INV_X4 U128 ( .A(big_endian), .ZN(U_addrdec_n40) );
  NAND2_X4 U129 ( .A1(U_dsdc_n1166), .A2(U_dsdc_n998), .ZN(n83) );
  INV_X4 U130 ( .A(U_dsdc_n601), .ZN(U_dsdc_DP_OP_1642_126_2028_n85) );
  AND2_X4 U131 ( .A1(U_dsdc_bm_row_addr_1__8_), .A2(U_dsdc_n604), .ZN(n86) );
  NAND2_X2 U132 ( .A1(U_dsdc_i_dqs), .A2(U_dsdc_i_dqs_d), .ZN(n88) );
endmodule


module DW_memctl ( hready_resp, hresp, hrdata, s_ras_n, s_cas_n, s_cke, 
        s_wr_data, s_addr, s_bank_addr, s_dout_valid, s_sel_n, s_dqm, s_we_n, 
        s_dqs, s_sa, s_scl, s_rd_ready, s_rd_start, s_rd_pop, s_rd_end, 
        s_rd_dqs_mask, s_cas_latency, s_read_pipe, s_sda_out, s_sda_oe_n, gpo, 
        debug_ad_bank_addr, debug_ad_row_addr, debug_ad_col_addr, 
        debug_ad_sf_bank_addr, debug_ad_sf_row_addr, debug_ad_sf_col_addr, 
        debug_hiu_addr, debug_sm_burst_done, debug_sm_pop_n, debug_sm_push_n, 
        debug_smc_cs, debug_ref_req, hclk, hclk_2x, hresetn, scan_mode, haddr, 
        hsel_mem, hsel_reg, hwrite, htrans, hsize, hburst, hready, hwdata, 
        s_rd_data, s_sda_in, gpi, remap, power_down, clear_sr_dp, big_endian
 );
  output [1:0] hresp;
  output [31:0] hrdata;
  output [15:0] s_wr_data;
  output [15:0] s_addr;
  output [1:0] s_bank_addr;
  output [1:0] s_dout_valid;
  output [0:0] s_sel_n;
  output [1:0] s_dqm;
  output [1:0] s_dqs;
  output [2:0] s_sa;
  output [2:0] s_cas_latency;
  output [2:0] s_read_pipe;
  output [7:0] gpo;
  output [1:0] debug_ad_bank_addr;
  output [15:0] debug_ad_row_addr;
  output [15:0] debug_ad_col_addr;
  output [1:0] debug_ad_sf_bank_addr;
  output [15:0] debug_ad_sf_row_addr;
  output [15:0] debug_ad_sf_col_addr;
  output [31:0] debug_hiu_addr;
  output [3:0] debug_smc_cs;
  input [31:0] haddr;
  input [1:0] htrans;
  input [2:0] hsize;
  input [2:0] hburst;
  input [31:0] hwdata;
  input [31:0] s_rd_data;
  input [7:0] gpi;
  input s_rd_ready, hclk, hclk_2x, hresetn, scan_mode, hsel_mem, hsel_reg,
         hwrite, hready, s_sda_in, remap, power_down, clear_sr_dp, big_endian;
  output hready_resp, s_ras_n, s_cas_n, s_cke, s_we_n, s_scl, s_rd_start,
         s_rd_pop, s_rd_end, s_rd_dqs_mask, s_sda_out, s_sda_oe_n,
         debug_sm_burst_done, debug_sm_pop_n, debug_sm_push_n, debug_ref_req;
  wire   hiu_wrap_burst, hiu_rw, hiu_terminate, miu_burst_done, miu_pop_n,
         miu_push_n, n2, n3, n4, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135,
         SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137,
         SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139,
         SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141,
         SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143,
         SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145,
         SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147,
         SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149,
         SYNOPSYS_UNCONNECTED_150;
  wire   [1:0] hiu_req;
  wire   [5:0] hiu_burst_size;
  wire   [31:0] hiu_data;
  wire   [3:0] hiu_haddr;
  wire   [2:0] hiu_hsize;
  wire   [31:0] miu_data;
  assign debug_smc_cs[0] = 1'b0;
  assign debug_smc_cs[1] = 1'b0;
  assign debug_smc_cs[2] = 1'b0;
  assign debug_smc_cs[3] = 1'b0;
  assign debug_sm_push_n = 1'b0;
  assign debug_sm_pop_n = 1'b0;
  assign debug_sm_burst_done = 1'b0;
  assign debug_hiu_addr[0] = 1'b0;
  assign debug_ad_sf_col_addr[0] = 1'b0;
  assign debug_ad_sf_col_addr[1] = 1'b0;
  assign debug_ad_sf_col_addr[2] = 1'b0;
  assign debug_ad_sf_col_addr[3] = 1'b0;
  assign debug_ad_sf_col_addr[4] = 1'b0;
  assign debug_ad_sf_col_addr[5] = 1'b0;
  assign debug_ad_sf_col_addr[6] = 1'b0;
  assign debug_ad_sf_col_addr[7] = 1'b0;
  assign debug_ad_sf_col_addr[8] = 1'b0;
  assign debug_ad_sf_col_addr[9] = 1'b0;
  assign debug_ad_sf_col_addr[10] = 1'b0;
  assign debug_ad_sf_col_addr[11] = 1'b0;
  assign debug_ad_sf_col_addr[12] = 1'b0;
  assign debug_ad_sf_col_addr[13] = 1'b0;
  assign debug_ad_sf_col_addr[14] = 1'b0;
  assign debug_ad_sf_col_addr[15] = 1'b0;
  assign debug_ad_sf_row_addr[0] = 1'b0;
  assign debug_ad_sf_row_addr[1] = 1'b0;
  assign debug_ad_sf_row_addr[2] = 1'b0;
  assign debug_ad_sf_row_addr[3] = 1'b0;
  assign debug_ad_sf_row_addr[4] = 1'b0;
  assign debug_ad_sf_row_addr[5] = 1'b0;
  assign debug_ad_sf_row_addr[6] = 1'b0;
  assign debug_ad_sf_row_addr[7] = 1'b0;
  assign debug_ad_sf_row_addr[8] = 1'b0;
  assign debug_ad_sf_row_addr[9] = 1'b0;
  assign debug_ad_sf_row_addr[10] = 1'b0;
  assign debug_ad_sf_row_addr[11] = 1'b0;
  assign debug_ad_sf_row_addr[12] = 1'b0;
  assign debug_ad_sf_row_addr[13] = 1'b0;
  assign debug_ad_sf_row_addr[14] = 1'b0;
  assign debug_ad_sf_row_addr[15] = 1'b0;
  assign debug_ad_sf_bank_addr[0] = 1'b0;
  assign debug_ad_sf_bank_addr[1] = 1'b0;
  assign hresp[0] = 1'b0;
  assign hresp[1] = 1'b0;

  INV_X4 U2 ( .A(n4), .ZN(n3) );
  INV_X1 U4 ( .A(big_endian), .ZN(n4) );
  DW_memctl_hiu U_hiu ( .hclk(hclk), .hresetn(hresetn), .hsel_mem(hsel_mem), 
        .hsel_reg(hsel_reg), .htrans(htrans), .hwrite(hwrite), .hsize(hsize), 
        .hburst(hburst), .hready(hready), .hready_resp(hready_resp), .hresp({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}), .haddr(haddr), 
        .hwdata(hwdata), .hrdata(hrdata), .hiu_req(hiu_req), .hiu_burst_size(
        hiu_burst_size), .hiu_wrap_burst(hiu_wrap_burst), .hiu_rw(hiu_rw), 
        .hiu_terminate(hiu_terminate), .hiu_addr({debug_hiu_addr[31:1], 
        SYNOPSYS_UNCONNECTED_3}), .hiu_data(hiu_data), .hiu_haddr(hiu_haddr), 
        .hiu_hsize(hiu_hsize), .miu_burst_done(miu_burst_done), .miu_push_n(
        miu_push_n), .miu_pop_n(miu_pop_n), .miu_data({miu_data[31:14], n2, 
        miu_data[12:0]}), .miu_data_width({1'b0, 1'b0}), .miu_col_width({1'b0, 
        1'b0, 1'b0, 1'b0}), .big_endian(n3) );
  DW_memctl_miu U_miu ( .hclk(hclk), .hclk_2x(hclk_2x), .hresetn(hresetn), 
        .scan_mode(scan_mode), .hiu_mem_req(hiu_req[1]), .hiu_reg_req(
        hiu_req[0]), .hiu_rw(hiu_rw), .hiu_burst_size(hiu_burst_size), 
        .hiu_wrapped_burst(hiu_wrap_burst), .hiu_terminate(hiu_terminate), 
        .hiu_addr({debug_hiu_addr[31:1], 1'b0}), .hiu_haddr(hiu_haddr), 
        .hiu_hsize(hiu_hsize), .hiu_wr_data(hiu_data), .s_rd_data(s_rd_data), 
        .miu_burst_done(miu_burst_done), .miu_pop_n(miu_pop_n), .miu_push_n(
        miu_push_n), .miu_col_addr_width({SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7}), .miu_data_width({SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9}), .m_addr(
        {SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25}), .s_addr(s_addr), 
        .s_bank_addr(s_bank_addr), .s_ras_n(s_ras_n), .s_cas_n(s_cas_n), 
        .s_sel_n(s_sel_n[0]), .s_cke(s_cke), .s_we_n(s_we_n), .s_wr_data(
        s_wr_data), .s_dqm(s_dqm), .s_dout_valid(s_dout_valid), .s_rd_ready(
        s_rd_ready), .s_rd_start(s_rd_start), .s_rd_pop(s_rd_pop), .s_rd_end(
        s_rd_end), .s_rd_dqs_mask(s_rd_dqs_mask), .s_cas_latency(s_cas_latency), .s_read_pipe(s_read_pipe), .sf_cas_latency({SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28}), .s_sa(s_sa), 
        .s_scl(s_scl), .s_dqs(s_dqs), .s_sda_out(s_sda_out), .s_sda_in(
        s_sda_in), .s_sda_oe_n(s_sda_oe_n), .sm_addr({SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51}), .sm_bs_n({
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55}), .sm_dout_valid({
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59}), .sm_wp_n({
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62}), .sm_rd_data({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .sm_wr_data({SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94}), .remap(1'b0), .sm_clken(1'b0), .sm_ready(
        1'b0), .sm_data_width_set0({1'b0, 1'b0, 1'b0}), .m_wr_data({
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, 
        SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, 
        SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110}), .m_dout_valid({
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112}), .s_ebi_gnt(1'b0), 
        .sm_ebi_gnt(1'b0), .power_down(power_down), .sf_power_down(1'b0), 
        .sm_power_down(1'b0), .clear_sr_dp(clear_sr_dp), .sf_clear_dp(1'b0), 
        .big_endian(n3), .miu_rd_data_out({miu_data[31:14], n2, miu_data[12:0]}), .gpi(gpi), .gpo(gpo), .debug_ad_bank_addr(debug_ad_bank_addr), 
        .debug_ad_row_addr(debug_ad_row_addr), .debug_ad_sf_bank_addr({
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114}), 
        .debug_ad_sf_row_addr({SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130}), .debug_ad_sf_col_addr({
        SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, 
        SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134, 
        SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136, 
        SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, 
        SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146}), .debug_smc_cs({
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150}), .debug_ref_req(
        debug_ref_req), .debug_ad_col_addr_15_(debug_ad_col_addr[15]), 
        .debug_ad_col_addr_14_(debug_ad_col_addr[14]), .debug_ad_col_addr_11_(
        debug_ad_col_addr[11]), .debug_ad_col_addr_10_(debug_ad_col_addr[10]), 
        .debug_ad_col_addr_9_(debug_ad_col_addr[9]), .debug_ad_col_addr_8_(
        debug_ad_col_addr[8]), .debug_ad_col_addr_7_(debug_ad_col_addr[7]), 
        .debug_ad_col_addr_6_(debug_ad_col_addr[6]), .debug_ad_col_addr_5_(
        debug_ad_col_addr[5]), .debug_ad_col_addr_4_(debug_ad_col_addr[4]), 
        .debug_ad_col_addr_3_(debug_ad_col_addr[3]), .debug_ad_col_addr_2_(
        debug_ad_col_addr[2]), .debug_ad_col_addr_1_(debug_ad_col_addr[1]), 
        .debug_ad_col_addr_0_(debug_ad_col_addr[0]), 
        .debug_ad_col_addr_13__BAR_BAR(debug_ad_col_addr[13]), 
        .debug_ad_col_addr_12__BAR_BAR(debug_ad_col_addr[12]) );
endmodule

