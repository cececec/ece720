
module cortexm0ds_logic ( hclk, hreset_n, haddr_o, hburst_o, hmastlock_o, 
        hprot_o, hsize_o, htrans_o, hwdata_o, hwrite_o, hrdata_i, hready_i, 
        hresp_i, nmi_i, irq_i, txev_o, rxev_i, lockup_o, sys_reset_req_o, 
        sleeping_o, vis_r0_o, vis_r1_o, vis_r2_o, vis_r3_o, vis_r4_o, vis_r5_o, 
        vis_r6_o, vis_r7_o, vis_r8_o, vis_r9_o, vis_r10_o, vis_r11_o, 
        vis_r12_o, vis_r14_o, vis_msp_o, vis_psp_o, vis_pc_o, vis_apsr_o, 
        vis_tbit_o, vis_ipsr_o, vis_control_o, vis_primask_o );
  output [31:0] haddr_o;
  output [2:0] hburst_o;
  output [3:0] hprot_o;
  output [2:0] hsize_o;
  output [1:0] htrans_o;
  output [31:0] hwdata_o;
  input [31:0] hrdata_i;
  input [15:0] irq_i;
  output [31:0] vis_r0_o;
  output [31:0] vis_r1_o;
  output [31:0] vis_r2_o;
  output [31:0] vis_r3_o;
  output [31:0] vis_r4_o;
  output [31:0] vis_r5_o;
  output [31:0] vis_r6_o;
  output [31:0] vis_r7_o;
  output [31:0] vis_r8_o;
  output [31:0] vis_r9_o;
  output [31:0] vis_r10_o;
  output [31:0] vis_r11_o;
  output [31:0] vis_r12_o;
  output [31:0] vis_r14_o;
  output [29:0] vis_msp_o;
  output [29:0] vis_psp_o;
  output [30:0] vis_pc_o;
  output [3:0] vis_apsr_o;
  output [5:0] vis_ipsr_o;
  input hclk, hreset_n, hready_i, hresp_i, nmi_i, rxev_i;
  output hmastlock_o, hwrite_o, txev_o, lockup_o, sys_reset_req_o, sleeping_o,
         vis_tbit_o, vis_control_o, vis_primask_o;
  wire   n8698, n8706, n9796, n9972, n10055, n10553, n11746, n11928, n11929,
         n11939, n11945, n11957, n11971, n13747, n13758, n13795, n13813,
         n13835, n13846, n13870, n13894, n13907, n13919, n13932, n13951,
         n13963, n13989, n14001, n14432, n14825, n14928, n14934, n14956,
         U811_Z_0, U810_Z_0, U809_Z_0, U806_Z_0, U805_Z_0, U804_Z_0, U803_Z_0,
         U802_Z_0, U801_Z_0, U800_Z_0, U799_Z_0, U798_Z_0, U797_Z_0, U795_Z_0,
         U792_Z_0, U791_Z_0, U790_Z_0, U789_Z_0, U788_Z_0, U787_Z_0, U786_Z_0,
         U785_Z_0, U784_Z_0, U783_Z_0, U782_Z_0, U781_Z_0, U780_Z_0, U779_Z_0,
         U778_Z_0, U777_Z_0, U776_Z_0, U775_Z_0, U774_Z_0, U773_Z_0, U772_Z_0,
         U771_Z_0, U770_Z_0, U769_Z_0, U768_Z_0, U767_Z_0, U766_Z_0, U765_Z_0,
         U764_Z_0, U763_Z_0, U762_Z_0, U761_Z_0, U760_Z_0, U756_Z_0, U755_Z_0,
         U754_Z_0, U752_Z_0, U751_Z_0, U750_Z_0, U749_Z_0, U748_Z_0, U747_Z_0,
         U746_Z_0, U745_Z_0, U744_Z_0, U743_Z_0, U742_Z_0, U741_Z_0, U740_Z_0,
         U739_Z_0, U738_Z_0, U737_Z_0, U736_Z_0, U735_Z_0, U734_Z_0, U733_Z_0,
         U732_Z_0, U731_Z_0, U730_Z_0, U729_Z_0, U728_Z_0, U727_Z_0, U726_Z_0,
         U725_Z_0, U724_Z_0, U723_Z_0, U722_Z_0, U721_Z_0, U720_Z_0, U719_Z_0,
         U718_Z_0, U717_Z_0, U716_Z_0, U715_Z_0, U714_Z_0, U713_Z_0, U712_Z_0,
         U711_Z_0, U710_Z_0, U709_Z_0, U708_Z_0, U707_Z_0, U706_Z_0, U705_Z_0,
         U704_Z_0, U703_Z_0, U702_Z_0, U701_Z_0, U700_Z_0, U699_Z_0, U698_Z_0,
         U697_Z_0, U696_Z_0, U695_Z_0, U694_Z_0, U693_Z_0, U692_Z_0, U691_Z_0,
         U687_Z_0, U686_Z_0, U685_Z_0, U684_Z_0, U683_Z_0, U682_Z_0, U681_Z_0,
         U680_Z_0, U679_Z_0, U678_Z_0, U677_Z_0, U676_Z_0, U675_Z_0, U674_Z_0,
         U673_Z_0, U672_Z_0, U671_Z_0, U670_Z_0, U669_Z_0, U668_Z_0, U667_Z_0,
         U666_Z_0, U665_Z_0, U664_Z_0, U663_Z_0, U662_Z_0, U661_Z_0, U660_Z_0,
         U659_Z_0, U658_Z_0, U657_Z_0, U656_Z_0, U655_Z_0, U654_Z_0, U653_Z_0,
         U652_Z_0, U651_Z_0, U650_Z_0, U649_Z_0, U648_Z_0, U647_Z_0, U646_Z_0,
         U645_Z_0, U644_Z_0, U643_Z_0, U642_Z_0, U641_Z_0, U640_Z_0, U639_Z_0,
         U638_Z_0, U637_Z_0, U636_Z_0, U635_Z_0, U634_Z_0, U633_Z_0, U632_Z_0,
         U631_Z_0, U630_Z_0, U629_Z_0, U628_Z_0, U627_Z_0, U626_Z_0, U625_Z_0,
         U624_Z_0, U623_Z_0, U622_Z_0, U621_Z_0, U620_Z_0, U619_Z_0, U618_Z_0,
         U617_Z_0, U614_Z_0, U613_Z_0, U612_Z_0, U611_Z_0, U610_Z_0, U609_Z_0,
         U608_Z_0, U607_Z_0, U606_Z_0, U605_Z_0, U604_Z_0, U603_Z_0, U602_Z_0,
         U601_Z_0, U600_Z_0, U599_Z_0, U598_Z_0, U597_Z_0, U596_Z_0, U595_Z_0,
         U594_Z_0, U593_Z_0, U592_Z_0, U591_Z_0, U590_Z_0, U589_Z_0, U588_Z_0,
         U587_Z_0, U586_Z_0, U585_Z_0, U584_Z_0, U583_Z_0, U582_Z_0, U581_Z_0,
         U580_Z_0, U579_Z_0, U578_Z_0, U577_Z_0, U576_Z_0, U575_Z_0, U574_Z_0,
         U573_Z_0, U572_Z_0, U571_Z_0, U570_Z_0, U569_Z_0, U568_Z_0, U567_Z_0,
         U566_Z_0, U565_Z_0, U564_Z_0, U563_Z_0, U562_Z_0, U561_Z_0, U560_Z_0,
         U559_Z_0, U558_Z_0, U557_Z_0, U556_Z_0, U555_Z_0, U554_Z_0, U553_Z_0,
         U552_Z_0, U551_Z_0, U550_Z_0, U549_Z_0, U548_Z_0, U547_Z_0, U546_Z_0,
         U545_Z_0, U544_Z_0, U543_Z_0, U542_Z_0, U541_Z_0, U540_Z_0, U539_Z_0,
         U538_Z_0, U537_Z_0, U536_Z_0, U535_Z_0, U534_Z_0, U533_Z_0, U532_Z_0,
         U531_Z_0, U530_Z_0, U529_Z_0, U528_Z_0, U527_Z_0, U526_Z_0, U525_Z_0,
         U524_Z_0, U523_Z_0, U522_Z_0, U521_Z_0, U520_Z_0, U519_Z_0, U518_Z_0,
         U517_Z_0, U516_Z_0, U515_Z_0, U514_Z_0, U513_Z_0, U512_Z_0, U511_Z_0,
         U510_Z_0, U509_Z_0, U508_Z_0, U507_Z_0, U506_Z_0, U505_Z_0, U504_Z_0,
         U503_Z_0, U502_Z_0, U501_Z_0, U500_Z_0, U499_Z_0, U498_Z_0, U497_Z_0,
         U496_Z_0, U495_Z_0, U494_Z_0, U493_Z_0, U492_Z_0, U491_Z_0, U490_Z_0,
         U489_Z_0, U488_Z_0, U487_Z_0, U486_Z_0, U483_Z_0, U482_Z_0, U481_Z_0,
         U480_Z_0, U479_Z_0, U478_Z_0, U477_Z_0, U476_Z_0, U475_Z_0, U474_Z_0,
         U473_Z_0, U472_Z_0, U471_Z_0, U470_Z_0, U469_Z_0, U468_Z_0, U467_Z_0,
         U466_Z_0, U465_Z_0, U464_Z_0, U463_Z_0, U462_Z_0, U461_Z_0, U460_Z_0,
         U459_Z_0, U458_Z_0, U457_Z_0, U456_Z_0, U455_Z_0, U454_Z_0, U453_Z_0,
         U452_Z_0, U449_Z_0, U448_Z_0, U447_Z_0, U446_Z_0, U445_Z_0, U444_Z_0,
         U443_Z_0, U442_Z_0, U441_Z_0, U440_Z_0, U439_Z_0, U438_Z_0, U437_Z_0,
         U436_Z_0, U435_Z_0, U434_Z_0, U433_Z_0, U432_Z_0, U431_Z_0, U430_Z_0,
         U429_Z_0, U428_Z_0, U427_Z_0, U426_Z_0, U425_Z_0, U424_Z_0, U423_Z_0,
         U422_Z_0, U421_Z_0, U420_Z_0, U419_Z_0, U418_Z_0, U415_Z_0, U414_Z_0,
         U413_Z_0, U412_Z_0, U411_Z_0, U410_Z_0, U409_Z_0, U408_Z_0, U407_Z_0,
         U406_Z_0, U405_Z_0, U404_Z_0, U403_Z_0, U402_Z_0, U401_Z_0, U400_Z_0,
         U399_Z_0, U398_Z_0, U397_Z_0, U396_Z_0, U395_Z_0, U394_Z_0, U393_Z_0,
         U392_Z_0, U391_Z_0, U390_Z_0, U389_Z_0, U388_Z_0, U387_Z_0, U386_Z_0,
         U385_Z_0, U384_Z_0, U383_Z_0, U382_Z_0, U381_Z_0, U380_Z_0, U379_Z_0,
         U378_Z_0, U377_Z_0, U376_Z_0, U375_Z_0, U374_Z_0, U373_Z_0, U372_Z_0,
         U371_Z_0, U370_Z_0, U369_Z_0, U368_Z_0, U367_Z_0, U366_Z_0, U365_Z_0,
         U364_Z_0, U363_Z_0, U362_Z_0, U361_Z_0, U360_Z_0, U359_Z_0, U358_Z_0,
         U357_Z_0, U356_Z_0, U355_Z_0, U354_Z_0, U353_Z_0, U352_Z_0, U349_Z_0,
         U348_Z_0, U347_Z_0, U346_Z_0, U345_Z_0, U344_Z_0, U343_Z_0, U342_Z_0,
         U341_Z_0, U340_Z_0, U339_Z_0, U338_Z_0, U337_Z_0, U336_Z_0, U335_Z_0,
         U334_Z_0, U333_Z_0, U332_Z_0, U331_Z_0, U330_Z_0, U329_Z_0, U328_Z_0,
         U327_Z_0, U326_Z_0, U325_Z_0, U324_Z_0, U323_Z_0, U322_Z_0, U321_Z_0,
         U320_Z_0, U319_Z_0, U318_Z_0, U317_Z_0, U315_Z_0, U314_Z_0, U313_Z_0,
         U312_Z_0, U311_Z_0, U310_Z_0, U309_Z_0, U308_Z_0, U307_Z_0, U306_Z_0,
         U305_Z_0, U304_Z_0, U303_Z_0, U302_Z_0, U301_Z_0, U300_Z_0, U299_Z_0,
         U298_Z_0, U297_Z_0, U296_Z_0, U295_Z_0, U294_Z_0, U293_Z_0, U292_Z_0,
         U291_Z_0, U290_Z_0, U289_Z_0, U288_Z_0, U287_Z_0, U286_Z_0, U285_Z_0,
         U284_Z_0, U283_Z_0, U282_Z_0, U281_Z_0, U280_Z_0, U279_Z_0, U278_Z_0,
         U277_Z_0, U276_Z_0, U275_Z_0, U274_Z_0, U273_Z_0, U272_Z_0, U271_Z_0,
         U270_Z_0, U269_Z_0, U268_Z_0, U265_Z_0, U264_Z_0, U263_Z_0, U262_Z_0,
         U261_Z_0, U260_Z_0, U259_Z_0, U258_Z_0, U257_Z_0, U256_Z_0, U255_Z_0,
         U254_Z_0, U253_Z_0, U252_Z_0, U251_Z_0, U250_Z_0, U247_Z_0, U246_Z_0,
         U245_Z_0, U244_Z_0, U243_Z_0, U242_Z_0, U241_Z_0, U240_Z_0, U239_Z_0,
         U238_Z_0, U237_Z_0, U236_Z_0, U235_Z_0, U234_Z_0, U233_Z_0, U232_Z_0,
         U229_Z_0, U227_Z_0, U189_Z_0, U186_Z_0, U180_Z_0, U175_Z_0, U163_Z_0,
         U158_Z_0, U144_Z_0, U134_Z_0, U122_Z_0, U121_Z_0, U105_Z_0, U98_Z_0,
         U97_Z_0, U4_DATA1_0, add_2073_SUM_1_, add_2073_SUM_7_,
         add_2073_SUM_31_, add_2073_B_1_, add_2073_A_2_, add_2073_A_3_,
         add_2073_A_4_, add_2073_A_5_, add_2073_A_6_, add_2073_A_7_,
         add_2073_A_8_, add_2073_A_9_, add_2073_A_10_, add_2073_A_11_,
         add_2073_A_12_, add_2073_A_13_, add_2073_A_14_, add_2073_A_15_,
         add_2073_A_16_, add_2073_A_17_, add_2073_A_18_, add_2073_A_19_,
         add_2073_A_20_, add_2073_A_21_, add_2073_A_22_, add_2073_A_23_,
         add_2073_A_24_, add_2073_A_25_, add_2073_A_26_, add_2073_A_27_,
         add_2073_A_28_, add_2073_A_29_, add_2073_A_30_, add_2073_A_31_,
         add_2073_A_32_, add_2082_B_1_, add_2082_B_4_, add_2082_A_1_,
         add_2082_A_2_, add_2082_A_3_, add_2082_A_4_, add_2082_A_5_,
         add_2082_A_6_, add_2082_A_7_, add_2082_A_8_, add_2082_A_9_,
         add_2082_A_10_, add_2082_A_11_, add_2082_A_12_, add_2082_A_13_,
         add_2082_A_14_, add_2082_A_15_, add_2082_A_16_, add_2082_A_17_,
         add_2082_A_18_, add_2082_A_19_, add_2082_A_20_, add_2082_A_21_,
         add_2082_A_22_, add_2082_A_23_, add_2082_A_24_, add_2082_A_25_,
         add_2082_A_26_, add_2082_A_27_, add_2082_A_28_, add_2082_A_29_,
         add_2082_A_30_, add_2082_A_31_, add_2072_SUM_1_, add_2072_SUM_2_,
         add_2072_SUM_3_, add_2072_SUM_4_, add_2072_SUM_5_, add_2072_SUM_6_,
         add_2072_SUM_7_, add_2072_SUM_8_, add_2072_SUM_9_, add_2072_SUM_10_,
         add_2072_SUM_11_, add_2072_SUM_12_, add_2072_SUM_13_,
         add_2072_SUM_14_, add_2072_SUM_15_, add_2072_SUM_16_,
         add_2072_SUM_17_, add_2072_SUM_18_, add_2072_SUM_19_,
         add_2072_SUM_20_, add_2072_SUM_21_, add_2072_SUM_22_,
         add_2072_SUM_23_, add_2072_SUM_24_, add_2072_SUM_25_,
         add_2072_SUM_26_, add_2072_SUM_27_, add_2072_SUM_28_, add_2071_SUM_1_,
         add_2071_SUM_2_, add_2071_SUM_3_, add_2071_SUM_4_, add_2071_SUM_5_,
         add_2071_SUM_6_, add_2071_SUM_7_, add_2071_SUM_8_, add_2071_SUM_9_,
         add_2071_SUM_10_, add_2071_SUM_11_, add_2071_SUM_12_,
         add_2071_SUM_13_, add_2071_SUM_14_, add_2071_SUM_15_,
         add_2071_SUM_16_, add_2071_SUM_17_, add_2071_SUM_18_,
         add_2071_SUM_19_, add_2071_SUM_20_, add_2071_SUM_21_,
         add_2071_SUM_22_, add_2071_SUM_23_, add_2071_SUM_24_,
         add_2071_SUM_25_, add_2071_SUM_26_, add_2071_SUM_27_,
         add_2071_SUM_28_, add_2071_SUM_29_, sub_2069_carry_2_,
         sub_2069_carry_3_, sub_2069_carry_4_, sub_2069_carry_5_,
         sub_2069_carry_6_, sub_2069_carry_7_, sub_2069_carry_8_,
         sub_2069_SUM_1_, sub_2069_SUM_2_, sub_2069_SUM_3_, sub_2069_SUM_4_,
         sub_2069_SUM_5_, sub_2069_SUM_6_, sub_2069_SUM_7_, sub_2069_SUM_8_,
         sub_2069_A_1_, sub_2069_A_2_, sub_2069_A_3_, sub_2069_A_4_,
         sub_2069_A_5_, sub_2069_A_6_, sub_2069_A_7_, sub_2069_A_8_,
         sub_2068_carry_2_, sub_2068_carry_3_, sub_2068_carry_4_,
         sub_2068_carry_5_, sub_2068_carry_6_, sub_2068_carry_7_,
         sub_2068_carry_8_, sub_2068_carry_9_, sub_2068_carry_10_,
         sub_2068_carry_11_, sub_2068_carry_12_, sub_2068_carry_13_,
         sub_2068_carry_14_, sub_2068_carry_15_, sub_2068_carry_16_,
         sub_2068_carry_17_, sub_2068_carry_18_, sub_2068_carry_19_,
         sub_2068_carry_20_, sub_2068_carry_21_, sub_2068_carry_22_,
         sub_2068_carry_23_, sub_2068_SUM_1_, sub_2068_SUM_2_, sub_2068_SUM_3_,
         sub_2068_SUM_4_, sub_2068_SUM_5_, sub_2068_SUM_6_, sub_2068_SUM_7_,
         sub_2068_SUM_8_, sub_2068_SUM_9_, sub_2068_SUM_10_, sub_2068_SUM_11_,
         sub_2068_SUM_12_, sub_2068_SUM_13_, sub_2068_SUM_14_,
         sub_2068_SUM_15_, sub_2068_SUM_16_, sub_2068_SUM_17_,
         sub_2068_SUM_18_, sub_2068_SUM_19_, sub_2068_SUM_20_,
         sub_2068_SUM_21_, sub_2068_SUM_22_, sub_2068_A_0_, sub_2068_A_1_,
         sub_2068_A_2_, sub_2068_A_3_, sub_2068_A_4_, sub_2068_A_5_,
         sub_2068_A_6_, sub_2068_A_7_, sub_2068_A_8_, sub_2068_A_9_,
         sub_2068_A_10_, sub_2068_A_11_, sub_2068_A_12_, sub_2068_A_13_,
         sub_2068_A_14_, sub_2068_A_15_, sub_2068_A_16_, sub_2068_A_17_,
         sub_2068_A_18_, sub_2068_A_19_, sub_2068_A_20_, sub_2068_A_21_,
         sub_2068_A_22_, sub_2068_A_23_, n2, n3, n4, n5, n6, n7, n8, n9, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n27, n28, n29, n30, n31, n33, n36, n37, n39, n40, n41, n42, n44, n45,
         n46, n48, n49, n50, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n76,
         n77, n78, n80, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n99, n100, n101, n102, n104, n105, n106,
         n108, n109, n110, n111, n113, n114, n115, n117, n118, n119, n120,
         n122, n123, n124, n126, n127, n128, n129, n131, n132, n133, n135,
         n136, n137, n138, n140, n141, n142, n144, n145, n146, n148, n149,
         n150, n152, n153, n154, n156, n157, n158, n159, n160, n161, n162,
         n164, n165, n166, n167, n168, n170, n171, n172, n173, n175, n176,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n264, n265, n266,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n314, n315, n316, n317, n318, n320, n322, n324, n325, n326, n327,
         n329, n330, n333, n334, n335, n336, n337, n338, n339, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n440, n442, n443,
         n444, n445, n446, n447, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n471, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n510, n511, n512, n514,
         n515, n516, n517, n518, n519, n520, n522, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n563, n564, n565, n566, n567, n568, n569, n570, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n788, n790, n791, n792, n793, n794, n795, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n863, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1625,
         n1626, n1627, n1628, n1629, n1630, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1750, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2172, n2173, n2174,
         n2175, n2176, n2181, n2182, n2183, n2184, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2209, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2271, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2297, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2402, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2433, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2452, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2481, n2484, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2507, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2531, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2562,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2585, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2612, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2639, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2705, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2738,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2764, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2787, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2809, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2833, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2856, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2881, n2882, n2883, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2961, n2964, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3022, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3041, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3134,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3155, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3199, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3233, n3234, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3592, n3593, n3597, n3598, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3634, n3645,
         n3646, n3647, n3650, n3655, n3656, n3657, n3660, n3665, n3666, n3667,
         n3670, n3675, n3676, n3677, n3678, n3681, n3686, n3687, n3688, n3691,
         n3696, n3697, n3698, n3701, n3706, n3707, n3708, n3711, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3883, n3888, n3889, n3890, n3893, n3898, n3899, n3900,
         n3903, n3908, n3909, n3910, n3913, n3918, n3919, n3920, n3921, n3924,
         n3929, n3930, n3931, n3934, n3939, n3940, n3941, n3944, n3949, n3950,
         n3951, n3954, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3977, n3982,
         n3983, n3984, n3987, n3992, n3993, n3994, n3997, n4002, n4003, n4004,
         n4007, n4012, n4013, n4014, n4015, n4018, n4023, n4024, n4025, n4028,
         n4033, n4034, n4035, n4038, n4043, n4044, n4045, n4046, n4049, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4084, n4089, n4090,
         n4091, n4094, n4099, n4100, n4101, n4104, n4109, n4110, n4111, n4114,
         n4119, n4120, n4121, n4122, n4125, n4130, n4131, n4132, n4133, n4134,
         n4137, n4142, n4143, n4144, n4145, n4148, n4153, n4154, n4155, n4156,
         n4157, n4158, n4161, n4162, n4163, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4210, n4211, n4216, n4221, n4224,
         n4227, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4410, n4411, n4412, n4413, n4414, n4420, n4421,
         n4422, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4466, n4467,
         n4468, n4469, n4472, n4474, n4475, n4476, n4479, n4480, n4481, n4482,
         n4484, n4486, n4487, n4488, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4755, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4804, n4806, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4819, n4820, n4821, n4822, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4843, n4845,
         n4846, n4847, n4848, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5165, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5243, n5244, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17212;
  wire   [33:3] add_2082_carry;
  wire   [29:2] add_2072_carry;
  wire   [30:2] add_2071_carry;

  XNOR2_X2 sub_2068_U1_A_1 ( .A(sub_2068_A_1_), .B(sub_2068_A_0_), .ZN(
        sub_2068_SUM_1_) );
  OR2_X1 sub_2068_U1_B_1 ( .A1(sub_2068_A_1_), .A2(sub_2068_A_0_), .ZN(
        sub_2068_carry_2_) );
  XNOR2_X2 sub_2068_U1_A_2 ( .A(sub_2068_A_2_), .B(sub_2068_carry_2_), .ZN(
        sub_2068_SUM_2_) );
  OR2_X1 sub_2068_U1_B_2 ( .A1(sub_2068_A_2_), .A2(sub_2068_carry_2_), .ZN(
        sub_2068_carry_3_) );
  XNOR2_X2 sub_2068_U1_A_3 ( .A(sub_2068_A_3_), .B(sub_2068_carry_3_), .ZN(
        sub_2068_SUM_3_) );
  OR2_X1 sub_2068_U1_B_3 ( .A1(sub_2068_A_3_), .A2(sub_2068_carry_3_), .ZN(
        sub_2068_carry_4_) );
  XNOR2_X2 sub_2068_U1_A_4 ( .A(sub_2068_A_4_), .B(sub_2068_carry_4_), .ZN(
        sub_2068_SUM_4_) );
  OR2_X1 sub_2068_U1_B_4 ( .A1(sub_2068_A_4_), .A2(sub_2068_carry_4_), .ZN(
        sub_2068_carry_5_) );
  XNOR2_X2 sub_2068_U1_A_5 ( .A(sub_2068_A_5_), .B(sub_2068_carry_5_), .ZN(
        sub_2068_SUM_5_) );
  OR2_X1 sub_2068_U1_B_5 ( .A1(sub_2068_A_5_), .A2(sub_2068_carry_5_), .ZN(
        sub_2068_carry_6_) );
  XNOR2_X2 sub_2068_U1_A_6 ( .A(sub_2068_A_6_), .B(sub_2068_carry_6_), .ZN(
        sub_2068_SUM_6_) );
  OR2_X1 sub_2068_U1_B_6 ( .A1(sub_2068_A_6_), .A2(sub_2068_carry_6_), .ZN(
        sub_2068_carry_7_) );
  XNOR2_X2 sub_2068_U1_A_7 ( .A(sub_2068_A_7_), .B(sub_2068_carry_7_), .ZN(
        sub_2068_SUM_7_) );
  OR2_X1 sub_2068_U1_B_7 ( .A1(sub_2068_A_7_), .A2(sub_2068_carry_7_), .ZN(
        sub_2068_carry_8_) );
  XNOR2_X2 sub_2068_U1_A_8 ( .A(sub_2068_A_8_), .B(sub_2068_carry_8_), .ZN(
        sub_2068_SUM_8_) );
  OR2_X1 sub_2068_U1_B_8 ( .A1(sub_2068_A_8_), .A2(sub_2068_carry_8_), .ZN(
        sub_2068_carry_9_) );
  XNOR2_X2 sub_2068_U1_A_9 ( .A(sub_2068_A_9_), .B(sub_2068_carry_9_), .ZN(
        sub_2068_SUM_9_) );
  OR2_X1 sub_2068_U1_B_9 ( .A1(sub_2068_A_9_), .A2(sub_2068_carry_9_), .ZN(
        sub_2068_carry_10_) );
  XNOR2_X2 sub_2068_U1_A_10 ( .A(sub_2068_A_10_), .B(sub_2068_carry_10_), .ZN(
        sub_2068_SUM_10_) );
  OR2_X1 sub_2068_U1_B_10 ( .A1(sub_2068_A_10_), .A2(sub_2068_carry_10_), .ZN(
        sub_2068_carry_11_) );
  XNOR2_X2 sub_2068_U1_A_11 ( .A(sub_2068_A_11_), .B(sub_2068_carry_11_), .ZN(
        sub_2068_SUM_11_) );
  OR2_X1 sub_2068_U1_B_11 ( .A1(sub_2068_A_11_), .A2(sub_2068_carry_11_), .ZN(
        sub_2068_carry_12_) );
  XNOR2_X2 sub_2068_U1_A_12 ( .A(sub_2068_A_12_), .B(sub_2068_carry_12_), .ZN(
        sub_2068_SUM_12_) );
  OR2_X1 sub_2068_U1_B_12 ( .A1(sub_2068_A_12_), .A2(sub_2068_carry_12_), .ZN(
        sub_2068_carry_13_) );
  XNOR2_X2 sub_2068_U1_A_13 ( .A(sub_2068_A_13_), .B(sub_2068_carry_13_), .ZN(
        sub_2068_SUM_13_) );
  OR2_X1 sub_2068_U1_B_13 ( .A1(sub_2068_A_13_), .A2(sub_2068_carry_13_), .ZN(
        sub_2068_carry_14_) );
  XNOR2_X2 sub_2068_U1_A_14 ( .A(sub_2068_A_14_), .B(sub_2068_carry_14_), .ZN(
        sub_2068_SUM_14_) );
  OR2_X1 sub_2068_U1_B_14 ( .A1(sub_2068_A_14_), .A2(sub_2068_carry_14_), .ZN(
        sub_2068_carry_15_) );
  XNOR2_X2 sub_2068_U1_A_15 ( .A(sub_2068_A_15_), .B(sub_2068_carry_15_), .ZN(
        sub_2068_SUM_15_) );
  OR2_X1 sub_2068_U1_B_15 ( .A1(sub_2068_A_15_), .A2(sub_2068_carry_15_), .ZN(
        sub_2068_carry_16_) );
  XNOR2_X2 sub_2068_U1_A_16 ( .A(sub_2068_A_16_), .B(sub_2068_carry_16_), .ZN(
        sub_2068_SUM_16_) );
  OR2_X1 sub_2068_U1_B_16 ( .A1(sub_2068_A_16_), .A2(sub_2068_carry_16_), .ZN(
        sub_2068_carry_17_) );
  XNOR2_X2 sub_2068_U1_A_17 ( .A(sub_2068_A_17_), .B(sub_2068_carry_17_), .ZN(
        sub_2068_SUM_17_) );
  OR2_X1 sub_2068_U1_B_17 ( .A1(sub_2068_A_17_), .A2(sub_2068_carry_17_), .ZN(
        sub_2068_carry_18_) );
  XNOR2_X2 sub_2068_U1_A_18 ( .A(sub_2068_A_18_), .B(sub_2068_carry_18_), .ZN(
        sub_2068_SUM_18_) );
  OR2_X1 sub_2068_U1_B_18 ( .A1(sub_2068_A_18_), .A2(sub_2068_carry_18_), .ZN(
        sub_2068_carry_19_) );
  XNOR2_X2 sub_2068_U1_A_19 ( .A(sub_2068_A_19_), .B(sub_2068_carry_19_), .ZN(
        sub_2068_SUM_19_) );
  OR2_X1 sub_2068_U1_B_19 ( .A1(sub_2068_A_19_), .A2(sub_2068_carry_19_), .ZN(
        sub_2068_carry_20_) );
  XNOR2_X2 sub_2068_U1_A_20 ( .A(sub_2068_A_20_), .B(sub_2068_carry_20_), .ZN(
        sub_2068_SUM_20_) );
  OR2_X1 sub_2068_U1_B_20 ( .A1(sub_2068_A_20_), .A2(sub_2068_carry_20_), .ZN(
        sub_2068_carry_21_) );
  XNOR2_X2 sub_2068_U1_A_21 ( .A(sub_2068_A_21_), .B(sub_2068_carry_21_), .ZN(
        sub_2068_SUM_21_) );
  OR2_X1 sub_2068_U1_B_21 ( .A1(sub_2068_A_21_), .A2(sub_2068_carry_21_), .ZN(
        sub_2068_carry_22_) );
  XNOR2_X2 sub_2068_U1_A_22 ( .A(sub_2068_A_22_), .B(sub_2068_carry_22_), .ZN(
        sub_2068_SUM_22_) );
  OR2_X1 sub_2068_U1_B_22 ( .A1(sub_2068_A_22_), .A2(sub_2068_carry_22_), .ZN(
        sub_2068_carry_23_) );
  XNOR2_X2 sub_2069_U1_A_1 ( .A(sub_2069_A_1_), .B(n5829), .ZN(sub_2069_SUM_1_) );
  OR2_X1 sub_2069_U1_B_1 ( .A1(sub_2069_A_1_), .A2(n5829), .ZN(
        sub_2069_carry_2_) );
  XNOR2_X2 sub_2069_U1_A_2 ( .A(sub_2069_A_2_), .B(sub_2069_carry_2_), .ZN(
        sub_2069_SUM_2_) );
  OR2_X1 sub_2069_U1_B_2 ( .A1(sub_2069_A_2_), .A2(sub_2069_carry_2_), .ZN(
        sub_2069_carry_3_) );
  XNOR2_X2 sub_2069_U1_A_3 ( .A(sub_2069_A_3_), .B(sub_2069_carry_3_), .ZN(
        sub_2069_SUM_3_) );
  OR2_X1 sub_2069_U1_B_3 ( .A1(sub_2069_A_3_), .A2(sub_2069_carry_3_), .ZN(
        sub_2069_carry_4_) );
  XNOR2_X2 sub_2069_U1_A_4 ( .A(sub_2069_A_4_), .B(sub_2069_carry_4_), .ZN(
        sub_2069_SUM_4_) );
  OR2_X1 sub_2069_U1_B_4 ( .A1(sub_2069_A_4_), .A2(sub_2069_carry_4_), .ZN(
        sub_2069_carry_5_) );
  XNOR2_X2 sub_2069_U1_A_5 ( .A(sub_2069_A_5_), .B(sub_2069_carry_5_), .ZN(
        sub_2069_SUM_5_) );
  OR2_X1 sub_2069_U1_B_5 ( .A1(sub_2069_A_5_), .A2(sub_2069_carry_5_), .ZN(
        sub_2069_carry_6_) );
  XNOR2_X2 sub_2069_U1_A_6 ( .A(sub_2069_A_6_), .B(sub_2069_carry_6_), .ZN(
        sub_2069_SUM_6_) );
  OR2_X1 sub_2069_U1_B_6 ( .A1(sub_2069_A_6_), .A2(sub_2069_carry_6_), .ZN(
        sub_2069_carry_7_) );
  XNOR2_X2 sub_2069_U1_A_7 ( .A(sub_2069_A_7_), .B(sub_2069_carry_7_), .ZN(
        sub_2069_SUM_7_) );
  OR2_X1 sub_2069_U1_B_7 ( .A1(sub_2069_A_7_), .A2(sub_2069_carry_7_), .ZN(
        sub_2069_carry_8_) );
  XNOR2_X2 sub_2069_U1_A_8 ( .A(sub_2069_A_8_), .B(sub_2069_carry_8_), .ZN(
        sub_2069_SUM_8_) );
  HA_X1 add_2071_U1_1_1 ( .A(vis_pc_o[1]), .B(vis_pc_o[0]), .CO(
        add_2071_carry[2]), .S(add_2071_SUM_1_) );
  HA_X1 add_2071_U1_1_2 ( .A(vis_pc_o[2]), .B(add_2071_carry[2]), .CO(
        add_2071_carry[3]), .S(add_2071_SUM_2_) );
  HA_X1 add_2071_U1_1_3 ( .A(vis_pc_o[3]), .B(add_2071_carry[3]), .CO(
        add_2071_carry[4]), .S(add_2071_SUM_3_) );
  HA_X1 add_2071_U1_1_4 ( .A(vis_pc_o[4]), .B(add_2071_carry[4]), .CO(
        add_2071_carry[5]), .S(add_2071_SUM_4_) );
  HA_X1 add_2071_U1_1_5 ( .A(vis_pc_o[5]), .B(add_2071_carry[5]), .CO(
        add_2071_carry[6]), .S(add_2071_SUM_5_) );
  HA_X1 add_2071_U1_1_6 ( .A(vis_pc_o[6]), .B(add_2071_carry[6]), .CO(
        add_2071_carry[7]), .S(add_2071_SUM_6_) );
  HA_X1 add_2071_U1_1_7 ( .A(vis_pc_o[7]), .B(add_2071_carry[7]), .CO(
        add_2071_carry[8]), .S(add_2071_SUM_7_) );
  HA_X1 add_2071_U1_1_8 ( .A(vis_pc_o[8]), .B(add_2071_carry[8]), .CO(
        add_2071_carry[9]), .S(add_2071_SUM_8_) );
  HA_X1 add_2071_U1_1_9 ( .A(vis_pc_o[9]), .B(add_2071_carry[9]), .CO(
        add_2071_carry[10]), .S(add_2071_SUM_9_) );
  HA_X1 add_2071_U1_1_10 ( .A(vis_pc_o[10]), .B(add_2071_carry[10]), .CO(
        add_2071_carry[11]), .S(add_2071_SUM_10_) );
  HA_X1 add_2071_U1_1_11 ( .A(vis_pc_o[11]), .B(add_2071_carry[11]), .CO(
        add_2071_carry[12]), .S(add_2071_SUM_11_) );
  HA_X1 add_2071_U1_1_12 ( .A(vis_pc_o[12]), .B(add_2071_carry[12]), .CO(
        add_2071_carry[13]), .S(add_2071_SUM_12_) );
  HA_X1 add_2071_U1_1_13 ( .A(vis_pc_o[13]), .B(add_2071_carry[13]), .CO(
        add_2071_carry[14]), .S(add_2071_SUM_13_) );
  HA_X1 add_2071_U1_1_14 ( .A(vis_pc_o[14]), .B(add_2071_carry[14]), .CO(
        add_2071_carry[15]), .S(add_2071_SUM_14_) );
  HA_X1 add_2071_U1_1_15 ( .A(vis_pc_o[15]), .B(add_2071_carry[15]), .CO(
        add_2071_carry[16]), .S(add_2071_SUM_15_) );
  HA_X1 add_2071_U1_1_16 ( .A(vis_pc_o[16]), .B(add_2071_carry[16]), .CO(
        add_2071_carry[17]), .S(add_2071_SUM_16_) );
  HA_X1 add_2071_U1_1_17 ( .A(vis_pc_o[17]), .B(add_2071_carry[17]), .CO(
        add_2071_carry[18]), .S(add_2071_SUM_17_) );
  HA_X1 add_2071_U1_1_18 ( .A(vis_pc_o[18]), .B(add_2071_carry[18]), .CO(
        add_2071_carry[19]), .S(add_2071_SUM_18_) );
  HA_X1 add_2071_U1_1_19 ( .A(vis_pc_o[19]), .B(add_2071_carry[19]), .CO(
        add_2071_carry[20]), .S(add_2071_SUM_19_) );
  HA_X1 add_2071_U1_1_20 ( .A(vis_pc_o[20]), .B(add_2071_carry[20]), .CO(
        add_2071_carry[21]), .S(add_2071_SUM_20_) );
  HA_X1 add_2071_U1_1_21 ( .A(vis_pc_o[21]), .B(add_2071_carry[21]), .CO(
        add_2071_carry[22]), .S(add_2071_SUM_21_) );
  HA_X1 add_2071_U1_1_22 ( .A(vis_pc_o[22]), .B(add_2071_carry[22]), .CO(
        add_2071_carry[23]), .S(add_2071_SUM_22_) );
  HA_X1 add_2071_U1_1_23 ( .A(vis_pc_o[23]), .B(add_2071_carry[23]), .CO(
        add_2071_carry[24]), .S(add_2071_SUM_23_) );
  HA_X1 add_2071_U1_1_24 ( .A(vis_pc_o[24]), .B(add_2071_carry[24]), .CO(
        add_2071_carry[25]), .S(add_2071_SUM_24_) );
  HA_X1 add_2071_U1_1_25 ( .A(vis_pc_o[25]), .B(add_2071_carry[25]), .CO(
        add_2071_carry[26]), .S(add_2071_SUM_25_) );
  HA_X1 add_2071_U1_1_26 ( .A(vis_pc_o[26]), .B(add_2071_carry[26]), .CO(
        add_2071_carry[27]), .S(add_2071_SUM_26_) );
  HA_X1 add_2071_U1_1_27 ( .A(vis_pc_o[27]), .B(add_2071_carry[27]), .CO(
        add_2071_carry[28]), .S(add_2071_SUM_27_) );
  HA_X1 add_2071_U1_1_28 ( .A(vis_pc_o[28]), .B(add_2071_carry[28]), .CO(
        add_2071_carry[29]), .S(add_2071_SUM_28_) );
  HA_X1 add_2071_U1_1_29 ( .A(vis_pc_o[29]), .B(add_2071_carry[29]), .CO(
        add_2071_carry[30]), .S(add_2071_SUM_29_) );
  HA_X1 add_2072_U1_1_1 ( .A(vis_pc_o[2]), .B(n5797), .CO(add_2072_carry[2]), 
        .S(add_2072_SUM_1_) );
  HA_X1 add_2072_U1_1_2 ( .A(vis_pc_o[3]), .B(add_2072_carry[2]), .CO(
        add_2072_carry[3]), .S(add_2072_SUM_2_) );
  HA_X1 add_2072_U1_1_3 ( .A(vis_pc_o[4]), .B(add_2072_carry[3]), .CO(
        add_2072_carry[4]), .S(add_2072_SUM_3_) );
  HA_X1 add_2072_U1_1_4 ( .A(vis_pc_o[5]), .B(add_2072_carry[4]), .CO(
        add_2072_carry[5]), .S(add_2072_SUM_4_) );
  HA_X1 add_2072_U1_1_5 ( .A(vis_pc_o[6]), .B(add_2072_carry[5]), .CO(
        add_2072_carry[6]), .S(add_2072_SUM_5_) );
  HA_X1 add_2072_U1_1_6 ( .A(vis_pc_o[7]), .B(add_2072_carry[6]), .CO(
        add_2072_carry[7]), .S(add_2072_SUM_6_) );
  HA_X1 add_2072_U1_1_7 ( .A(vis_pc_o[8]), .B(add_2072_carry[7]), .CO(
        add_2072_carry[8]), .S(add_2072_SUM_7_) );
  HA_X1 add_2072_U1_1_8 ( .A(vis_pc_o[9]), .B(add_2072_carry[8]), .CO(
        add_2072_carry[9]), .S(add_2072_SUM_8_) );
  HA_X1 add_2072_U1_1_9 ( .A(vis_pc_o[10]), .B(add_2072_carry[9]), .CO(
        add_2072_carry[10]), .S(add_2072_SUM_9_) );
  HA_X1 add_2072_U1_1_10 ( .A(vis_pc_o[11]), .B(add_2072_carry[10]), .CO(
        add_2072_carry[11]), .S(add_2072_SUM_10_) );
  HA_X1 add_2072_U1_1_11 ( .A(vis_pc_o[12]), .B(add_2072_carry[11]), .CO(
        add_2072_carry[12]), .S(add_2072_SUM_11_) );
  HA_X1 add_2072_U1_1_12 ( .A(vis_pc_o[13]), .B(add_2072_carry[12]), .CO(
        add_2072_carry[13]), .S(add_2072_SUM_12_) );
  HA_X1 add_2072_U1_1_13 ( .A(vis_pc_o[14]), .B(add_2072_carry[13]), .CO(
        add_2072_carry[14]), .S(add_2072_SUM_13_) );
  HA_X1 add_2072_U1_1_14 ( .A(vis_pc_o[15]), .B(add_2072_carry[14]), .CO(
        add_2072_carry[15]), .S(add_2072_SUM_14_) );
  HA_X1 add_2072_U1_1_15 ( .A(vis_pc_o[16]), .B(add_2072_carry[15]), .CO(
        add_2072_carry[16]), .S(add_2072_SUM_15_) );
  HA_X1 add_2072_U1_1_16 ( .A(vis_pc_o[17]), .B(add_2072_carry[16]), .CO(
        add_2072_carry[17]), .S(add_2072_SUM_16_) );
  HA_X1 add_2072_U1_1_17 ( .A(vis_pc_o[18]), .B(add_2072_carry[17]), .CO(
        add_2072_carry[18]), .S(add_2072_SUM_17_) );
  HA_X1 add_2072_U1_1_18 ( .A(vis_pc_o[19]), .B(add_2072_carry[18]), .CO(
        add_2072_carry[19]), .S(add_2072_SUM_18_) );
  HA_X1 add_2072_U1_1_19 ( .A(vis_pc_o[20]), .B(add_2072_carry[19]), .CO(
        add_2072_carry[20]), .S(add_2072_SUM_19_) );
  HA_X1 add_2072_U1_1_20 ( .A(vis_pc_o[21]), .B(add_2072_carry[20]), .CO(
        add_2072_carry[21]), .S(add_2072_SUM_20_) );
  HA_X1 add_2072_U1_1_21 ( .A(vis_pc_o[22]), .B(add_2072_carry[21]), .CO(
        add_2072_carry[22]), .S(add_2072_SUM_21_) );
  HA_X1 add_2072_U1_1_22 ( .A(vis_pc_o[23]), .B(add_2072_carry[22]), .CO(
        add_2072_carry[23]), .S(add_2072_SUM_22_) );
  HA_X1 add_2072_U1_1_23 ( .A(vis_pc_o[24]), .B(add_2072_carry[23]), .CO(
        add_2072_carry[24]), .S(add_2072_SUM_23_) );
  HA_X1 add_2072_U1_1_24 ( .A(vis_pc_o[25]), .B(add_2072_carry[24]), .CO(
        add_2072_carry[25]), .S(add_2072_SUM_24_) );
  HA_X1 add_2072_U1_1_25 ( .A(vis_pc_o[26]), .B(add_2072_carry[25]), .CO(
        add_2072_carry[26]), .S(add_2072_SUM_25_) );
  HA_X1 add_2072_U1_1_26 ( .A(vis_pc_o[27]), .B(add_2072_carry[26]), .CO(
        add_2072_carry[27]), .S(add_2072_SUM_26_) );
  HA_X1 add_2072_U1_1_27 ( .A(vis_pc_o[28]), .B(add_2072_carry[27]), .CO(
        add_2072_carry[28]), .S(add_2072_SUM_27_) );
  HA_X1 add_2072_U1_1_28 ( .A(vis_pc_o[29]), .B(add_2072_carry[28]), .CO(
        add_2072_carry[29]), .S(add_2072_SUM_28_) );
  FA_X1 add_2082_U1_2 ( .A(add_2082_A_2_), .B(n5822), .CI(n16691), .CO(
        add_2082_carry[3]), .S(add_2073_A_2_) );
  FA_X1 add_2082_U1_3 ( .A(add_2082_A_3_), .B(n5806), .CI(add_2082_carry[3]), 
        .CO(add_2082_carry[4]), .S(add_2073_A_3_) );
  FA_X1 add_2082_U1_4 ( .A(add_2082_A_4_), .B(add_2082_B_4_), .CI(
        add_2082_carry[4]), .CO(add_2082_carry[5]), .S(add_2073_A_4_) );
  FA_X1 add_2082_U1_5 ( .A(add_2082_A_5_), .B(n5801), .CI(add_2082_carry[5]), 
        .CO(add_2082_carry[6]), .S(add_2073_A_5_) );
  FA_X1 add_2082_U1_6 ( .A(add_2082_A_6_), .B(n5802), .CI(add_2082_carry[6]), 
        .CO(add_2082_carry[7]), .S(add_2073_A_6_) );
  FA_X1 add_2082_U1_7 ( .A(add_2082_A_7_), .B(n5817), .CI(add_2082_carry[7]), 
        .CO(add_2082_carry[8]), .S(add_2073_A_7_) );
  FA_X1 add_2082_U1_8 ( .A(add_2082_A_8_), .B(n5821), .CI(add_2082_carry[8]), 
        .CO(add_2082_carry[9]), .S(add_2073_A_8_) );
  FA_X1 add_2082_U1_9 ( .A(add_2082_A_9_), .B(n5819), .CI(add_2082_carry[9]), 
        .CO(add_2082_carry[10]), .S(add_2073_A_9_) );
  FA_X1 add_2082_U1_10 ( .A(add_2082_A_10_), .B(n5805), .CI(add_2082_carry[10]), .CO(add_2082_carry[11]), .S(add_2073_A_10_) );
  FA_X1 add_2082_U1_11 ( .A(add_2082_A_11_), .B(n5804), .CI(add_2082_carry[11]), .CO(add_2082_carry[12]), .S(add_2073_A_11_) );
  FA_X1 add_2082_U1_12 ( .A(add_2082_A_12_), .B(n5820), .CI(add_2082_carry[12]), .CO(add_2082_carry[13]), .S(add_2073_A_12_) );
  FA_X1 add_2082_U1_13 ( .A(add_2082_A_13_), .B(n5807), .CI(add_2082_carry[13]), .CO(add_2082_carry[14]), .S(add_2073_A_13_) );
  FA_X1 add_2082_U1_14 ( .A(add_2082_A_14_), .B(n5808), .CI(add_2082_carry[14]), .CO(add_2082_carry[15]), .S(add_2073_A_14_) );
  FA_X1 add_2082_U1_15 ( .A(add_2082_A_15_), .B(n5809), .CI(add_2082_carry[15]), .CO(add_2082_carry[16]), .S(add_2073_A_15_) );
  FA_X1 add_2082_U1_16 ( .A(add_2082_A_16_), .B(n5818), .CI(add_2082_carry[16]), .CO(add_2082_carry[17]), .S(add_2073_A_16_) );
  FA_X1 add_2082_U1_17 ( .A(add_2082_A_17_), .B(n5810), .CI(add_2082_carry[17]), .CO(add_2082_carry[18]), .S(add_2073_A_17_) );
  FA_X1 add_2082_U1_18 ( .A(add_2082_A_18_), .B(n5811), .CI(add_2082_carry[18]), .CO(add_2082_carry[19]), .S(add_2073_A_18_) );
  FA_X1 add_2082_U1_19 ( .A(add_2082_A_19_), .B(n5812), .CI(add_2082_carry[19]), .CO(add_2082_carry[20]), .S(add_2073_A_19_) );
  FA_X1 add_2082_U1_20 ( .A(add_2082_A_20_), .B(n5813), .CI(add_2082_carry[20]), .CO(add_2082_carry[21]), .S(add_2073_A_20_) );
  FA_X1 add_2082_U1_21 ( .A(add_2082_A_21_), .B(n5814), .CI(add_2082_carry[21]), .CO(add_2082_carry[22]), .S(add_2073_A_21_) );
  FA_X1 add_2082_U1_22 ( .A(add_2082_A_22_), .B(n5815), .CI(add_2082_carry[22]), .CO(add_2082_carry[23]), .S(add_2073_A_22_) );
  FA_X1 add_2082_U1_23 ( .A(add_2082_A_23_), .B(n5816), .CI(add_2082_carry[23]), .CO(add_2082_carry[24]), .S(add_2073_A_23_) );
  FA_X1 add_2082_U1_24 ( .A(add_2082_A_24_), .B(n5803), .CI(add_2082_carry[24]), .CO(add_2082_carry[25]), .S(add_2073_A_24_) );
  FA_X1 add_2082_U1_25 ( .A(add_2082_A_25_), .B(U163_Z_0), .CI(
        add_2082_carry[25]), .CO(add_2082_carry[26]), .S(add_2073_A_25_) );
  FA_X1 add_2082_U1_26 ( .A(add_2082_A_26_), .B(n4951), .CI(add_2082_carry[26]), .CO(add_2082_carry[27]), .S(add_2073_A_26_) );
  FA_X1 add_2082_U1_27 ( .A(add_2082_A_27_), .B(n4952), .CI(add_2082_carry[27]), .CO(add_2082_carry[28]), .S(add_2073_A_27_) );
  FA_X1 add_2082_U1_28 ( .A(add_2082_A_28_), .B(U175_Z_0), .CI(
        add_2082_carry[28]), .CO(add_2082_carry[29]), .S(add_2073_A_28_) );
  FA_X1 add_2082_U1_29 ( .A(add_2082_A_29_), .B(U189_Z_0), .CI(
        add_2082_carry[29]), .CO(add_2082_carry[30]), .S(add_2073_A_29_) );
  FA_X1 add_2082_U1_30 ( .A(add_2082_A_30_), .B(U158_Z_0), .CI(
        add_2082_carry[30]), .CO(add_2082_carry[31]), .S(add_2073_A_30_) );
  FA_X1 add_2082_U1_31 ( .A(add_2082_A_31_), .B(U180_Z_0), .CI(
        add_2082_carry[31]), .CO(add_2082_carry[32]), .S(add_2073_A_31_) );
  FA_X1 add_2082_U1_32 ( .A(n4949), .B(U186_Z_0), .CI(add_2082_carry[32]), 
        .CO(add_2082_carry[33]), .S(add_2073_A_32_) );
  NOR2_X1 U3 ( .A1(n5034), .A2(n2), .ZN(sub_2069_A_8_) );
  NOR2_X1 U4 ( .A1(n5034), .A2(n3), .ZN(sub_2069_A_7_) );
  NOR2_X1 U5 ( .A1(n5034), .A2(n4), .ZN(sub_2069_A_6_) );
  NOR2_X1 U6 ( .A1(n5034), .A2(n5), .ZN(sub_2069_A_5_) );
  NOR2_X1 U8 ( .A1(n5034), .A2(n6), .ZN(sub_2069_A_4_) );
  NOR2_X1 U9 ( .A1(n5034), .A2(n7), .ZN(sub_2069_A_3_) );
  NOR2_X1 U10 ( .A1(n5034), .A2(n8), .ZN(sub_2069_A_2_) );
  NOR2_X1 U11 ( .A1(n5034), .A2(n9), .ZN(sub_2069_A_1_) );
  OAI21_X1 U13 ( .B1(n11), .B2(n12), .A(n4746), .ZN(n5654) );
  NAND4_X1 U14 ( .A1(n13), .A2(n14), .A3(hwdata_o[2]), .A4(n15), .ZN(n12) );
  NOR4_X1 U15 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n15) );
  INV_X1 U16 ( .A(n20), .ZN(n16) );
  NAND4_X1 U17 ( .A1(n21), .A2(hwdata_o[17]), .A3(n22), .A4(n23), .ZN(n11) );
  NOR4_X1 U18 ( .A1(hwdata_o[29]), .A2(hwdata_o[30]), .A3(n24), .A4(n25), .ZN(
        n23) );
  OAI221_X1 U19 ( .B1(n16644), .B2(n27), .C1(n28), .C2(n29), .A(n30), .ZN(
        n5655) );
  AOI221_X1 U20 ( .B1(n31), .B2(vis_pc_o[30]), .C1(n33), .C2(n5006), .A(n17120), .ZN(n30) );
  AND2_X1 U21 ( .A1(n17117), .A2(add_2071_carry[30]), .ZN(n33) );
  OAI21_X1 U22 ( .B1(add_2071_carry[30]), .B2(n36), .A(n37), .ZN(n31) );
  OAI211_X1 U24 ( .C1(n39), .C2(n29), .A(n40), .B(n41), .ZN(n5656) );
  AOI22_X1 U25 ( .A1(add_2071_SUM_6_), .A2(n17117), .B1(n17112), .B2(
        vis_pc_o[6]), .ZN(n41) );
  AOI21_X1 U27 ( .B1(n16726), .B2(n17116), .A(n17120), .ZN(n40) );
  OAI211_X1 U28 ( .C1(n44), .C2(n29), .A(n45), .B(n46), .ZN(n5657) );
  AOI22_X1 U29 ( .A1(add_2071_SUM_22_), .A2(n17117), .B1(n17111), .B2(
        vis_pc_o[22]), .ZN(n46) );
  AOI21_X1 U31 ( .B1(n16705), .B2(n17114), .A(n17120), .ZN(n45) );
  OAI211_X1 U32 ( .C1(n48), .C2(n29), .A(n49), .B(n50), .ZN(n5658) );
  AOI22_X1 U33 ( .A1(add_2071_SUM_14_), .A2(n17118), .B1(n17111), .B2(
        vis_pc_o[14]), .ZN(n50) );
  AOI21_X1 U34 ( .B1(n16715), .B2(n17114), .A(n17120), .ZN(n49) );
  OAI211_X1 U35 ( .C1(n5601), .C2(n37), .A(n52), .B(n53), .ZN(n5659) );
  AOI222_X1 U36 ( .A1(add_2071_SUM_19_), .A2(n17117), .B1(n16706), .B2(n17114), 
        .C1(n54), .C2(n55), .ZN(n53) );
  OAI211_X1 U37 ( .C1(n5573), .C2(n37), .A(n52), .B(n56), .ZN(n5660) );
  AOI222_X1 U38 ( .A1(add_2071_SUM_20_), .A2(n17117), .B1(n16668), .B2(n17114), 
        .C1(n54), .C2(n57), .ZN(n56) );
  INV_X1 U39 ( .A(n58), .ZN(n57) );
  OAI211_X1 U40 ( .C1(n5238), .C2(n37), .A(n52), .B(n59), .ZN(n5661) );
  AOI222_X1 U41 ( .A1(add_2071_SUM_21_), .A2(n17117), .B1(n16702), .B2(n17114), 
        .C1(n54), .C2(n60), .ZN(n59) );
  INV_X1 U42 ( .A(n61), .ZN(n60) );
  OAI211_X1 U43 ( .C1(n5237), .C2(n37), .A(n52), .B(n62), .ZN(n5662) );
  AOI222_X1 U44 ( .A1(add_2071_SUM_17_), .A2(n17117), .B1(n16672), .B2(n17114), 
        .C1(n54), .C2(n63), .ZN(n62) );
  INV_X1 U45 ( .A(n64), .ZN(n63) );
  OAI211_X1 U46 ( .C1(n5236), .C2(n37), .A(n52), .B(n65), .ZN(n5663) );
  AOI222_X1 U47 ( .A1(add_2071_SUM_16_), .A2(n17117), .B1(n16710), .B2(n17114), 
        .C1(n54), .C2(n66), .ZN(n65) );
  OAI211_X1 U48 ( .C1(n5235), .C2(n37), .A(n52), .B(n67), .ZN(n5664) );
  AOI222_X1 U49 ( .A1(add_2071_SUM_15_), .A2(n17117), .B1(n16711), .B2(n17114), 
        .C1(n54), .C2(n68), .ZN(n67) );
  OAI211_X1 U50 ( .C1(n5114), .C2(n37), .A(n52), .B(n69), .ZN(n5665) );
  AOI222_X1 U51 ( .A1(add_2071_SUM_18_), .A2(n17117), .B1(n16709), .B2(n17114), 
        .C1(n54), .C2(n70), .ZN(n69) );
  AOI21_X1 U52 ( .B1(n54), .B2(n71), .A(n17120), .ZN(n52) );
  OAI211_X1 U53 ( .C1(n72), .C2(n29), .A(n73), .B(n74), .ZN(n5666) );
  AOI22_X1 U54 ( .A1(add_2071_SUM_28_), .A2(n17117), .B1(n17111), .B2(
        vis_pc_o[28]), .ZN(n74) );
  AOI21_X1 U55 ( .B1(n16693), .B2(n17115), .A(n17120), .ZN(n73) );
  OAI211_X1 U56 ( .C1(n76), .C2(n29), .A(n77), .B(n78), .ZN(n5667) );
  AOI22_X1 U57 ( .A1(add_2071_SUM_27_), .A2(n17118), .B1(n17111), .B2(
        vis_pc_o[27]), .ZN(n78) );
  AOI21_X1 U58 ( .B1(n16695), .B2(n17115), .A(n17121), .ZN(n77) );
  OAI22_X1 U59 ( .A1(n80), .A2(n17126), .B1(n82), .B2(n83), .ZN(n5668) );
  AOI21_X1 U61 ( .B1(n84), .B2(n85), .A(n17127), .ZN(n82) );
  AOI221_X1 U62 ( .B1(n86), .B2(n87), .C1(n88), .C2(n89), .A(n90), .ZN(n80) );
  AND3_X1 U63 ( .A1(n91), .A2(n92), .A3(n84), .ZN(n90) );
  OAI33_X1 U64 ( .A1(n27), .A2(U186_Z_0), .A3(n4949), .B1(n93), .B2(n16688), 
        .B3(n94), .ZN(n91) );
  INV_X1 U65 ( .A(n76), .ZN(n87) );
  OAI211_X1 U66 ( .C1(n95), .C2(n29), .A(n96), .B(n97), .ZN(n5669) );
  AOI22_X1 U67 ( .A1(add_2071_SUM_26_), .A2(n17118), .B1(n17111), .B2(
        vis_pc_o[26]), .ZN(n97) );
  AOI21_X1 U69 ( .B1(n16698), .B2(n17115), .A(n17120), .ZN(n96) );
  INV_X1 U70 ( .A(n99), .ZN(n95) );
  OAI211_X1 U71 ( .C1(n100), .C2(n29), .A(n101), .B(n102), .ZN(n5670) );
  AOI22_X1 U72 ( .A1(add_2071_SUM_25_), .A2(n17118), .B1(n17111), .B2(
        vis_pc_o[25]), .ZN(n102) );
  AOI21_X1 U74 ( .B1(n16663), .B2(n17115), .A(n17120), .ZN(n101) );
  OAI211_X1 U75 ( .C1(n104), .C2(n29), .A(n105), .B(n106), .ZN(n5671) );
  AOI22_X1 U76 ( .A1(add_2071_SUM_24_), .A2(n17118), .B1(n17111), .B2(
        vis_pc_o[24]), .ZN(n106) );
  AOI21_X1 U78 ( .B1(n16655), .B2(n17115), .A(n17120), .ZN(n105) );
  INV_X1 U79 ( .A(n108), .ZN(n104) );
  OAI211_X1 U80 ( .C1(n109), .C2(n29), .A(n110), .B(n111), .ZN(n5672) );
  AOI22_X1 U81 ( .A1(add_2071_SUM_23_), .A2(n17118), .B1(n17111), .B2(
        vis_pc_o[23]), .ZN(n111) );
  AOI21_X1 U82 ( .B1(n16701), .B2(n17115), .A(n17120), .ZN(n110) );
  OAI211_X1 U83 ( .C1(n113), .C2(n29), .A(n114), .B(n115), .ZN(n5673) );
  AOI22_X1 U84 ( .A1(add_2071_SUM_29_), .A2(n17118), .B1(n17111), .B2(
        vis_pc_o[29]), .ZN(n115) );
  AOI21_X1 U86 ( .B1(add_2073_SUM_31_), .B2(n17115), .A(n17121), .ZN(n114) );
  INV_X1 U87 ( .A(n117), .ZN(n113) );
  OAI211_X1 U88 ( .C1(n118), .C2(n29), .A(n119), .B(n120), .ZN(n5674) );
  AOI22_X1 U89 ( .A1(add_2071_SUM_12_), .A2(n17118), .B1(n17111), .B2(
        vis_pc_o[12]), .ZN(n120) );
  AOI21_X1 U91 ( .B1(n16679), .B2(n17115), .A(n17121), .ZN(n119) );
  OAI211_X1 U92 ( .C1(n122), .C2(n29), .A(n123), .B(n124), .ZN(n5675) );
  AOI22_X1 U93 ( .A1(add_2071_SUM_10_), .A2(n17118), .B1(n17111), .B2(
        vis_pc_o[10]), .ZN(n124) );
  AOI21_X1 U95 ( .B1(n16719), .B2(n17115), .A(n17121), .ZN(n123) );
  INV_X1 U96 ( .A(n126), .ZN(n122) );
  OAI211_X1 U97 ( .C1(n127), .C2(n29), .A(n128), .B(n129), .ZN(n5676) );
  AOI22_X1 U98 ( .A1(add_2071_SUM_8_), .A2(n17118), .B1(n17112), .B2(
        vis_pc_o[8]), .ZN(n129) );
  AOI21_X1 U100 ( .B1(n16727), .B2(n17115), .A(n17121), .ZN(n128) );
  OAI211_X1 U101 ( .C1(n131), .C2(n29), .A(n132), .B(n133), .ZN(n5677) );
  AOI22_X1 U102 ( .A1(add_2071_SUM_13_), .A2(n17118), .B1(n17112), .B2(
        vis_pc_o[13]), .ZN(n133) );
  AOI21_X1 U104 ( .B1(n16658), .B2(n17115), .A(n17121), .ZN(n132) );
  INV_X1 U105 ( .A(n135), .ZN(n131) );
  OAI211_X1 U106 ( .C1(n136), .C2(n29), .A(n137), .B(n138), .ZN(n5678) );
  AOI22_X1 U107 ( .A1(add_2071_SUM_11_), .A2(n17118), .B1(n17112), .B2(
        vis_pc_o[11]), .ZN(n138) );
  AOI21_X1 U109 ( .B1(n16653), .B2(n17116), .A(n17121), .ZN(n137) );
  OAI211_X1 U110 ( .C1(n140), .C2(n29), .A(n141), .B(n142), .ZN(n5679) );
  AOI22_X1 U111 ( .A1(add_2071_SUM_9_), .A2(n17119), .B1(n17112), .B2(
        vis_pc_o[9]), .ZN(n142) );
  AOI21_X1 U113 ( .B1(n16723), .B2(n17116), .A(n17121), .ZN(n141) );
  OAI211_X1 U114 ( .C1(n144), .C2(n29), .A(n145), .B(n146), .ZN(n5680) );
  AOI22_X1 U115 ( .A1(add_2071_SUM_7_), .A2(n17119), .B1(n17112), .B2(
        vis_pc_o[7]), .ZN(n146) );
  AOI21_X1 U116 ( .B1(n16722), .B2(n17115), .A(n17121), .ZN(n145) );
  OAI211_X1 U117 ( .C1(n148), .C2(n29), .A(n149), .B(n150), .ZN(n5681) );
  AOI22_X1 U118 ( .A1(add_2071_SUM_5_), .A2(n17119), .B1(n17112), .B2(
        vis_pc_o[5]), .ZN(n150) );
  AOI21_X1 U119 ( .B1(add_2073_SUM_7_), .B2(n17116), .A(n17121), .ZN(n149) );
  OAI211_X1 U120 ( .C1(n152), .C2(n29), .A(n153), .B(n154), .ZN(n5682) );
  AOI22_X1 U121 ( .A1(add_2071_SUM_4_), .A2(n17119), .B1(n17112), .B2(
        vis_pc_o[4]), .ZN(n154) );
  AOI21_X1 U122 ( .B1(n16731), .B2(n17116), .A(n17121), .ZN(n153) );
  OAI222_X1 U123 ( .A1(n152), .A2(n156), .B1(n5240), .B2(n157), .C1(n158), 
        .C2(n159), .ZN(n5683) );
  OAI211_X1 U125 ( .C1(n160), .C2(n29), .A(n161), .B(n162), .ZN(n5684) );
  AOI22_X1 U126 ( .A1(add_2071_SUM_3_), .A2(n17119), .B1(n17112), .B2(
        vis_pc_o[3]), .ZN(n162) );
  AOI21_X1 U127 ( .B1(n16730), .B2(n17116), .A(n17121), .ZN(n161) );
  OAI222_X1 U128 ( .A1(n160), .A2(n156), .B1(n157), .B2(n164), .C1(n158), .C2(
        n165), .ZN(n5685) );
  OAI211_X1 U129 ( .C1(n166), .C2(n29), .A(n167), .B(n168), .ZN(n5686) );
  AOI22_X1 U130 ( .A1(add_2071_SUM_2_), .A2(n17119), .B1(n17112), .B2(
        vis_pc_o[2]), .ZN(n168) );
  AOI21_X1 U131 ( .B1(n16682), .B2(n17116), .A(n17121), .ZN(n167) );
  OAI222_X1 U132 ( .A1(n166), .A2(n156), .B1(n5099), .B2(n157), .C1(n158), 
        .C2(n170), .ZN(n5687) );
  OAI211_X1 U133 ( .C1(n171), .C2(n29), .A(n172), .B(n173), .ZN(n5688) );
  AOI22_X1 U134 ( .A1(add_2071_SUM_1_), .A2(n17117), .B1(n17112), .B2(
        vis_pc_o[1]), .ZN(n173) );
  AOI21_X1 U136 ( .B1(n16729), .B2(n17114), .A(n17120), .ZN(n172) );
  OAI222_X1 U138 ( .A1(n171), .A2(n156), .B1(n157), .B2(n175), .C1(n158), .C2(
        n176), .ZN(n5689) );
  OAI221_X1 U139 ( .B1(n36), .B2(vis_pc_o[0]), .C1(n4973), .C2(n37), .A(n178), 
        .ZN(n5690) );
  AOI221_X1 U140 ( .B1(n54), .B2(n179), .C1(n16732), .C2(n17114), .A(n17120), 
        .ZN(n178) );
  OAI221_X1 U142 ( .B1(n181), .B2(n182), .C1(n183), .C2(n184), .A(n185), .ZN(
        n180) );
  OR2_X1 U143 ( .A1(n186), .A2(n5234), .ZN(n182) );
  NAND2_X1 U146 ( .A1(n189), .A2(n37), .ZN(n36) );
  OAI222_X1 U147 ( .A1(n190), .A2(n156), .B1(n5025), .B2(n157), .C1(n158), 
        .C2(n191), .ZN(n5691) );
  OAI222_X1 U148 ( .A1(n192), .A2(n156), .B1(n4966), .B2(n157), .C1(n158), 
        .C2(n186), .ZN(n5692) );
  NAND2_X1 U149 ( .A1(n193), .A2(n194), .ZN(n157) );
  NAND2_X1 U150 ( .A1(n158), .A2(n195), .ZN(n156) );
  INV_X1 U151 ( .A(n196), .ZN(n158) );
  NAND2_X1 U152 ( .A1(n197), .A2(n198), .ZN(n5693) );
  OAI221_X1 U153 ( .B1(n199), .B2(n200), .C1(n201), .C2(n202), .A(n203), .ZN(
        n198) );
  INV_X1 U154 ( .A(n204), .ZN(n197) );
  OAI21_X1 U155 ( .B1(n205), .B2(n202), .A(n206), .ZN(n5694) );
  OAI221_X1 U156 ( .B1(n207), .B2(n200), .C1(n208), .C2(n202), .A(n209), .ZN(
        n206) );
  OAI21_X1 U157 ( .B1(n210), .B2(n211), .A(n212), .ZN(n5695) );
  OAI21_X1 U158 ( .B1(n213), .B2(n210), .A(n214), .ZN(n212) );
  OAI21_X1 U160 ( .B1(n215), .B2(n211), .A(n216), .ZN(n5696) );
  OAI21_X1 U161 ( .B1(n215), .B2(n213), .A(n217), .ZN(n216) );
  OAI21_X1 U162 ( .B1(n211), .B2(n218), .A(n219), .ZN(n5697) );
  OAI21_X1 U163 ( .B1(n213), .B2(n218), .A(n220), .ZN(n219) );
  OAI21_X1 U164 ( .B1(n211), .B2(n221), .A(n222), .ZN(n5698) );
  OAI21_X1 U165 ( .B1(n213), .B2(n221), .A(n223), .ZN(n222) );
  OAI21_X1 U166 ( .B1(n211), .B2(n224), .A(n225), .ZN(n5699) );
  OAI21_X1 U167 ( .B1(n213), .B2(n224), .A(n4799), .ZN(n225) );
  OAI21_X1 U168 ( .B1(n211), .B2(n226), .A(n227), .ZN(n5700) );
  OAI21_X1 U169 ( .B1(n213), .B2(n226), .A(n228), .ZN(n227) );
  OAI21_X1 U170 ( .B1(n211), .B2(n229), .A(n230), .ZN(n5701) );
  OAI21_X1 U171 ( .B1(n213), .B2(n229), .A(n231), .ZN(n230) );
  OAI22_X1 U172 ( .A1(n232), .A2(n211), .B1(n4796), .B2(n233), .ZN(n5702) );
  NOR2_X1 U173 ( .A1(n232), .A2(n213), .ZN(n233) );
  OAI22_X1 U174 ( .A1(n234), .A2(n211), .B1(n5578), .B2(n235), .ZN(n5703) );
  NOR2_X1 U175 ( .A1(n234), .A2(n213), .ZN(n235) );
  OAI22_X1 U176 ( .A1(n236), .A2(n211), .B1(n5537), .B2(n237), .ZN(n5704) );
  NOR2_X1 U177 ( .A1(n236), .A2(n213), .ZN(n237) );
  OAI22_X1 U178 ( .A1(n238), .A2(n211), .B1(n5570), .B2(n239), .ZN(n5705) );
  NOR2_X1 U179 ( .A1(n238), .A2(n213), .ZN(n239) );
  OAI22_X1 U180 ( .A1(n240), .A2(n211), .B1(n4795), .B2(n241), .ZN(n5706) );
  NOR2_X1 U181 ( .A1(n240), .A2(n213), .ZN(n241) );
  OAI22_X1 U182 ( .A1(n242), .A2(n211), .B1(n243), .B2(n244), .ZN(n5707) );
  NOR2_X1 U183 ( .A1(n242), .A2(n213), .ZN(n243) );
  OAI22_X1 U184 ( .A1(n211), .A2(n245), .B1(n5538), .B2(n246), .ZN(n5708) );
  NOR2_X1 U185 ( .A1(n213), .A2(n245), .ZN(n246) );
  OAI22_X1 U186 ( .A1(n211), .A2(n247), .B1(n5539), .B2(n248), .ZN(n5709) );
  NOR2_X1 U187 ( .A1(n213), .A2(n247), .ZN(n248) );
  OAI22_X1 U188 ( .A1(n211), .A2(n249), .B1(n5540), .B2(n250), .ZN(n5710) );
  NOR2_X1 U189 ( .A1(n213), .A2(n249), .ZN(n250) );
  OAI211_X1 U192 ( .C1(n4905), .C2(n17122), .A(n254), .B(n255), .ZN(n5711) );
  OAI21_X1 U193 ( .B1(haddr_o[7]), .B2(haddr_o[2]), .A(n256), .ZN(n254) );
  OAI33_X1 U194 ( .A1(n257), .A2(n5068), .A3(n258), .B1(n259), .B2(n5516), 
        .B3(n260), .ZN(n5712) );
  NOR3_X1 U195 ( .A1(n253), .A2(n251), .A3(n261), .ZN(n257) );
  OAI221_X1 U196 ( .B1(n262), .B2(n17109), .C1(n264), .C2(n17107), .A(n266), 
        .ZN(n5713) );
  NAND2_X1 U199 ( .A1(sub_2068_SUM_22_), .A2(n17106), .ZN(n269) );
  OAI221_X1 U201 ( .B1(n5625), .B2(n17109), .C1(n270), .C2(n17107), .A(n271), 
        .ZN(n5715) );
  NAND2_X1 U202 ( .A1(sub_2068_SUM_21_), .A2(n17106), .ZN(n271) );
  OAI221_X1 U203 ( .B1(n5618), .B2(n17109), .C1(n272), .C2(n265), .A(n273), 
        .ZN(n5716) );
  NAND2_X1 U204 ( .A1(sub_2068_SUM_20_), .A2(n17106), .ZN(n273) );
  OAI221_X1 U205 ( .B1(n5033), .B2(n17109), .C1(n274), .C2(n265), .A(n275), 
        .ZN(n5717) );
  NAND2_X1 U206 ( .A1(sub_2068_SUM_19_), .A2(n17106), .ZN(n275) );
  OAI221_X1 U207 ( .B1(n5067), .B2(n17109), .C1(n276), .C2(n265), .A(n277), 
        .ZN(n5718) );
  NAND2_X1 U208 ( .A1(sub_2068_SUM_18_), .A2(n17106), .ZN(n277) );
  OAI221_X1 U209 ( .B1(n5639), .B2(n17109), .C1(n278), .C2(n17107), .A(n279), 
        .ZN(n5719) );
  NAND2_X1 U210 ( .A1(sub_2068_SUM_17_), .A2(n17106), .ZN(n279) );
  NAND2_X1 U212 ( .A1(sub_2068_SUM_16_), .A2(n17106), .ZN(n281) );
  OAI221_X1 U214 ( .B1(n5505), .B2(n17109), .C1(n282), .C2(n265), .A(n283), 
        .ZN(n5721) );
  NAND2_X1 U215 ( .A1(sub_2068_SUM_15_), .A2(n17106), .ZN(n283) );
  OAI221_X1 U216 ( .B1(n5506), .B2(n17109), .C1(n284), .C2(n265), .A(n285), 
        .ZN(n5722) );
  NAND2_X1 U217 ( .A1(sub_2068_SUM_14_), .A2(n17106), .ZN(n285) );
  OAI221_X1 U218 ( .B1(n5600), .B2(n17109), .C1(n286), .C2(n265), .A(n287), 
        .ZN(n5723) );
  NAND2_X1 U219 ( .A1(sub_2068_SUM_13_), .A2(n17106), .ZN(n287) );
  OAI221_X1 U220 ( .B1(n5507), .B2(n17110), .C1(n288), .C2(n17107), .A(n289), 
        .ZN(n5724) );
  NAND2_X1 U221 ( .A1(sub_2068_SUM_12_), .A2(n17106), .ZN(n289) );
  NAND2_X1 U223 ( .A1(sub_2068_SUM_11_), .A2(n17105), .ZN(n291) );
  NAND2_X1 U226 ( .A1(sub_2068_SUM_10_), .A2(n17105), .ZN(n293) );
  OAI221_X1 U228 ( .B1(n5579), .B2(n17110), .C1(n294), .C2(n17107), .A(n295), 
        .ZN(n5727) );
  NAND2_X1 U229 ( .A1(sub_2068_SUM_9_), .A2(n17105), .ZN(n295) );
  OAI221_X1 U230 ( .B1(n5581), .B2(n17110), .C1(n296), .C2(n17107), .A(n297), 
        .ZN(n5728) );
  NAND2_X1 U231 ( .A1(sub_2068_SUM_8_), .A2(n17105), .ZN(n297) );
  OAI221_X1 U232 ( .B1(n5520), .B2(n17110), .C1(n298), .C2(n17107), .A(n299), 
        .ZN(n5729) );
  NAND2_X1 U233 ( .A1(sub_2068_SUM_7_), .A2(n17105), .ZN(n299) );
  NAND2_X1 U235 ( .A1(sub_2068_SUM_6_), .A2(n17105), .ZN(n301) );
  NAND2_X1 U238 ( .A1(sub_2068_SUM_5_), .A2(n17105), .ZN(n303) );
  NAND2_X1 U241 ( .A1(sub_2068_SUM_4_), .A2(n17105), .ZN(n305) );
  OAI221_X1 U243 ( .B1(n5513), .B2(n17110), .C1(n306), .C2(n17107), .A(n307), 
        .ZN(n5733) );
  NAND2_X1 U244 ( .A1(sub_2068_SUM_3_), .A2(n17105), .ZN(n307) );
  OAI221_X1 U245 ( .B1(n5512), .B2(n17110), .C1(n308), .C2(n265), .A(n309), 
        .ZN(n5734) );
  NAND2_X1 U246 ( .A1(sub_2068_SUM_2_), .A2(n17105), .ZN(n309) );
  OAI221_X1 U247 ( .B1(n5511), .B2(n17109), .C1(n310), .C2(n265), .A(n311), 
        .ZN(n5735) );
  NAND2_X1 U248 ( .A1(sub_2068_SUM_1_), .A2(n17105), .ZN(n311) );
  OAI222_X1 U249 ( .A1(n5510), .A2(n17110), .B1(sub_2068_A_0_), .B2(n16647), 
        .C1(n260), .C2(n17107), .ZN(n5736) );
  INV_X1 U252 ( .A(n315), .ZN(n258) );
  NOR2_X1 U255 ( .A1(n259), .A2(sub_2068_A_0_), .ZN(n314) );
  NAND2_X1 U256 ( .A1(n5516), .A2(n315), .ZN(n265) );
  NAND2_X1 U257 ( .A1(n316), .A2(n253), .ZN(n315) );
  OAI221_X1 U258 ( .B1(n317), .B2(n17103), .C1(n4971), .C2(n17102), .A(n320), 
        .ZN(n5737) );
  AOI22_X1 U259 ( .A1(n16738), .A2(vis_pc_o[23]), .B1(n322), .B2(vis_tbit_o), 
        .ZN(n320) );
  OAI221_X1 U261 ( .B1(n186), .B2(n324), .C1(n5101), .C2(n17101), .A(n325), 
        .ZN(n5738) );
  OAI21_X1 U262 ( .B1(n326), .B2(n327), .A(n17104), .ZN(n325) );
  AOI21_X1 U263 ( .B1(n329), .B2(n330), .A(n4922), .ZN(n326) );
  NAND3_X1 U264 ( .A1(n16657), .A2(n16686), .A3(n333), .ZN(n330) );
  OAI221_X1 U265 ( .B1(n334), .B2(n335), .C1(n16803), .C2(n336), .A(n337), 
        .ZN(n5739) );
  AOI222_X1 U266 ( .A1(n338), .A2(n339), .B1(n16646), .B2(hrdata_i[30]), .C1(
        n341), .C2(hrdata_i[14]), .ZN(n337) );
  OAI221_X1 U268 ( .B1(n3), .B2(n334), .C1(n16795), .C2(n336), .A(n342), .ZN(
        n5740) );
  AOI222_X1 U269 ( .A1(n338), .A2(n343), .B1(n16646), .B2(hrdata_i[28]), .C1(
        n341), .C2(hrdata_i[12]), .ZN(n342) );
  OAI221_X1 U271 ( .B1(n4), .B2(n334), .C1(n16814), .C2(n336), .A(n344), .ZN(
        n5741) );
  AOI222_X1 U272 ( .A1(n338), .A2(n345), .B1(n16646), .B2(hrdata_i[27]), .C1(
        n341), .C2(hrdata_i[11]), .ZN(n344) );
  OAI221_X1 U274 ( .B1(n5), .B2(n334), .C1(n16815), .C2(n336), .A(n346), .ZN(
        n5742) );
  AOI222_X1 U275 ( .A1(n338), .A2(n347), .B1(n16646), .B2(hrdata_i[26]), .C1(
        n341), .C2(hrdata_i[10]), .ZN(n346) );
  OAI221_X1 U277 ( .B1(n6), .B2(n334), .C1(n16796), .C2(n336), .A(n348), .ZN(
        n5743) );
  AOI222_X1 U278 ( .A1(n338), .A2(n349), .B1(n16646), .B2(hrdata_i[25]), .C1(
        n341), .C2(hrdata_i[9]), .ZN(n348) );
  OAI221_X1 U280 ( .B1(n7), .B2(n334), .C1(n16797), .C2(n336), .A(n350), .ZN(
        n5744) );
  AOI222_X1 U281 ( .A1(n338), .A2(n351), .B1(n16646), .B2(hrdata_i[24]), .C1(
        n341), .C2(hrdata_i[8]), .ZN(n350) );
  OAI221_X1 U283 ( .B1(n8), .B2(n334), .C1(n16799), .C2(n336), .A(n352), .ZN(
        n5745) );
  AOI222_X1 U284 ( .A1(n338), .A2(n353), .B1(n16646), .B2(hrdata_i[23]), .C1(
        n341), .C2(hrdata_i[7]), .ZN(n352) );
  OAI221_X1 U286 ( .B1(n9), .B2(n334), .C1(n16801), .C2(n336), .A(n354), .ZN(
        n5746) );
  AOI222_X1 U287 ( .A1(n338), .A2(n355), .B1(n16646), .B2(hrdata_i[22]), .C1(
        n341), .C2(hrdata_i[6]), .ZN(n354) );
  OAI221_X1 U289 ( .B1(n5240), .B2(n334), .C1(n5244), .C2(n336), .A(n356), 
        .ZN(n5747) );
  AOI222_X1 U290 ( .A1(n338), .A2(n357), .B1(n16646), .B2(hrdata_i[21]), .C1(
        n341), .C2(hrdata_i[5]), .ZN(n356) );
  OAI221_X1 U292 ( .B1(n164), .B2(n334), .C1(n5243), .C2(n336), .A(n358), .ZN(
        n5748) );
  AOI222_X1 U293 ( .A1(n338), .A2(n359), .B1(n16646), .B2(hrdata_i[20]), .C1(
        n341), .C2(hrdata_i[4]), .ZN(n358) );
  OAI221_X1 U295 ( .B1(n5099), .B2(n334), .C1(n16794), .C2(n336), .A(n360), 
        .ZN(n5749) );
  AOI222_X1 U296 ( .A1(n338), .A2(n361), .B1(n16646), .B2(hrdata_i[19]), .C1(
        n341), .C2(hrdata_i[3]), .ZN(n360) );
  OAI221_X1 U298 ( .B1(n175), .B2(n334), .C1(n5241), .C2(n336), .A(n362), .ZN(
        n5750) );
  AOI222_X1 U299 ( .A1(n338), .A2(n363), .B1(n16646), .B2(hrdata_i[18]), .C1(
        n341), .C2(hrdata_i[2]), .ZN(n362) );
  OAI221_X1 U301 ( .B1(n5025), .B2(n334), .C1(n5026), .C2(n336), .A(n364), 
        .ZN(n5751) );
  AOI222_X1 U302 ( .A1(n338), .A2(n365), .B1(n16646), .B2(hrdata_i[17]), .C1(
        n341), .C2(hrdata_i[1]), .ZN(n364) );
  OAI221_X1 U304 ( .B1(n4966), .B2(n334), .C1(n4967), .C2(n336), .A(n366), 
        .ZN(n5752) );
  AOI222_X1 U305 ( .A1(n338), .A2(n367), .B1(n16646), .B2(hrdata_i[16]), .C1(
        n341), .C2(hrdata_i[0]), .ZN(n366) );
  OAI221_X1 U307 ( .B1(n2), .B2(n334), .C1(n16807), .C2(n336), .A(n368), .ZN(
        n5753) );
  AOI222_X1 U308 ( .A1(n338), .A2(n369), .B1(n16646), .B2(hrdata_i[29]), .C1(
        n341), .C2(hrdata_i[13]), .ZN(n368) );
  OAI221_X1 U310 ( .B1(n334), .B2(n370), .C1(n16811), .C2(n336), .A(n371), 
        .ZN(n5754) );
  AOI222_X1 U311 ( .A1(n338), .A2(n372), .B1(n16646), .B2(hrdata_i[31]), .C1(
        n341), .C2(hrdata_i[15]), .ZN(n371) );
  NAND2_X1 U314 ( .A1(n16869), .A2(vis_pc_o[0]), .ZN(n374) );
  OAI22_X1 U317 ( .A1(n335), .A2(n379), .B1(n380), .B2(n381), .ZN(n5755) );
  INV_X1 U318 ( .A(hrdata_i[14]), .ZN(n380) );
  OAI221_X1 U320 ( .B1(n382), .B2(n381), .C1(n2), .C2(n379), .A(n383), .ZN(
        n5756) );
  NAND2_X1 U321 ( .A1(sub_2069_SUM_8_), .A2(n384), .ZN(n383) );
  OAI221_X1 U322 ( .B1(n385), .B2(n381), .C1(n3), .C2(n379), .A(n386), .ZN(
        n5757) );
  NAND2_X1 U323 ( .A1(sub_2069_SUM_7_), .A2(n384), .ZN(n386) );
  INV_X1 U324 ( .A(hrdata_i[12]), .ZN(n385) );
  OAI221_X1 U325 ( .B1(n387), .B2(n381), .C1(n4), .C2(n379), .A(n388), .ZN(
        n5758) );
  NAND2_X1 U326 ( .A1(sub_2069_SUM_6_), .A2(n384), .ZN(n388) );
  INV_X1 U327 ( .A(hrdata_i[11]), .ZN(n387) );
  OAI221_X1 U328 ( .B1(n389), .B2(n381), .C1(n5), .C2(n379), .A(n390), .ZN(
        n5759) );
  NAND2_X1 U329 ( .A1(sub_2069_SUM_5_), .A2(n384), .ZN(n390) );
  INV_X1 U330 ( .A(hrdata_i[10]), .ZN(n389) );
  OAI221_X1 U331 ( .B1(n391), .B2(n381), .C1(n6), .C2(n379), .A(n392), .ZN(
        n5760) );
  NAND2_X1 U332 ( .A1(sub_2069_SUM_4_), .A2(n384), .ZN(n392) );
  OAI221_X1 U333 ( .B1(n393), .B2(n381), .C1(n7), .C2(n379), .A(n394), .ZN(
        n5761) );
  NAND2_X1 U334 ( .A1(sub_2069_SUM_3_), .A2(n384), .ZN(n394) );
  OAI221_X1 U335 ( .B1(n395), .B2(n381), .C1(n8), .C2(n379), .A(n396), .ZN(
        n5762) );
  NAND2_X1 U336 ( .A1(sub_2069_SUM_2_), .A2(n384), .ZN(n396) );
  INV_X1 U337 ( .A(hrdata_i[7]), .ZN(n395) );
  OAI221_X1 U338 ( .B1(n397), .B2(n381), .C1(n9), .C2(n379), .A(n398), .ZN(
        n5763) );
  NAND2_X1 U339 ( .A1(sub_2069_SUM_1_), .A2(n384), .ZN(n398) );
  AOI21_X1 U340 ( .B1(n399), .B2(n5648), .A(n400), .ZN(n384) );
  OR4_X1 U341 ( .A1(n401), .A2(n402), .A3(n403), .A4(n404), .ZN(n399) );
  XOR2_X1 U342 ( .A(n405), .B(n406), .Z(n404) );
  NOR2_X1 U343 ( .A1(n5034), .A2(n164), .ZN(n406) );
  XOR2_X1 U344 ( .A(n4804), .B(n407), .Z(n402) );
  OAI221_X1 U345 ( .B1(n408), .B2(n409), .C1(n5025), .C2(n410), .A(n411), .ZN(
        n401) );
  AOI21_X1 U346 ( .B1(n412), .B2(n413), .A(n414), .ZN(n411) );
  XOR2_X1 U347 ( .A(n415), .B(n416), .Z(n414) );
  AOI21_X1 U348 ( .B1(n4966), .B2(n417), .A(n410), .ZN(n409) );
  AOI211_X1 U349 ( .C1(n4966), .C2(n417), .A(n5025), .B(n5034), .ZN(n408) );
  OAI22_X1 U350 ( .A1(n5240), .A2(n418), .B1(n419), .B2(n381), .ZN(n5764) );
  INV_X1 U351 ( .A(hrdata_i[5]), .ZN(n419) );
  OAI222_X1 U352 ( .A1(n164), .A2(n418), .B1(n420), .B2(n381), .C1(n421), .C2(
        n422), .ZN(n5765) );
  OAI222_X1 U354 ( .A1(n5099), .A2(n418), .B1(n423), .B2(n381), .C1(n424), 
        .C2(n422), .ZN(n5766) );
  OAI222_X1 U355 ( .A1(n175), .A2(n418), .B1(n425), .B2(n381), .C1(n426), .C2(
        n422), .ZN(n5767) );
  OAI222_X1 U356 ( .A1(n5025), .A2(n418), .B1(n427), .B2(n381), .C1(n428), 
        .C2(n422), .ZN(n5768) );
  INV_X1 U357 ( .A(n410), .ZN(n428) );
  OAI222_X1 U358 ( .A1(n4966), .A2(n418), .B1(n429), .B2(n381), .C1(n412), 
        .C2(n422), .ZN(n5769) );
  OAI21_X1 U360 ( .B1(n430), .B2(n431), .A(n422), .ZN(n418) );
  OAI221_X1 U361 ( .B1(n432), .B2(n433), .C1(n5254), .C2(n434), .A(n435), .ZN(
        n5770) );
  AOI21_X1 U362 ( .B1(n436), .B2(n437), .A(n433), .ZN(n434) );
  AOI221_X1 U363 ( .B1(n438), .B2(n16734), .C1(n440), .C2(n16817), .A(n442), 
        .ZN(n432) );
  OAI33_X1 U364 ( .A1(n443), .A2(n16795), .A3(n444), .B1(n16681), .B2(n16814), 
        .B3(n445), .ZN(n442) );
  OAI221_X1 U365 ( .B1(n446), .B2(n433), .C1(n5162), .C2(n447), .A(n435), .ZN(
        n5771) );
  AOI222_X1 U366 ( .A1(n440), .A2(n16798), .B1(n449), .B2(n17098), .C1(n450), 
        .C2(n451), .ZN(n446) );
  OAI221_X1 U367 ( .B1(n5253), .B2(n452), .C1(n453), .C2(n433), .A(n435), .ZN(
        n5772) );
  AOI222_X1 U368 ( .A1(n440), .A2(n16657), .B1(n449), .B2(n16817), .C1(n450), 
        .C2(n454), .ZN(n453) );
  AOI21_X1 U369 ( .B1(n436), .B2(n455), .A(n433), .ZN(n452) );
  OAI221_X1 U370 ( .B1(n5003), .B2(n456), .C1(n457), .C2(n433), .A(n435), .ZN(
        n5773) );
  NAND2_X1 U371 ( .A1(n447), .A2(n458), .ZN(n435) );
  OAI21_X1 U372 ( .B1(n16799), .B2(n459), .A(n460), .ZN(n458) );
  INV_X1 U373 ( .A(n433), .ZN(n447) );
  AOI222_X1 U374 ( .A1(n440), .A2(n17098), .B1(n449), .B2(n16657), .C1(n450), 
        .C2(n461), .ZN(n457) );
  NAND3_X1 U375 ( .A1(n462), .A2(n463), .A3(n464), .ZN(n450) );
  AOI21_X1 U376 ( .B1(n465), .B2(n466), .A(n438), .ZN(n464) );
  NAND2_X1 U377 ( .A1(n467), .A2(n468), .ZN(n438) );
  NAND3_X1 U378 ( .A1(n469), .A2(n16725), .A3(n471), .ZN(n467) );
  AOI21_X1 U379 ( .B1(n16733), .B2(n16657), .A(n443), .ZN(n471) );
  OAI211_X1 U380 ( .C1(n473), .C2(n474), .A(n16819), .B(n475), .ZN(n463) );
  NAND3_X1 U381 ( .A1(n16816), .A2(n16725), .A3(n476), .ZN(n462) );
  OAI221_X1 U382 ( .B1(n477), .B2(n443), .C1(n478), .C2(n479), .A(n480), .ZN(
        n449) );
  AOI22_X1 U383 ( .A1(n16819), .A2(n481), .B1(n482), .B2(n466), .ZN(n480) );
  INV_X1 U384 ( .A(n445), .ZN(n481) );
  NOR2_X1 U385 ( .A1(n483), .A2(n484), .ZN(n445) );
  NOR2_X1 U386 ( .A1(n485), .A2(n16795), .ZN(n477) );
  AOI21_X1 U387 ( .B1(n436), .B2(n486), .A(n433), .ZN(n456) );
  NAND2_X1 U388 ( .A1(n17124), .A2(n487), .ZN(n433) );
  NAND4_X1 U389 ( .A1(n488), .A2(n489), .A3(n490), .A4(n491), .ZN(n487) );
  NOR4_X1 U390 ( .A1(n492), .A2(n493), .A3(n494), .A4(n495), .ZN(n491) );
  OAI221_X1 U391 ( .B1(n496), .B2(n497), .C1(n498), .C2(n499), .A(n500), .ZN(
        n492) );
  NAND4_X1 U392 ( .A1(n483), .A2(n501), .A3(n502), .A4(n503), .ZN(n500) );
  AOI21_X1 U393 ( .B1(n504), .B2(n16817), .A(n505), .ZN(n496) );
  AOI221_X1 U394 ( .B1(n506), .B2(n507), .C1(n508), .C2(n16802), .A(n510), 
        .ZN(n490) );
  OAI211_X1 U395 ( .C1(n16733), .C2(n329), .A(n511), .B(n512), .ZN(n508) );
  NAND3_X1 U396 ( .A1(n16733), .A2(n16871), .A3(n16811), .ZN(n511) );
  AOI21_X1 U397 ( .B1(n514), .B2(n17097), .A(n515), .ZN(n436) );
  OAI22_X1 U398 ( .A1(n16854), .A2(n17122), .B1(n516), .B2(n17126), .ZN(n5774)
         );
  NOR4_X1 U399 ( .A1(n517), .A2(n518), .A3(n519), .A4(n520), .ZN(n516) );
  OAI221_X1 U400 ( .B1(n16858), .B2(n522), .C1(n16864), .C2(n524), .A(n525), 
        .ZN(n520) );
  AOI22_X1 U401 ( .A1(n526), .A2(n527), .B1(n528), .B2(n529), .ZN(n525) );
  OAI221_X1 U402 ( .B1(n16795), .B2(n530), .C1(n531), .C2(n532), .A(n533), 
        .ZN(n519) );
  AOI222_X1 U403 ( .A1(n534), .A2(n535), .B1(n536), .B2(n537), .C1(n16819), 
        .C2(n538), .ZN(n533) );
  INV_X1 U404 ( .A(n539), .ZN(n538) );
  AOI221_X1 U405 ( .B1(n540), .B2(n541), .C1(n542), .C2(n543), .A(n544), .ZN(
        n539) );
  OR2_X1 U406 ( .A1(n545), .A2(n546), .ZN(n544) );
  NAND3_X1 U407 ( .A1(n547), .A2(n548), .A3(n549), .ZN(n537) );
  NAND3_X1 U408 ( .A1(n550), .A2(n16797), .A3(n551), .ZN(n549) );
  INV_X1 U409 ( .A(n552), .ZN(n536) );
  AOI211_X1 U410 ( .C1(n466), .C2(n553), .A(n554), .B(n555), .ZN(n531) );
  AOI21_X1 U411 ( .B1(n556), .B2(n557), .A(n558), .ZN(n555) );
  OAI21_X1 U412 ( .B1(n559), .B2(n16824), .A(n16862), .ZN(n557) );
  NAND2_X1 U413 ( .A1(n560), .A2(n561), .ZN(n554) );
  NAND3_X1 U414 ( .A1(n16819), .A2(n16839), .A3(n563), .ZN(n561) );
  OAI21_X1 U415 ( .B1(n564), .B2(n565), .A(n566), .ZN(n560) );
  INV_X1 U416 ( .A(n567), .ZN(n564) );
  OAI21_X1 U417 ( .B1(n568), .B2(n569), .A(n570), .ZN(n553) );
  NAND3_X1 U418 ( .A1(n16833), .A2(n16826), .A3(n5228), .ZN(n570) );
  AOI221_X1 U419 ( .B1(n572), .B2(n573), .C1(n574), .C2(n473), .A(n575), .ZN(
        n530) );
  OAI33_X1 U420 ( .A1(n576), .A2(n5243), .A3(n577), .B1(n578), .B2(n579), .B3(
        n580), .ZN(n575) );
  NAND2_X1 U421 ( .A1(n16680), .A2(n581), .ZN(n578) );
  OAI22_X1 U422 ( .A1(n16797), .A2(n582), .B1(n16796), .B2(n583), .ZN(n581) );
  OAI21_X1 U423 ( .B1(n16801), .B2(n16812), .A(n16798), .ZN(n573) );
  OAI221_X1 U424 ( .B1(n584), .B2(n585), .C1(n16866), .C2(n586), .A(n587), 
        .ZN(n518) );
  AOI222_X1 U425 ( .A1(n588), .A2(n589), .B1(n590), .B2(n591), .C1(n592), .C2(
        n593), .ZN(n587) );
  OAI22_X1 U426 ( .A1(n594), .A2(n16734), .B1(n595), .B2(n596), .ZN(n593) );
  AOI221_X1 U427 ( .B1(n597), .B2(n16862), .C1(n16833), .C2(n598), .A(n599), 
        .ZN(n595) );
  OAI21_X1 U428 ( .B1(n16680), .B2(n16839), .A(n600), .ZN(n598) );
  OAI21_X1 U429 ( .B1(n601), .B2(n602), .A(n483), .ZN(n600) );
  INV_X1 U430 ( .A(n603), .ZN(n601) );
  OAI21_X1 U431 ( .B1(n604), .B2(n605), .A(n606), .ZN(n591) );
  INV_X1 U432 ( .A(n607), .ZN(n588) );
  AOI222_X1 U433 ( .A1(n608), .A2(n563), .B1(n609), .B2(n610), .C1(n611), .C2(
        n589), .ZN(n586) );
  AOI221_X1 U434 ( .B1(n612), .B2(n5228), .C1(n613), .C2(n614), .A(n615), .ZN(
        n584) );
  NOR2_X1 U435 ( .A1(n616), .A2(n617), .ZN(n613) );
  NAND4_X1 U436 ( .A1(n618), .A2(n619), .A3(n620), .A4(n621), .ZN(n517) );
  AOI21_X1 U437 ( .B1(n574), .B2(n622), .A(n623), .ZN(n621) );
  NOR4_X1 U438 ( .A1(n624), .A2(n579), .A3(n503), .A4(n625), .ZN(n623) );
  OAI21_X1 U439 ( .B1(n16812), .B2(n626), .A(n627), .ZN(n622) );
  AOI21_X1 U440 ( .B1(n628), .B2(n16657), .A(n629), .ZN(n626) );
  NAND4_X1 U441 ( .A1(n630), .A2(n631), .A3(n483), .A4(n632), .ZN(n620) );
  OAI22_X1 U442 ( .A1(n16869), .A2(n17122), .B1(n633), .B2(n17126), .ZN(n5775)
         );
  NOR4_X1 U443 ( .A1(n634), .A2(n635), .A3(n636), .A4(n637), .ZN(n633) );
  OAI221_X1 U444 ( .B1(n638), .B2(n639), .C1(n640), .C2(n641), .A(n642), .ZN(
        n637) );
  OAI222_X1 U445 ( .A1(n643), .A2(n644), .B1(n16829), .B2(n646), .C1(n647), 
        .C2(n648), .ZN(n636) );
  INV_X1 U446 ( .A(n535), .ZN(n647) );
  OAI21_X1 U447 ( .B1(n649), .B2(n514), .A(n650), .ZN(n535) );
  AOI221_X1 U448 ( .B1(n16861), .B2(n651), .C1(n16823), .C2(n16828), .A(n652), 
        .ZN(n643) );
  OAI33_X1 U449 ( .A1(n653), .A2(n16853), .A3(n16836), .B1(n654), .B2(n16810), 
        .B3(n655), .ZN(n652) );
  OAI222_X1 U450 ( .A1(n656), .A2(n552), .B1(n657), .B2(n610), .C1(n658), .C2(
        n576), .ZN(n635) );
  INV_X1 U451 ( .A(n577), .ZN(n658) );
  NAND3_X1 U452 ( .A1(n16800), .A2(n659), .A3(n16801), .ZN(n577) );
  AOI222_X1 U453 ( .A1(n660), .A2(n195), .B1(n609), .B2(n16836), .C1(n590), 
        .C2(n661), .ZN(n657) );
  OAI221_X1 U454 ( .B1(n662), .B2(n663), .C1(n664), .C2(n665), .A(n666), .ZN(
        n661) );
  NAND2_X1 U455 ( .A1(n667), .A2(n16850), .ZN(n665) );
  NAND2_X1 U456 ( .A1(n16680), .A2(n16834), .ZN(n663) );
  AOI222_X1 U457 ( .A1(n16796), .A2(n17098), .B1(n17099), .B2(n668), .C1(
        n16815), .C2(n669), .ZN(n656) );
  OR3_X1 U458 ( .A1(n670), .A2(n671), .A3(n672), .ZN(n634) );
  OAI33_X1 U459 ( .A1(n650), .A2(n4956), .A3(n16864), .B1(n514), .B2(n16845), 
        .B3(n673), .ZN(n672) );
  NOR4_X1 U460 ( .A1(n485), .A2(n674), .A3(n16808), .A4(n459), .ZN(n671) );
  NOR4_X1 U461 ( .A1(n676), .A2(n17098), .A3(n443), .A4(n677), .ZN(n670) );
  AOI21_X1 U462 ( .B1(n678), .B2(n504), .A(n679), .ZN(n676) );
  INV_X1 U463 ( .A(n680), .ZN(n678) );
  OAI221_X1 U464 ( .B1(n191), .B2(n324), .C1(n5255), .C2(n17101), .A(n681), 
        .ZN(n5776) );
  AOI21_X1 U465 ( .B1(n16738), .B2(vis_pc_o[0]), .A(n682), .ZN(n681) );
  NOR4_X1 U466 ( .A1(n683), .A2(n628), .A3(n684), .A4(n17103), .ZN(n682) );
  INV_X1 U467 ( .A(n638), .ZN(n628) );
  OAI221_X1 U469 ( .B1(n685), .B2(n17126), .C1(n16833), .C2(n17122), .A(n686), 
        .ZN(n5777) );
  NAND3_X1 U470 ( .A1(n529), .A2(n16851), .A3(n687), .ZN(n686) );
  NOR4_X1 U471 ( .A1(n688), .A2(n689), .A3(n690), .A4(n691), .ZN(n685) );
  OAI22_X1 U472 ( .A1(n692), .A2(n693), .B1(n5230), .B2(n694), .ZN(n691) );
  INV_X1 U473 ( .A(n695), .ZN(n693) );
  OAI33_X1 U474 ( .A1(n696), .A2(n5165), .A3(n605), .B1(n677), .B2(n697), .B3(
        n478), .ZN(n690) );
  OAI221_X1 U475 ( .B1(n698), .B2(n16808), .C1(n16864), .C2(n699), .A(n700), 
        .ZN(n689) );
  INV_X1 U476 ( .A(n701), .ZN(n700) );
  NOR4_X1 U477 ( .A1(n702), .A2(n703), .A3(n704), .A4(n705), .ZN(n698) );
  AOI21_X1 U478 ( .B1(n706), .B2(n707), .A(n16807), .ZN(n705) );
  NAND4_X1 U479 ( .A1(n485), .A2(n708), .A3(n709), .A4(n710), .ZN(n707) );
  NOR3_X1 U480 ( .A1(n659), .A2(n711), .A3(n712), .ZN(n710) );
  INV_X1 U481 ( .A(n444), .ZN(n485) );
  NAND3_X1 U482 ( .A1(n475), .A2(n16813), .A3(n629), .ZN(n706) );
  NOR3_X1 U483 ( .A1(n711), .A2(n580), .A3(n582), .ZN(n704) );
  OAI33_X1 U484 ( .A1(n713), .A2(n714), .A3(n715), .B1(n478), .B2(n716), .B3(
        n503), .ZN(n703) );
  AOI22_X1 U485 ( .A1(n16814), .A2(n717), .B1(n718), .B2(n679), .ZN(n716) );
  INV_X1 U486 ( .A(n719), .ZN(n717) );
  AOI211_X1 U487 ( .C1(n720), .C2(n721), .A(n16804), .B(n722), .ZN(n719) );
  OAI221_X1 U488 ( .B1(n556), .B2(n723), .C1(n724), .C2(n725), .A(n726), .ZN(
        n702) );
  AOI22_X1 U489 ( .A1(n727), .A2(n728), .B1(n729), .B2(n730), .ZN(n726) );
  AOI221_X1 U490 ( .B1(n731), .B2(n333), .C1(n732), .C2(n733), .A(n734), .ZN(
        n724) );
  INV_X1 U491 ( .A(n735), .ZN(n733) );
  AOI21_X1 U492 ( .B1(n16733), .B2(n505), .A(n736), .ZN(n735) );
  NAND4_X1 U493 ( .A1(n737), .A2(n738), .A3(n739), .A4(n740), .ZN(n688) );
  NOR4_X1 U494 ( .A1(n741), .A2(n742), .A3(n493), .A4(n545), .ZN(n740) );
  NOR3_X1 U495 ( .A1(n16828), .A2(n16836), .A3(n594), .ZN(n545) );
  NAND3_X1 U496 ( .A1(n16826), .A2(n16856), .A3(n744), .ZN(n739) );
  OAI21_X1 U497 ( .B1(n16820), .B2(n745), .A(n640), .ZN(n744) );
  NAND3_X1 U498 ( .A1(n16824), .A2(n16821), .A3(n746), .ZN(n737) );
  OAI22_X1 U499 ( .A1(n747), .A2(n17126), .B1(n17097), .B2(n748), .ZN(n5778)
         );
  AOI211_X1 U500 ( .C1(n16680), .C2(n16853), .A(n17126), .B(n534), .ZN(n748)
         );
  AOI211_X1 U501 ( .C1(n526), .C2(n16821), .A(n749), .B(n750), .ZN(n747) );
  OAI22_X1 U502 ( .A1(n499), .A2(n692), .B1(n751), .B2(n696), .ZN(n750) );
  OAI211_X1 U503 ( .C1(n752), .C2(n753), .A(n754), .B(n755), .ZN(n749) );
  OAI211_X1 U504 ( .C1(n756), .C2(n757), .A(n503), .B(n16802), .ZN(n754) );
  NOR2_X1 U505 ( .A1(n758), .A2(n759), .ZN(n756) );
  AOI21_X1 U506 ( .B1(n543), .B2(n760), .A(n761), .ZN(n752) );
  NOR3_X1 U507 ( .A1(n762), .A2(n16841), .A3(n16864), .ZN(n761) );
  OAI22_X1 U508 ( .A1(n764), .A2(n765), .B1(n5256), .B2(n766), .ZN(n5779) );
  AOI21_X1 U509 ( .B1(n767), .B2(n768), .A(n765), .ZN(n766) );
  AOI221_X1 U510 ( .B1(n769), .B2(n403), .C1(n770), .C2(n659), .A(n771), .ZN(
        n764) );
  OAI22_X1 U511 ( .A1(n16816), .A2(n772), .B1(n5243), .B2(n773), .ZN(n771) );
  OAI22_X1 U513 ( .A1(n774), .A2(n765), .B1(n16810), .B2(n775), .ZN(n5780) );
  AOI21_X1 U514 ( .B1(n767), .B2(n776), .A(n765), .ZN(n775) );
  NOR3_X1 U515 ( .A1(n777), .A2(n778), .A3(n779), .ZN(n774) );
  INV_X1 U516 ( .A(n780), .ZN(n779) );
  AOI22_X1 U517 ( .A1(n781), .A2(n770), .B1(n4806), .B2(n769), .ZN(n780) );
  AOI21_X1 U518 ( .B1(n782), .B2(n783), .A(n5034), .ZN(n769) );
  NOR2_X1 U519 ( .A1(n784), .A2(n785), .ZN(n783) );
  OAI33_X1 U520 ( .A1(n786), .A2(n16957), .A3(n788), .B1(n16659), .B2(n16815), 
        .B3(n790), .ZN(n778) );
  AOI21_X1 U521 ( .B1(n791), .B2(n466), .A(n792), .ZN(n790) );
  XNOR2_X1 U522 ( .A(n793), .B(n654), .ZN(n786) );
  NAND2_X1 U523 ( .A1(n794), .A2(n795), .ZN(n654) );
  NAND2_X1 U524 ( .A1(n17097), .A2(n16671), .ZN(n793) );
  OAI221_X1 U525 ( .B1(n16794), .B2(n773), .C1(n16796), .C2(n772), .A(n460), 
        .ZN(n777) );
  AOI21_X1 U526 ( .B1(n797), .B2(n798), .A(n799), .ZN(n460) );
  INV_X1 U527 ( .A(n800), .ZN(n773) );
  OAI22_X1 U528 ( .A1(n16851), .A2(n17122), .B1(n801), .B2(n17126), .ZN(n5781)
         );
  NOR2_X1 U529 ( .A1(n802), .A2(n803), .ZN(n801) );
  OAI211_X1 U530 ( .C1(n804), .C2(n16821), .A(n805), .B(n806), .ZN(n803) );
  AOI22_X1 U531 ( .A1(n807), .A2(n808), .B1(n809), .B2(n16826), .ZN(n806) );
  OAI21_X1 U532 ( .B1(n810), .B2(n811), .A(n16855), .ZN(n805) );
  OAI33_X1 U533 ( .A1(n514), .A2(n16828), .A3(n16841), .B1(n640), .B2(n812), 
        .B3(n16858), .ZN(n811) );
  AOI21_X1 U534 ( .B1(n5165), .B2(n16851), .A(n813), .ZN(n810) );
  NOR4_X1 U535 ( .A1(n814), .A2(n815), .A3(n816), .A4(n817), .ZN(n804) );
  OAI221_X1 U536 ( .B1(n499), .B2(n818), .C1(n819), .C2(n16813), .A(n820), 
        .ZN(n817) );
  AOI22_X1 U537 ( .A1(n821), .A2(n822), .B1(n629), .B2(n16659), .ZN(n820) );
  OAI211_X1 U538 ( .C1(n823), .C2(n16659), .A(n824), .B(n825), .ZN(n816) );
  AOI22_X1 U539 ( .A1(n826), .A2(n16871), .B1(n543), .B2(n827), .ZN(n825) );
  OAI211_X1 U540 ( .C1(n16802), .C2(n625), .A(n16680), .B(n828), .ZN(n826) );
  AOI221_X1 U541 ( .B1(n821), .B2(n829), .C1(n16811), .C2(n830), .A(n831), 
        .ZN(n828) );
  NOR3_X1 U542 ( .A1(n711), .A2(n16801), .A3(n832), .ZN(n831) );
  OAI22_X1 U543 ( .A1(n16803), .A2(n582), .B1(n833), .B2(n625), .ZN(n830) );
  NAND3_X1 U544 ( .A1(n833), .A2(n16657), .A3(n834), .ZN(n829) );
  OAI21_X1 U545 ( .B1(n835), .B2(n731), .A(n474), .ZN(n824) );
  NOR3_X1 U546 ( .A1(n16674), .A2(n16796), .A3(n16798), .ZN(n835) );
  AOI221_X1 U547 ( .B1(n474), .B2(n16683), .C1(n505), .C2(n791), .A(n684), 
        .ZN(n823) );
  INV_X1 U548 ( .A(n329), .ZN(n474) );
  OAI211_X1 U549 ( .C1(n838), .C2(n610), .A(n839), .B(n840), .ZN(n815) );
  AOI22_X1 U550 ( .A1(n841), .A2(n473), .B1(n842), .B2(n597), .ZN(n840) );
  AOI21_X1 U551 ( .B1(n16841), .B2(n606), .A(n16838), .ZN(n842) );
  AOI21_X1 U552 ( .B1(n843), .B2(n832), .A(n16814), .ZN(n841) );
  NAND3_X1 U553 ( .A1(n16815), .A2(n16686), .A3(n730), .ZN(n839) );
  AOI21_X1 U554 ( .B1(n844), .B2(n632), .A(n845), .ZN(n838) );
  NOR3_X1 U555 ( .A1(n846), .A2(n585), .A3(n617), .ZN(n845) );
  OR4_X1 U556 ( .A1(n847), .A2(n484), .A3(n482), .A4(n848), .ZN(n814) );
  NOR3_X1 U557 ( .A1(n849), .A2(n16871), .A3(n567), .ZN(n847) );
  OAI211_X1 U558 ( .C1(n850), .C2(n851), .A(n852), .B(n853), .ZN(n802) );
  NOR3_X1 U559 ( .A1(n854), .A2(n855), .A3(n856), .ZN(n853) );
  NOR3_X1 U560 ( .A1(n664), .A2(n715), .A3(n857), .ZN(n856) );
  NOR3_X1 U561 ( .A1(n650), .A2(n604), .A3(n849), .ZN(n854) );
  OAI21_X1 U562 ( .B1(n858), .B2(n807), .A(n16862), .ZN(n852) );
  NOR3_X1 U563 ( .A1(n859), .A2(n16819), .A3(n860), .ZN(n858) );
  AOI21_X1 U564 ( .B1(n597), .B2(n861), .A(n599), .ZN(n850) );
  NOR3_X1 U565 ( .A1(n16680), .A2(n16866), .A3(n16847), .ZN(n599) );
  OAI21_X1 U566 ( .B1(n16830), .B2(n16841), .A(n863), .ZN(n861) );
  OAI221_X1 U567 ( .B1(n5006), .B2(n16792), .C1(n4948), .C2(n324), .A(n865), 
        .ZN(n5782) );
  AOI22_X1 U568 ( .A1(n17104), .A2(haddr_o[31]), .B1(n866), .B2(n867), .ZN(
        n865) );
  INV_X1 U569 ( .A(n868), .ZN(n5783) );
  AOI221_X1 U570 ( .B1(haddr_o[9]), .B2(n17104), .C1(n869), .C2(n866), .A(n870), .ZN(n868) );
  OAI22_X1 U571 ( .A1(n16792), .A2(n4814), .B1(n324), .B2(n5546), .ZN(n870) );
  AOI22_X1 U573 ( .A1(n16738), .A2(vis_pc_o[2]), .B1(n322), .B2(vis_ipsr_o[3]), 
        .ZN(n872) );
  INV_X1 U574 ( .A(haddr_o[3]), .ZN(n871) );
  INV_X1 U575 ( .A(n873), .ZN(n5785) );
  AOI221_X1 U576 ( .B1(haddr_o[30]), .B2(n17104), .C1(n874), .C2(n866), .A(
        n875), .ZN(n873) );
  OAI22_X1 U577 ( .A1(n16793), .A2(n4817), .B1(n324), .B2(n4954), .ZN(n875) );
  AOI22_X1 U579 ( .A1(n16738), .A2(vis_pc_o[1]), .B1(n322), .B2(vis_ipsr_o[2]), 
        .ZN(n877) );
  OAI221_X1 U580 ( .B1(n878), .B2(n17103), .C1(n5626), .C2(n17101), .A(n879), 
        .ZN(n5787) );
  AOI22_X1 U581 ( .A1(n16738), .A2(vis_pc_o[27]), .B1(n322), .B2(vis_apsr_o[0]), .ZN(n879) );
  OAI221_X1 U583 ( .B1(n5239), .B2(n16793), .C1(n4953), .C2(n324), .A(n880), 
        .ZN(n5788) );
  AOI22_X1 U584 ( .A1(n17104), .A2(haddr_o[29]), .B1(n866), .B2(n881), .ZN(
        n880) );
  OAI221_X1 U585 ( .B1(n882), .B2(n17126), .C1(n16862), .C2(n17122), .A(n883), 
        .ZN(n5789) );
  NAND3_X1 U586 ( .A1(n4974), .A2(n592), .A3(n884), .ZN(n883) );
  NOR4_X1 U587 ( .A1(n885), .A2(n886), .A3(n887), .A4(n888), .ZN(n882) );
  OAI33_X1 U588 ( .A1(n653), .A2(n851), .A3(n532), .B1(n889), .B2(n16847), 
        .B3(n503), .ZN(n888) );
  NAND2_X1 U589 ( .A1(n631), .A2(n483), .ZN(n889) );
  NOR3_X1 U590 ( .A1(n650), .A2(n714), .A3(n715), .ZN(n887) );
  NAND4_X1 U591 ( .A1(n890), .A2(n618), .A3(n891), .A4(n892), .ZN(n886) );
  NAND3_X1 U592 ( .A1(n893), .A2(n894), .A3(n895), .ZN(n885) );
  AOI221_X1 U593 ( .B1(n809), .B2(n728), .C1(n649), .C2(n799), .A(n896), .ZN(
        n895) );
  AOI22_X1 U594 ( .A1(n897), .A2(n898), .B1(n899), .B2(n16864), .ZN(n894) );
  OAI21_X1 U595 ( .B1(n813), .B2(n900), .A(n522), .ZN(n899) );
  NAND2_X1 U596 ( .A1(n16838), .A2(n610), .ZN(n900) );
  OAI22_X1 U597 ( .A1(n762), .A2(n673), .B1(n846), .B2(n901), .ZN(n898) );
  NAND2_X1 U598 ( .A1(n632), .A2(n16856), .ZN(n901) );
  AOI22_X1 U599 ( .A1(n466), .A2(n902), .B1(n16819), .B2(n903), .ZN(n893) );
  NAND4_X1 U600 ( .A1(n904), .A2(n905), .A3(n906), .A4(n907), .ZN(n903) );
  NOR3_X1 U601 ( .A1(n908), .A2(n909), .A3(n910), .ZN(n907) );
  NOR3_X1 U602 ( .A1(n911), .A2(n715), .A3(n859), .ZN(n910) );
  OAI33_X1 U603 ( .A1(n694), .A2(n16853), .A3(n651), .B1(n912), .B2(n16832), 
        .B3(n16871), .ZN(n908) );
  AOI222_X1 U604 ( .A1(n708), .A2(n913), .B1(n914), .B2(n915), .C1(n597), .C2(
        n916), .ZN(n906) );
  OAI21_X1 U605 ( .B1(n917), .B2(n918), .A(n919), .ZN(n916) );
  OAI21_X1 U606 ( .B1(n714), .B2(n653), .A(n16867), .ZN(n915) );
  OAI22_X1 U607 ( .A1(n16795), .A2(n920), .B1(n16807), .B2(n921), .ZN(n913) );
  AOI22_X1 U608 ( .A1(n5243), .A2(n922), .B1(n923), .B2(n17098), .ZN(n921) );
  AOI221_X1 U609 ( .B1(n720), .B2(n16733), .C1(n721), .C2(n16815), .A(n924), 
        .ZN(n920) );
  XOR2_X1 U610 ( .A(n17098), .B(n731), .Z(n924) );
  AOI221_X1 U611 ( .B1(n4974), .B2(n925), .C1(n483), .C2(n926), .A(n927), .ZN(
        n905) );
  AOI21_X1 U612 ( .B1(n928), .B2(n16816), .A(n580), .ZN(n927) );
  XOR2_X1 U613 ( .A(n16798), .B(n16796), .Z(n928) );
  OAI211_X1 U614 ( .C1(n16847), .C2(n711), .A(n929), .B(n16854), .ZN(n926) );
  NAND3_X1 U615 ( .A1(n930), .A2(n596), .A3(n16862), .ZN(n929) );
  OAI221_X1 U616 ( .B1(n819), .B2(n931), .C1(n932), .C2(n582), .A(n933), .ZN(
        n925) );
  AOI21_X1 U617 ( .B1(n934), .B2(n935), .A(n494), .ZN(n933) );
  INV_X1 U618 ( .A(n627), .ZN(n494) );
  NAND2_X1 U619 ( .A1(n936), .A2(n16814), .ZN(n627) );
  OAI211_X1 U620 ( .C1(n16800), .C2(n16657), .A(n937), .B(n938), .ZN(n935) );
  AOI221_X1 U621 ( .B1(n721), .B2(n16815), .C1(n668), .C2(n16817), .A(n939), 
        .ZN(n938) );
  XOR2_X1 U622 ( .A(n17098), .B(n469), .Z(n937) );
  AOI222_X1 U623 ( .A1(n934), .A2(n16659), .B1(n684), .B2(n475), .C1(n16797), 
        .C2(n482), .ZN(n904) );
  INV_X1 U624 ( .A(n940), .ZN(n684) );
  NAND4_X1 U625 ( .A1(n941), .A2(n819), .A3(n512), .A4(n942), .ZN(n902) );
  AOI221_X1 U626 ( .B1(n822), .B2(n16683), .C1(n943), .C2(n16734), .A(n944), 
        .ZN(n942) );
  NOR3_X1 U627 ( .A1(n945), .A2(n16862), .A3(n16659), .ZN(n944) );
  OAI221_X1 U628 ( .B1(haddr_o[4]), .B2(n946), .C1(n5502), .C2(n17122), .A(
        n255), .ZN(n5790) );
  OAI221_X1 U629 ( .B1(n947), .B2(n946), .C1(n5149), .C2(n17122), .A(n255), 
        .ZN(n5791) );
  XOR2_X1 U630 ( .A(haddr_o[3]), .B(n948), .Z(n947) );
  OAI211_X1 U631 ( .C1(n5096), .C2(n17122), .A(n949), .B(n255), .ZN(n5792) );
  OAI21_X1 U632 ( .B1(haddr_o[5]), .B2(haddr_o[3]), .A(n256), .ZN(n949) );
  OAI221_X1 U633 ( .B1(haddr_o[8]), .B2(n946), .C1(n5017), .C2(n17122), .A(
        n255), .ZN(n5793) );
  OAI21_X1 U634 ( .B1(n950), .B2(n951), .A(n256), .ZN(n255) );
  NAND4_X1 U635 ( .A1(haddr_o[15]), .A2(n952), .A3(n953), .A4(n954), .ZN(n951)
         );
  NOR4_X1 U636 ( .A1(n955), .A2(n956), .A3(n957), .A4(n958), .ZN(n954) );
  AOI22_X1 U637 ( .A1(n959), .A2(n960), .B1(n961), .B2(n962), .ZN(n958) );
  NOR4_X1 U638 ( .A1(haddr_o[9]), .A2(haddr_o[7]), .A3(haddr_o[6]), .A4(
        haddr_o[5]), .ZN(n962) );
  AOI221_X1 U639 ( .B1(haddr_o[8]), .B2(n963), .C1(n964), .C2(haddr_o[11]), 
        .A(n965), .ZN(n961) );
  NOR3_X1 U640 ( .A1(haddr_o[10]), .A2(haddr_o[4]), .A3(haddr_o[3]), .ZN(n965)
         );
  NAND3_X1 U641 ( .A1(haddr_o[8]), .A2(haddr_o[2]), .A3(haddr_o[10]), .ZN(n964) );
  NOR3_X1 U642 ( .A1(n966), .A2(haddr_o[6]), .A3(haddr_o[3]), .ZN(n960) );
  AOI21_X1 U643 ( .B1(n876), .B2(n967), .A(n968), .ZN(n966) );
  AOI21_X1 U644 ( .B1(n969), .B2(n970), .A(n971), .ZN(n959) );
  XNOR2_X1 U645 ( .A(haddr_o[9]), .B(haddr_o[8]), .ZN(n971) );
  NAND4_X1 U646 ( .A1(n967), .A2(n968), .A3(n876), .A4(n972), .ZN(n970) );
  NOR2_X1 U647 ( .A1(haddr_o[10]), .A2(haddr_o[11]), .ZN(n972) );
  NOR3_X1 U649 ( .A1(haddr_o[16]), .A2(haddr_o[18]), .A3(haddr_o[17]), .ZN(
        n953) );
  NAND4_X1 U650 ( .A1(n973), .A2(n317), .A3(n974), .A4(n975), .ZN(n950) );
  NOR4_X1 U651 ( .A1(haddr_o[22]), .A2(haddr_o[21]), .A3(haddr_o[20]), .A4(
        haddr_o[19]), .ZN(n975) );
  NOR3_X1 U652 ( .A1(haddr_o[25]), .A2(haddr_o[27]), .A3(haddr_o[26]), .ZN(
        n974) );
  NAND2_X1 U653 ( .A1(n976), .A2(n977), .ZN(n5794) );
  NAND3_X1 U654 ( .A1(n978), .A2(n979), .A3(n980), .ZN(n977) );
  OAI21_X1 U655 ( .B1(n981), .B2(n16808), .A(n17127), .ZN(n976) );
  AOI21_X1 U656 ( .B1(n982), .B2(n983), .A(n984), .ZN(n981) );
  AOI211_X1 U657 ( .C1(n728), .C2(n985), .A(n986), .B(n987), .ZN(n983) );
  NOR3_X1 U658 ( .A1(n699), .A2(n16853), .A3(n16839), .ZN(n987) );
  INV_X1 U659 ( .A(n988), .ZN(n986) );
  OAI21_X1 U660 ( .B1(n989), .B2(n655), .A(n891), .ZN(n985) );
  AOI222_X1 U661 ( .A1(n990), .A2(n757), .B1(n991), .B2(n992), .C1(n993), .C2(
        n16864), .ZN(n982) );
  OAI22_X1 U662 ( .A1(n994), .A2(n558), .B1(n16848), .B2(n995), .ZN(n993) );
  OAI22_X1 U663 ( .A1(n16842), .A2(n624), .B1(n996), .B2(n616), .ZN(n992) );
  AOI222_X1 U664 ( .A1(n526), .A2(n997), .B1(n998), .B2(n16851), .C1(n563), 
        .C2(n16836), .ZN(n996) );
  OAI22_X1 U665 ( .A1(n5231), .A2(n17123), .B1(n17127), .B2(n999), .ZN(n5795)
         );
  OAI21_X1 U666 ( .B1(n430), .B2(n431), .A(n1000), .ZN(n5796) );
  NAND4_X1 U667 ( .A1(n430), .A2(n1001), .A3(n334), .A4(n1002), .ZN(n1000) );
  OAI21_X1 U668 ( .B1(n5233), .B2(n1003), .A(n1004), .ZN(n5797) );
  NAND2_X1 U669 ( .A1(n1005), .A2(n1006), .ZN(n5798) );
  OAI211_X1 U670 ( .C1(n189), .C2(n1007), .A(n1008), .B(n17124), .ZN(n1006) );
  OAI21_X1 U671 ( .B1(n189), .B2(n17111), .A(n1009), .ZN(n1005) );
  INV_X1 U672 ( .A(n37), .ZN(n42) );
  INV_X1 U673 ( .A(n1010), .ZN(n189) );
  OAI21_X1 U674 ( .B1(n5229), .B2(n1011), .A(n1012), .ZN(n5799) );
  NOR3_X1 U675 ( .A1(n200), .A2(n186), .A3(n181), .ZN(n1011) );
  OAI22_X1 U676 ( .A1(n4947), .A2(n17123), .B1(n1013), .B2(n17126), .ZN(n5800)
         );
  NOR4_X1 U677 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
  OAI33_X1 U678 ( .A1(n843), .A2(n1018), .A3(n552), .B1(n1019), .B2(n16795), 
        .B3(n1020), .ZN(n1017) );
  NOR2_X1 U679 ( .A1(n16812), .A2(n1021), .ZN(n1020) );
  AOI21_X1 U680 ( .B1(n1022), .B2(n16798), .A(n922), .ZN(n1018) );
  INV_X1 U681 ( .A(n712), .ZN(n922) );
  NOR3_X1 U682 ( .A1(n699), .A2(n16839), .A3(n1023), .ZN(n1016) );
  NAND3_X1 U683 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1015) );
  OAI211_X1 U684 ( .C1(n333), .C2(n465), .A(n16804), .B(n574), .ZN(n1026) );
  OAI211_X1 U685 ( .C1(n1027), .C2(n514), .A(n1028), .B(n1029), .ZN(n1014) );
  AOI222_X1 U686 ( .A1(n563), .A2(n1030), .B1(n991), .B2(n1031), .C1(n728), 
        .C2(n1032), .ZN(n1029) );
  OAI22_X1 U687 ( .A1(n16830), .A2(n650), .B1(n808), .B2(n1033), .ZN(n1032) );
  NAND2_X1 U688 ( .A1(n528), .A2(n1034), .ZN(n1033) );
  OAI21_X1 U689 ( .B1(n994), .B2(n1035), .A(n646), .ZN(n1031) );
  OAI221_X1 U690 ( .B1(n610), .B2(n699), .C1(n499), .C2(n692), .A(n1036), .ZN(
        n1030) );
  INV_X1 U691 ( .A(n1037), .ZN(n1036) );
  OAI22_X1 U692 ( .A1(n16820), .A2(n193), .B1(n422), .B2(n1038), .ZN(n5823) );
  OAI21_X1 U693 ( .B1(n1039), .B2(n1040), .A(n17125), .ZN(n1038) );
  NOR2_X1 U694 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
  AOI21_X1 U695 ( .B1(n1043), .B2(n641), .A(n196), .ZN(n193) );
  OAI22_X1 U696 ( .A1(n1044), .A2(n1045), .B1(n1046), .B2(n1047), .ZN(n5824)
         );
  INV_X1 U697 ( .A(n1048), .ZN(n1046) );
  INV_X1 U698 ( .A(n1047), .ZN(n1044) );
  NAND2_X1 U699 ( .A1(n17124), .A2(n1049), .ZN(n1047) );
  OAI21_X1 U700 ( .B1(n1050), .B2(n930), .A(n1051), .ZN(n5825) );
  OAI21_X1 U701 ( .B1(n1052), .B2(n200), .A(n1053), .ZN(n1051) );
  OAI21_X1 U702 ( .B1(n5234), .B2(n1054), .A(n1055), .ZN(n5826) );
  OAI211_X1 U703 ( .C1(n1056), .C2(n1057), .A(n16808), .B(n5167), .ZN(n1055)
         );
  NOR3_X1 U704 ( .A1(vis_pc_o[1]), .A2(n16806), .A3(n196), .ZN(n1057) );
  NAND2_X1 U705 ( .A1(n17124), .A2(n1058), .ZN(n196) );
  NOR4_X1 U706 ( .A1(n186), .A2(n181), .A3(n1059), .A4(n1058), .ZN(n1056) );
  OAI22_X1 U707 ( .A1(n1054), .A2(n184), .B1(n1059), .B2(n1060), .ZN(n5827) );
  OAI21_X1 U708 ( .B1(n1061), .B2(n1062), .A(n16808), .ZN(n1060) );
  NOR2_X1 U709 ( .A1(n5167), .A2(n5228), .ZN(n1062) );
  NOR3_X1 U710 ( .A1(n1063), .A2(n183), .A3(n1058), .ZN(n1061) );
  OAI22_X1 U712 ( .A1(n5230), .A2(n17123), .B1(n1064), .B2(n17126), .ZN(n5828)
         );
  AOI22_X1 U713 ( .A1(n1065), .A2(n181), .B1(n183), .B2(n1066), .ZN(n1064) );
  OAI21_X1 U714 ( .B1(n1067), .B2(n1068), .A(n5229), .ZN(n1065) );
  INV_X1 U715 ( .A(n1069), .ZN(n1068) );
  OAI22_X1 U716 ( .A1(n19), .A2(n1070), .B1(n4826), .B2(n1071), .ZN(n4854) );
  OAI22_X1 U717 ( .A1(n19), .A2(n16781), .B1(n5515), .B2(n17095), .ZN(n4855)
         );
  OAI22_X1 U718 ( .A1(n247), .A2(n17094), .B1(n5505), .B2(n17095), .ZN(n4856)
         );
  OAI22_X1 U719 ( .A1(n229), .A2(n17094), .B1(n5520), .B2(n17095), .ZN(n4857)
         );
  OAI22_X1 U720 ( .A1(n245), .A2(n16781), .B1(n5506), .B2(n17095), .ZN(n4858)
         );
  OAI22_X1 U721 ( .A1(n226), .A2(n16781), .B1(n5517), .B2(n17095), .ZN(n4859)
         );
  OAI22_X1 U722 ( .A1(n5516), .A2(n1074), .B1(n249), .B2(n1075), .ZN(n4860) );
  OAI22_X1 U723 ( .A1(n249), .A2(n17094), .B1(n5510), .B2(n17095), .ZN(n4861)
         );
  OAI22_X1 U724 ( .A1(n5503), .A2(n1076), .B1(n1077), .B2(n1078), .ZN(n4862)
         );
  OAI22_X1 U725 ( .A1(n5168), .A2(n1079), .B1(n221), .B2(n1080), .ZN(n4863) );
  OAI22_X1 U726 ( .A1(n4829), .A2(n1079), .B1(n215), .B2(n1080), .ZN(n4864) );
  OAI22_X1 U727 ( .A1(n240), .A2(n16781), .B1(n5507), .B2(n17095), .ZN(n4865)
         );
  OAI22_X1 U728 ( .A1(n236), .A2(n16781), .B1(n5508), .B2(n17095), .ZN(n4866)
         );
  OAI22_X1 U729 ( .A1(n221), .A2(n16781), .B1(n5509), .B2(n17095), .ZN(n4867)
         );
  OAI22_X1 U730 ( .A1(n210), .A2(n16781), .B1(n5511), .B2(n17095), .ZN(n4868)
         );
  OAI22_X1 U731 ( .A1(n215), .A2(n16781), .B1(n5512), .B2(n17095), .ZN(n4869)
         );
  OAI22_X1 U732 ( .A1(n218), .A2(n16781), .B1(n5513), .B2(n17095), .ZN(n4870)
         );
  OAI22_X1 U733 ( .A1(n224), .A2(n16781), .B1(n5514), .B2(n17095), .ZN(n4871)
         );
  OAI22_X1 U734 ( .A1(n238), .A2(n17094), .B1(n5571), .B2(n17095), .ZN(n4872)
         );
  OAI22_X1 U735 ( .A1(n242), .A2(n17094), .B1(n5600), .B2(n17095), .ZN(n4873)
         );
  OAI22_X1 U736 ( .A1(n4833), .A2(n1074), .B1(n210), .B2(n1075), .ZN(n4874) );
  INV_X1 U737 ( .A(n1074), .ZN(n1075) );
  NOR3_X1 U738 ( .A1(n251), .A2(n5007), .A3(n261), .ZN(n1074) );
  OAI21_X1 U739 ( .B1(n4834), .B2(n17123), .A(n1081), .ZN(n4875) );
  NAND4_X1 U740 ( .A1(n1082), .A2(n422), .A3(n1083), .A4(n1084), .ZN(n1081) );
  AOI221_X1 U741 ( .B1(n1085), .B2(n651), .C1(n1086), .C2(n1087), .A(n17126), 
        .ZN(n1084) );
  OAI22_X1 U743 ( .A1(n16854), .A2(n696), .B1(n1088), .B2(n16826), .ZN(n1085)
         );
  INV_X1 U744 ( .A(n1089), .ZN(n1083) );
  AOI21_X1 U745 ( .B1(n590), .B2(n1090), .A(n1091), .ZN(n1089) );
  AOI221_X1 U746 ( .B1(n16864), .B2(n1092), .C1(n1093), .C2(n1087), .A(n1094), 
        .ZN(n1091) );
  NAND3_X1 U747 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1082) );
  OAI22_X1 U748 ( .A1(n5829), .A2(n1059), .B1(n5165), .B2(n687), .ZN(n4876) );
  OAI21_X1 U749 ( .B1(n1098), .B2(n1099), .A(n194), .ZN(n5829) );
  NAND4_X1 U750 ( .A1(n7), .A2(n8), .A3(n9), .A4(n2), .ZN(n1099) );
  NAND4_X1 U755 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n1098) );
  OAI21_X1 U760 ( .B1(n4843), .B2(n17123), .A(n1100), .ZN(n4878) );
  OAI21_X1 U761 ( .B1(n1101), .B2(n1102), .A(n17125), .ZN(n1100) );
  NOR3_X1 U762 ( .A1(n1103), .A2(n16821), .A3(n1104), .ZN(n1102) );
  NOR4_X1 U763 ( .A1(n532), .A2(n556), .A3(n616), .A4(n568), .ZN(n1101) );
  OAI21_X1 U764 ( .B1(n4845), .B2(n17123), .A(n1105), .ZN(n4879) );
  OAI211_X1 U765 ( .C1(n1106), .C2(n1009), .A(n1107), .B(n17124), .ZN(n1105)
         );
  OAI22_X1 U766 ( .A1(n181), .A2(n1059), .B1(n5228), .B2(n687), .ZN(n4880) );
  OAI22_X1 U767 ( .A1(n373), .A2(n1108), .B1(n4847), .B2(n1109), .ZN(n4881) );
  OAI22_X1 U768 ( .A1(n4848), .A2(n1079), .B1(n210), .B2(n1080), .ZN(n4882) );
  INV_X1 U769 ( .A(n1080), .ZN(n1079) );
  NAND3_X1 U770 ( .A1(n1110), .A2(n253), .A3(n1111), .ZN(n1080) );
  OAI22_X1 U771 ( .A1(n1077), .A2(n1070), .B1(n5097), .B2(n1071), .ZN(n4883)
         );
  OAI22_X1 U772 ( .A1(n232), .A2(n17094), .B1(n5581), .B2(n17095), .ZN(n4884)
         );
  OAI22_X1 U773 ( .A1(n1112), .A2(n17094), .B1(n5639), .B2(n17095), .ZN(n4885)
         );
  OAI22_X1 U774 ( .A1(n5167), .A2(n17123), .B1(n1113), .B2(n17126), .ZN(n4886)
         );
  OAI22_X1 U775 ( .A1(n1114), .A2(n17094), .B1(n5033), .B2(n17095), .ZN(n4887)
         );
  OAI22_X1 U776 ( .A1(n1115), .A2(n17094), .B1(n5067), .B2(n17095), .ZN(n4888)
         );
  OAI22_X1 U777 ( .A1(n234), .A2(n17094), .B1(n5579), .B2(n17095), .ZN(n4889)
         );
  OAI22_X1 U778 ( .A1(n1116), .A2(n17094), .B1(n5625), .B2(n17095), .ZN(n4890)
         );
  OAI22_X1 U779 ( .A1(n1117), .A2(n17094), .B1(n5618), .B2(n17095), .ZN(n4891)
         );
  OAI22_X1 U780 ( .A1(n1118), .A2(n17094), .B1(n5074), .B2(n17095), .ZN(n4892)
         );
  AOI21_X1 U781 ( .B1(n17092), .B2(n1120), .A(n1121), .ZN(n4902) );
  AOI21_X1 U782 ( .B1(n17092), .B2(n1122), .A(n1123), .ZN(n4903) );
  AOI221_X1 U783 ( .B1(n1124), .B2(hwdata_o[9]), .C1(n1125), .C2(n1126), .A(
        n1127), .ZN(n4904) );
  OAI21_X1 U784 ( .B1(n1128), .B2(n1129), .A(irq_i[9]), .ZN(n1127) );
  OAI22_X1 U786 ( .A1(n4777), .A2(n1109), .B1(n1130), .B2(n1131), .ZN(n4906)
         );
  INV_X1 U787 ( .A(hrdata_i[16]), .ZN(n1130) );
  OAI22_X1 U788 ( .A1(n4778), .A2(n1109), .B1(n1132), .B2(n1131), .ZN(n4907)
         );
  INV_X1 U789 ( .A(hrdata_i[17]), .ZN(n1132) );
  OAI22_X1 U790 ( .A1(n4779), .A2(n1109), .B1(n1133), .B2(n1131), .ZN(n4908)
         );
  INV_X1 U791 ( .A(hrdata_i[18]), .ZN(n1133) );
  OAI22_X1 U792 ( .A1(n4780), .A2(n1109), .B1(n1134), .B2(n1131), .ZN(n4909)
         );
  INV_X1 U793 ( .A(hrdata_i[19]), .ZN(n1134) );
  OAI22_X1 U794 ( .A1(n4781), .A2(n1109), .B1(n1135), .B2(n1131), .ZN(n4910)
         );
  INV_X1 U795 ( .A(hrdata_i[20]), .ZN(n1135) );
  OAI22_X1 U796 ( .A1(n4782), .A2(n1109), .B1(n1136), .B2(n1131), .ZN(n4911)
         );
  INV_X1 U797 ( .A(hrdata_i[21]), .ZN(n1136) );
  OAI22_X1 U798 ( .A1(n4783), .A2(n1109), .B1(n1137), .B2(n1131), .ZN(n4912)
         );
  INV_X1 U799 ( .A(hrdata_i[22]), .ZN(n1137) );
  OAI22_X1 U800 ( .A1(n4784), .A2(n1109), .B1(n1138), .B2(n1131), .ZN(n4913)
         );
  INV_X1 U801 ( .A(hrdata_i[23]), .ZN(n1138) );
  OAI22_X1 U802 ( .A1(n4785), .A2(n1109), .B1(n1139), .B2(n1131), .ZN(n4914)
         );
  INV_X1 U803 ( .A(hrdata_i[24]), .ZN(n1139) );
  OAI22_X1 U804 ( .A1(n4786), .A2(n1109), .B1(n1140), .B2(n1131), .ZN(n4915)
         );
  OAI22_X1 U805 ( .A1(n4787), .A2(n1109), .B1(n1141), .B2(n1131), .ZN(n4916)
         );
  INV_X1 U806 ( .A(hrdata_i[26]), .ZN(n1141) );
  OAI22_X1 U807 ( .A1(n4788), .A2(n1109), .B1(n1142), .B2(n1131), .ZN(n4917)
         );
  OAI22_X1 U808 ( .A1(n4789), .A2(n1109), .B1(n1143), .B2(n1131), .ZN(n4918)
         );
  OAI22_X1 U809 ( .A1(n4790), .A2(n1109), .B1(n1144), .B2(n1131), .ZN(n4919)
         );
  OAI22_X1 U810 ( .A1(n4791), .A2(n1109), .B1(n1145), .B2(n1131), .ZN(n4920)
         );
  OAI22_X1 U811 ( .A1(n4792), .A2(n1109), .B1(n1146), .B2(n1131), .ZN(n4921)
         );
  INV_X1 U813 ( .A(hrdata_i[31]), .ZN(n1146) );
  OAI222_X1 U816 ( .A1(n1149), .A2(n17103), .B1(n4820), .B2(n16793), .C1(n4762), .C2(n17101), .ZN(n4925) );
  INV_X1 U818 ( .A(n1151), .ZN(n4927) );
  AOI222_X1 U819 ( .A1(haddr_o[6]), .A2(n17104), .B1(vis_pc_o[5]), .B2(n16738), 
        .C1(n1152), .C2(n866), .ZN(n1151) );
  OAI222_X1 U821 ( .A1(n1153), .A2(n318), .B1(n5238), .B2(n16793), .C1(n4764), 
        .C2(n17100), .ZN(n4928) );
  OAI222_X1 U822 ( .A1(n1154), .A2(n318), .B1(n5573), .B2(n16792), .C1(n4765), 
        .C2(n17101), .ZN(n4929) );
  OAI222_X1 U823 ( .A1(n1155), .A2(n318), .B1(n5601), .B2(n16793), .C1(n4766), 
        .C2(n17101), .ZN(n4930) );
  OAI222_X1 U824 ( .A1(n1156), .A2(n318), .B1(n5114), .B2(n16793), .C1(n4767), 
        .C2(n17101), .ZN(n4931) );
  INV_X1 U825 ( .A(haddr_o[19]), .ZN(n1156) );
  OAI222_X1 U826 ( .A1(n1157), .A2(n318), .B1(n5237), .B2(n16792), .C1(n4768), 
        .C2(n17100), .ZN(n4932) );
  OAI222_X1 U827 ( .A1(n1158), .A2(n318), .B1(n5236), .B2(n16792), .C1(n4769), 
        .C2(n17100), .ZN(n4933) );
  OAI222_X1 U828 ( .A1(n1159), .A2(n318), .B1(n5235), .B2(n16793), .C1(n4770), 
        .C2(n17100), .ZN(n4934) );
  OAI222_X1 U831 ( .A1(n952), .A2(n318), .B1(n4812), .B2(n16793), .C1(n4830), 
        .C2(n17100), .ZN(n4937) );
  INV_X1 U833 ( .A(haddr_o[11]), .ZN(n963) );
  OAI222_X1 U834 ( .A1(n948), .A2(n17103), .B1(n4811), .B2(n16793), .C1(n4771), 
        .C2(n17100), .ZN(n4939) );
  INV_X1 U835 ( .A(n1160), .ZN(n4940) );
  AOI222_X1 U836 ( .A1(haddr_o[8]), .A2(n17104), .B1(vis_pc_o[7]), .B2(n16738), 
        .C1(n1161), .C2(n866), .ZN(n1160) );
  INV_X1 U838 ( .A(n1162), .ZN(n4941) );
  AOI222_X1 U839 ( .A1(haddr_o[15]), .A2(n17104), .B1(vis_pc_o[14]), .B2(
        n16738), .C1(n1163), .C2(n866), .ZN(n1162) );
  AOI22_X1 U844 ( .A1(n16738), .A2(vis_pc_o[4]), .B1(n322), .B2(vis_ipsr_o[5]), 
        .ZN(n1164) );
  AOI22_X1 U847 ( .A1(n16738), .A2(vis_pc_o[3]), .B1(n322), .B2(vis_ipsr_o[4]), 
        .ZN(n1165) );
  INV_X1 U848 ( .A(n324), .ZN(n322) );
  NAND2_X1 U849 ( .A1(n784), .A2(n17102), .ZN(n324) );
  NAND2_X1 U853 ( .A1(n17102), .A2(n1166), .ZN(n318) );
  OAI211_X1 U854 ( .C1(n16841), .C2(n692), .A(n1167), .B(n762), .ZN(n1166) );
  OAI21_X1 U855 ( .B1(n16659), .B2(n931), .A(n17097), .ZN(n1167) );
  AOI222_X1 U859 ( .A1(n1172), .A2(n1173), .B1(n1174), .B2(n16851), .C1(n16819), .C2(n1175), .ZN(n1171) );
  OAI221_X1 U860 ( .B1(n16811), .B2(n1176), .C1(n846), .C2(n1027), .A(n1177), 
        .ZN(n1175) );
  OAI211_X1 U861 ( .C1(n16839), .C2(n1178), .A(n1179), .B(n1180), .ZN(n1168)
         );
  NOR3_X1 U862 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
  AOI211_X1 U863 ( .C1(n679), .C2(n548), .A(n479), .B(n478), .ZN(n1183) );
  NOR3_X1 U864 ( .A1(n580), .A2(n16795), .A3(n1184), .ZN(n1181) );
  NAND3_X1 U865 ( .A1(n16854), .A2(n16848), .A3(n506), .ZN(n1179) );
  OAI22_X1 U866 ( .A1(n4846), .A2(n1185), .B1(hprot_o[3]), .B2(n1186), .ZN(
        n4945) );
  INV_X1 U867 ( .A(n1185), .ZN(n1186) );
  NOR2_X1 U868 ( .A1(n999), .A2(n17127), .ZN(n1185) );
  OAI21_X1 U869 ( .B1(n17127), .B2(n200), .A(n194), .ZN(n5649) );
  INV_X1 U870 ( .A(n422), .ZN(n5648) );
  OAI22_X1 U871 ( .A1(n5504), .A2(n1076), .B1(n1078), .B2(n1187), .ZN(n5650)
         );
  INV_X1 U872 ( .A(n1078), .ZN(n1076) );
  NAND3_X1 U873 ( .A1(n1188), .A2(n253), .A3(n1189), .ZN(n1078) );
  OAI22_X1 U874 ( .A1(n1070), .A2(n1187), .B1(n5098), .B2(n1071), .ZN(n5651)
         );
  OAI22_X1 U875 ( .A1(n1190), .A2(n1070), .B1(n4961), .B2(n1071), .ZN(n5652)
         );
  INV_X1 U876 ( .A(n1070), .ZN(n1071) );
  NAND2_X1 U877 ( .A1(n1191), .A2(n253), .ZN(n1070) );
  OAI22_X1 U878 ( .A1(n1190), .A2(n17094), .B1(n17095), .B2(n262), .ZN(n5653)
         );
  AOI21_X1 U881 ( .B1(n16837), .B2(n17127), .A(n1192), .ZN(n9972) );
  NOR4_X1 U882 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
  OAI221_X1 U883 ( .B1(n1197), .B2(n1198), .C1(n16856), .C2(n988), .A(n1199), 
        .ZN(n1196) );
  AOI21_X1 U884 ( .B1(n1200), .B2(n16820), .A(n1201), .ZN(n1199) );
  AOI22_X1 U885 ( .A1(n1202), .A2(n1203), .B1(n630), .B2(n469), .ZN(n1197) );
  OAI211_X1 U886 ( .C1(n16814), .C2(n16674), .A(n669), .B(n17099), .ZN(n1203)
         );
  OAI221_X1 U887 ( .B1(n16803), .B2(n1204), .C1(n1205), .C2(n1087), .A(n1206), 
        .ZN(n1195) );
  AOI221_X1 U888 ( .B1(n844), .B2(n1207), .C1(n714), .C2(n1208), .A(n1209), 
        .ZN(n1206) );
  NOR3_X1 U889 ( .A1(n1210), .A2(n16871), .A3(n16864), .ZN(n1209) );
  OAI22_X1 U890 ( .A1(n818), .A2(n1211), .B1(n846), .B2(n1212), .ZN(n1208) );
  NAND2_X1 U891 ( .A1(n1213), .A2(n16862), .ZN(n1212) );
  INV_X1 U892 ( .A(n1214), .ZN(n844) );
  OR2_X1 U893 ( .A1(n1092), .A2(n16854), .ZN(n1087) );
  AOI222_X1 U894 ( .A1(n550), .A2(n732), .B1(n1215), .B2(n630), .C1(n1216), 
        .C2(n708), .ZN(n1204) );
  NOR2_X1 U895 ( .A1(n16869), .A2(n16686), .ZN(n1215) );
  OAI221_X1 U896 ( .B1(n797), .B2(n1217), .C1(n1218), .C2(n945), .A(n1219), 
        .ZN(n1194) );
  AOI22_X1 U897 ( .A1(n1220), .A2(n16813), .B1(n16814), .B2(n482), .ZN(n1219)
         );
  OAI221_X1 U898 ( .B1(n1221), .B2(n713), .C1(n1222), .C2(n16659), .A(n1223), 
        .ZN(n1193) );
  AOI222_X1 U899 ( .A1(n597), .A2(n1224), .B1(n914), .B2(n1225), .C1(n821), 
        .C2(n1226), .ZN(n1223) );
  OAI21_X1 U900 ( .B1(n1227), .B2(n1228), .A(n941), .ZN(n1226) );
  NOR3_X1 U901 ( .A1(n1229), .A2(n5244), .A3(n16799), .ZN(n1227) );
  OAI21_X1 U902 ( .B1(n16674), .B2(n781), .A(n16815), .ZN(n1229) );
  OAI21_X1 U903 ( .B1(n649), .B2(n1230), .A(n1231), .ZN(n1225) );
  NAND4_X1 U904 ( .A1(n1232), .A2(n610), .A3(n16839), .A4(n16867), .ZN(n1231)
         );
  NAND2_X1 U905 ( .A1(n994), .A2(n1043), .ZN(n1232) );
  OAI222_X1 U906 ( .A1(n585), .A2(n1233), .B1(n16837), .B2(n1234), .C1(n16829), 
        .C2(n617), .ZN(n1224) );
  AOI221_X1 U907 ( .B1(n473), .B2(n16803), .C1(n333), .C2(n16817), .A(n1235), 
        .ZN(n1222) );
  OAI221_X1 U908 ( .B1(n1236), .B2(n941), .C1(n16813), .C2(n638), .A(n1237), 
        .ZN(n1235) );
  NAND3_X1 U909 ( .A1(n469), .A2(n16871), .A3(n1202), .ZN(n1237) );
  INV_X1 U910 ( .A(n711), .ZN(n1202) );
  NAND2_X1 U911 ( .A1(n16803), .A2(n16871), .ZN(n638) );
  AOI221_X1 U912 ( .B1(n16796), .B2(n1238), .C1(n16801), .C2(n16657), .A(n1239), .ZN(n1236) );
  OR2_X1 U913 ( .A1(n833), .A2(n718), .ZN(n1239) );
  AOI221_X1 U914 ( .B1(n526), .B2(n664), .C1(n16845), .C2(n16839), .A(n1240), 
        .ZN(n1221) );
  OAI21_X1 U915 ( .B1(n1104), .B2(n16839), .A(n567), .ZN(n1240) );
  NAND2_X1 U916 ( .A1(n16845), .A2(n753), .ZN(n567) );
  AOI22_X1 U917 ( .A1(n1241), .A2(n1242), .B1(n16823), .B2(n17126), .ZN(n9796)
         );
  NOR4_X1 U918 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1242) );
  OAI33_X1 U919 ( .A1(n552), .A2(n16804), .A3(n1247), .B1(n677), .B2(n1248), 
        .B3(n16821), .ZN(n1246) );
  AOI21_X1 U920 ( .B1(n1249), .B2(n473), .A(n734), .ZN(n1248) );
  INV_X1 U921 ( .A(n1176), .ZN(n734) );
  NAND2_X1 U922 ( .A1(n934), .A2(n16683), .ZN(n1176) );
  NOR2_X1 U923 ( .A1(n931), .A2(n16686), .ZN(n1249) );
  NOR3_X1 U924 ( .A1(n1250), .A2(n1251), .A3(n720), .ZN(n1247) );
  INV_X1 U925 ( .A(n547), .ZN(n1251) );
  NAND3_X1 U926 ( .A1(n16799), .A2(n17098), .A3(n731), .ZN(n547) );
  OAI33_X1 U927 ( .A1(n668), .A2(n17098), .A3(n16657), .B1(n16687), .B2(n16800), .B3(n718), .ZN(n1250) );
  NAND3_X1 U928 ( .A1(n934), .A2(n16807), .A3(n574), .ZN(n552) );
  OAI33_X1 U929 ( .A1(n580), .A2(n1252), .A3(n616), .B1(n569), .B2(n579), .B3(
        n723), .ZN(n1245) );
  AOI21_X1 U930 ( .B1(n16725), .B2(n16802), .A(n1253), .ZN(n1252) );
  NOR3_X1 U931 ( .A1(n583), .A2(n16807), .A3(n16796), .ZN(n1253) );
  OAI33_X1 U932 ( .A1(n1254), .A2(n851), .A3(n759), .B1(n1255), .B2(n576), 
        .B3(n659), .ZN(n1244) );
  NAND3_X1 U933 ( .A1(n709), .A2(n540), .A3(n1256), .ZN(n576) );
  NOR3_X1 U934 ( .A1(n443), .A2(n16797), .A3(n444), .ZN(n1256) );
  OAI21_X1 U935 ( .B1(n16801), .B2(n5243), .A(n16799), .ZN(n1255) );
  OAI211_X1 U936 ( .C1(n1257), .C2(n16808), .A(n1258), .B(n1259), .ZN(n1243)
         );
  NAND4_X1 U937 ( .A1(n574), .A2(n16804), .A3(n1260), .A4(n16813), .ZN(n1259)
         );
  OAI21_X1 U938 ( .B1(n1261), .B2(n843), .A(n478), .ZN(n1260) );
  INV_X1 U939 ( .A(n639), .ZN(n574) );
  NAND2_X1 U940 ( .A1(n475), .A2(n1262), .ZN(n639) );
  INV_X1 U941 ( .A(n1263), .ZN(n1258) );
  AOI211_X1 U942 ( .C1(n1264), .C2(n1265), .A(n1266), .B(n1182), .ZN(n1257) );
  NOR2_X1 U943 ( .A1(n459), .A2(n731), .ZN(n1182) );
  OAI22_X1 U944 ( .A1(n16797), .A2(n459), .B1(n16825), .B2(n640), .ZN(n1266)
         );
  NAND2_X1 U945 ( .A1(n631), .A2(n482), .ZN(n459) );
  NOR2_X1 U946 ( .A1(n16813), .A2(n1267), .ZN(n1264) );
  NOR4_X1 U947 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1241) );
  INV_X1 U948 ( .A(n1028), .ZN(n1270) );
  AOI221_X1 U949 ( .B1(n16862), .B2(n1174), .C1(n528), .C2(n534), .A(n1272), 
        .ZN(n1028) );
  INV_X1 U950 ( .A(n857), .ZN(n1174) );
  OAI21_X1 U951 ( .B1(n1273), .B2(n610), .A(n642), .ZN(n1269) );
  AOI221_X1 U952 ( .B1(n695), .B2(n612), .C1(n1021), .C2(n572), .A(n1274), 
        .ZN(n642) );
  NOR3_X1 U953 ( .A1(n443), .A2(n16725), .A3(n677), .ZN(n1274) );
  INV_X1 U954 ( .A(n1019), .ZN(n572) );
  NAND4_X1 U955 ( .A1(n540), .A2(n476), .A3(n505), .A4(n16797), .ZN(n1019) );
  AOI211_X1 U956 ( .C1(n660), .C2(n1275), .A(n1276), .B(n1277), .ZN(n1273) );
  NOR3_X1 U957 ( .A1(n1027), .A2(n16821), .A3(n846), .ZN(n1277) );
  NOR4_X1 U958 ( .A1(n16828), .A2(n650), .A3(n912), .A4(n664), .ZN(n1276) );
  OAI21_X1 U959 ( .B1(n16839), .B2(n860), .A(n607), .ZN(n1275) );
  OAI221_X1 U960 ( .B1(n1278), .B2(n644), .C1(n605), .C2(n1279), .A(n1280), 
        .ZN(n1268) );
  AOI22_X1 U961 ( .A1(n751), .A2(n1281), .B1(n827), .B2(n1282), .ZN(n1280) );
  OAI22_X1 U962 ( .A1(n16825), .A2(n692), .B1(n16854), .B2(n1035), .ZN(n1282)
         );
  NAND2_X1 U963 ( .A1(n699), .A2(n644), .ZN(n1281) );
  OAI22_X1 U964 ( .A1(n5257), .A2(n1283), .B1(n1284), .B2(n765), .ZN(n8706) );
  AOI22_X1 U965 ( .A1(n770), .A2(n16674), .B1(n800), .B2(n659), .ZN(n1284) );
  NAND2_X1 U966 ( .A1(n1285), .A2(n443), .ZN(n770) );
  AOI21_X1 U967 ( .B1(n767), .B2(n1286), .A(n765), .ZN(n1283) );
  OAI22_X1 U968 ( .A1(n5258), .A2(n1287), .B1(n1288), .B2(n765), .ZN(n8698) );
  AOI22_X1 U969 ( .A1(n1289), .A2(n16798), .B1(n800), .B2(n16674), .ZN(n1288)
         );
  OAI21_X1 U970 ( .B1(n819), .B2(n1184), .A(n892), .ZN(n800) );
  OAI21_X1 U971 ( .B1(n16816), .B2(n443), .A(n1285), .ZN(n1289) );
  INV_X1 U972 ( .A(n1290), .ZN(n1285) );
  OAI211_X1 U973 ( .C1(n16821), .C2(n945), .A(n1291), .B(n1292), .ZN(n1290) );
  AOI21_X1 U974 ( .B1(n541), .B2(n631), .A(n1293), .ZN(n1292) );
  INV_X1 U975 ( .A(n468), .ZN(n1293) );
  NAND2_X1 U976 ( .A1(n1220), .A2(n631), .ZN(n468) );
  AOI21_X1 U977 ( .B1(n767), .B2(n1294), .A(n765), .ZN(n1287) );
  OAI21_X1 U978 ( .B1(n1295), .B2(n1296), .A(n17125), .ZN(n765) );
  OAI211_X1 U979 ( .C1(n16683), .C2(n1297), .A(n489), .B(n1298), .ZN(n1296) );
  INV_X1 U980 ( .A(n1299), .ZN(n1298) );
  AOI221_X1 U981 ( .B1(n1300), .B2(n543), .C1(n914), .C2(n1301), .A(n1302), 
        .ZN(n489) );
  INV_X1 U982 ( .A(n1303), .ZN(n1301) );
  OAI221_X1 U983 ( .B1(n696), .B2(n1304), .C1(n498), .C2(n673), .A(n1305), 
        .ZN(n1295) );
  AOI22_X1 U984 ( .A1(n1306), .A2(n195), .B1(n809), .B2(n990), .ZN(n1305) );
  NAND2_X1 U985 ( .A1(n1042), .A2(n808), .ZN(n1304) );
  OAI211_X1 U986 ( .C1(n851), .C2(n1307), .A(n1308), .B(n1309), .ZN(n767) );
  AOI221_X1 U988 ( .B1(n1314), .B2(n249), .C1(n1315), .C2(n1316), .A(n1317), 
        .ZN(n1313) );
  INV_X1 U989 ( .A(irq_i[0]), .ZN(n1312) );
  NAND2_X1 U990 ( .A1(n17093), .A2(n1318), .ZN(n1311) );
  OAI221_X1 U991 ( .B1(n373), .B2(n430), .C1(n379), .C2(n1319), .A(n400), .ZN(
        n14934) );
  INV_X1 U992 ( .A(n379), .ZN(n430) );
  OAI211_X1 U993 ( .C1(n4847), .C2(n378), .A(n1320), .B(n1321), .ZN(n14928) );
  INV_X1 U994 ( .A(n1322), .ZN(n1321) );
  OAI22_X1 U995 ( .A1(n1319), .A2(n334), .B1(n336), .B2(n4974), .ZN(n1322) );
  NAND3_X1 U998 ( .A1(n377), .A2(n375), .A3(n336), .ZN(n1320) );
  NAND3_X1 U999 ( .A1(n5231), .A2(n1323), .A3(n336), .ZN(n378) );
  OAI211_X1 U1001 ( .C1(n1054), .C2(n1324), .A(n1107), .B(n1325), .ZN(n376) );
  INV_X1 U1002 ( .A(n1326), .ZN(n1107) );
  NOR3_X1 U1003 ( .A1(n1108), .A2(n1327), .A3(n1106), .ZN(n1324) );
  NOR2_X1 U1004 ( .A1(n17126), .A2(n16869), .ZN(n1054) );
  OAI21_X1 U1005 ( .B1(n4973), .B2(n1002), .A(n1001), .ZN(n1323) );
  OAI221_X1 U1007 ( .B1(n1328), .B2(n1329), .C1(n1330), .C2(n1331), .A(n1332), 
        .ZN(n14825) );
  NAND3_X1 U1008 ( .A1(n1331), .A2(vis_tbit_o), .A3(n1329), .ZN(n1332) );
  NAND4_X1 U1009 ( .A1(n37), .A2(n1333), .A3(n1010), .A4(n185), .ZN(n1331) );
  NAND2_X1 U1010 ( .A1(n187), .A2(n188), .ZN(n1010) );
  OAI211_X1 U1011 ( .C1(n16847), .C2(n797), .A(n1334), .B(n1335), .ZN(n1333)
         );
  AOI22_X1 U1012 ( .A1(n16829), .A2(n16842), .B1(n16836), .B2(n16856), .ZN(
        n1335) );
  INV_X1 U1014 ( .A(n1336), .ZN(n1330) );
  NAND2_X1 U1015 ( .A1(n86), .A2(n17124), .ZN(n1329) );
  NOR2_X1 U1016 ( .A1(n1336), .A2(n1337), .ZN(n1328) );
  OAI22_X1 U1017 ( .A1(n187), .A2(n16785), .B1(n192), .B2(n188), .ZN(n1336) );
  OAI211_X1 U1018 ( .C1(n370), .C2(n379), .A(n1339), .B(n400), .ZN(n14432) );
  NAND3_X1 U1019 ( .A1(hrdata_i[15]), .A2(n379), .A3(n373), .ZN(n1339) );
  INV_X1 U1020 ( .A(n377), .ZN(n373) );
  NAND3_X1 U1021 ( .A1(n984), .A2(vis_tbit_o), .A3(n4846), .ZN(n377) );
  INV_X1 U1023 ( .A(hresp_i), .ZN(n984) );
  NAND4_X1 U1025 ( .A1(n1109), .A2(n1327), .A3(n1001), .A4(n16868), .ZN(n1340)
         );
  INV_X1 U1026 ( .A(n1003), .ZN(n1327) );
  NAND2_X1 U1028 ( .A1(n17124), .A2(n375), .ZN(n1108) );
  INV_X1 U1029 ( .A(n431), .ZN(n400) );
  NAND2_X1 U1030 ( .A1(n5034), .A2(n422), .ZN(n431) );
  AOI21_X1 U1032 ( .B1(n5229), .B2(n1342), .A(n1343), .ZN(n1341) );
  NAND3_X1 U1033 ( .A1(n1069), .A2(n1344), .A3(n1345), .ZN(n1342) );
  AOI22_X1 U1034 ( .A1(n1048), .A2(n1049), .B1(vis_primask_o), .B2(n1346), 
        .ZN(n1345) );
  INV_X1 U1035 ( .A(n1049), .ZN(n1346) );
  OAI33_X1 U1036 ( .A1(n16656), .A2(n16810), .A3(n1348), .B1(n1349), .B2(
        n16823), .B3(n1350), .ZN(n1049) );
  NAND2_X1 U1037 ( .A1(n897), .A2(n751), .ZN(n1349) );
  OAI21_X1 U1038 ( .B1(n1351), .B2(n1348), .A(n1352), .ZN(n1048) );
  NAND3_X1 U1039 ( .A1(n751), .A2(n1353), .A3(n897), .ZN(n1352) );
  INV_X1 U1040 ( .A(n1354), .ZN(n1351) );
  INV_X1 U1041 ( .A(n1067), .ZN(n1344) );
  OAI211_X1 U1042 ( .C1(n1355), .C2(n1356), .A(n1357), .B(n1358), .ZN(n1069)
         );
  OAI21_X1 U1043 ( .B1(n1359), .B2(n1360), .A(n1361), .ZN(n1357) );
  NAND4_X1 U1044 ( .A1(n1362), .A2(n1363), .A3(n1364), .A4(n1365), .ZN(n1361)
         );
  INV_X1 U1045 ( .A(n1366), .ZN(n1364) );
  OAI21_X1 U1046 ( .B1(n1052), .B2(n5503), .A(n1367), .ZN(n1366) );
  AOI211_X1 U1047 ( .C1(n1355), .C2(n1368), .A(n1369), .B(n1370), .ZN(n1360)
         );
  AOI211_X1 U1048 ( .C1(n1355), .C2(n1371), .A(n1372), .B(n1373), .ZN(n1359)
         );
  INV_X1 U1049 ( .A(n1374), .ZN(n1356) );
  OAI22_X1 U1050 ( .A1(n1372), .A2(n1371), .B1(n1368), .B2(n1370), .ZN(n1374)
         );
  NOR3_X1 U1052 ( .A1(n1375), .A2(n1376), .A3(n1377), .ZN(n14001) );
  AOI21_X1 U1053 ( .B1(n17092), .B2(n1378), .A(n1379), .ZN(n1377) );
  AOI211_X1 U1055 ( .C1(n1314), .C2(n247), .A(n1317), .B(n1380), .ZN(n1376) );
  AOI21_X1 U1056 ( .B1(hwdata_o[15]), .B2(n1124), .A(n1378), .ZN(n1380) );
  INV_X1 U1057 ( .A(irq_i[15]), .ZN(n1375) );
  INV_X1 U1059 ( .A(irq_i[13]), .ZN(n1383) );
  OAI22_X1 U1060 ( .A1(n1384), .A2(n1314), .B1(n242), .B2(n1385), .ZN(n1382)
         );
  NAND2_X1 U1061 ( .A1(n17093), .A2(n1386), .ZN(n1381) );
  AOI221_X1 U1063 ( .B1(n1314), .B2(n218), .C1(n1390), .C2(n1391), .A(n1317), 
        .ZN(n1389) );
  INV_X1 U1064 ( .A(irq_i[3]), .ZN(n1388) );
  NAND2_X1 U1065 ( .A1(n17093), .A2(n1392), .ZN(n1387) );
  AOI221_X1 U1067 ( .B1(n1314), .B2(n215), .C1(n1396), .C2(n1397), .A(n1317), 
        .ZN(n1395) );
  INV_X1 U1068 ( .A(irq_i[2]), .ZN(n1394) );
  NAND2_X1 U1069 ( .A1(n17093), .A2(n1398), .ZN(n1393) );
  AOI221_X1 U1071 ( .B1(n1314), .B2(n229), .C1(n1402), .C2(n1403), .A(n1317), 
        .ZN(n1401) );
  INV_X1 U1072 ( .A(irq_i[7]), .ZN(n1400) );
  NAND2_X1 U1073 ( .A1(n17093), .A2(n1404), .ZN(n1399) );
  AOI221_X1 U1075 ( .B1(n1314), .B2(n226), .C1(n1408), .C2(n1409), .A(n1317), 
        .ZN(n1407) );
  INV_X1 U1076 ( .A(irq_i[6]), .ZN(n1406) );
  NAND2_X1 U1077 ( .A1(n17093), .A2(n1410), .ZN(n1405) );
  AOI221_X1 U1079 ( .B1(n1314), .B2(n224), .C1(n1415), .C2(n1416), .A(n1317), 
        .ZN(n1414) );
  INV_X1 U1080 ( .A(irq_i[5]), .ZN(n1413) );
  NAND2_X1 U1081 ( .A1(n17093), .A2(n1419), .ZN(n1412) );
  AOI221_X1 U1083 ( .B1(n221), .B2(n1314), .C1(n1423), .C2(n1424), .A(n1317), 
        .ZN(n1422) );
  INV_X1 U1084 ( .A(irq_i[4]), .ZN(n1421) );
  NAND2_X1 U1085 ( .A1(n17093), .A2(n1425), .ZN(n1420) );
  OAI21_X1 U1087 ( .B1(n183), .B2(n1314), .A(nmi_i), .ZN(n1427) );
  INV_X1 U1088 ( .A(n1429), .ZN(n1426) );
  AOI221_X1 U1089 ( .B1(n1124), .B2(hwdata_o[11]), .C1(n1125), .C2(n1430), .A(
        n1431), .ZN(n13846) );
  OAI21_X1 U1090 ( .B1(n1432), .B2(n4755), .A(irq_i[11]), .ZN(n1431) );
  INV_X1 U1092 ( .A(irq_i[10]), .ZN(n1435) );
  OAI22_X1 U1093 ( .A1(n1436), .A2(n1314), .B1(n236), .B2(n1385), .ZN(n1434)
         );
  NAND2_X1 U1094 ( .A1(n17093), .A2(n1122), .ZN(n1433) );
  INV_X1 U1096 ( .A(irq_i[8]), .ZN(n1440) );
  OAI22_X1 U1097 ( .A1(n1441), .A2(n1314), .B1(n232), .B2(n1385), .ZN(n1439)
         );
  NAND2_X1 U1098 ( .A1(n17093), .A2(n1120), .ZN(n1438) );
  INV_X1 U1099 ( .A(n1441), .ZN(n1120) );
  OAI22_X1 U1101 ( .A1(n1445), .A2(n1314), .B1(n240), .B2(n1385), .ZN(n1443)
         );
  NAND2_X1 U1102 ( .A1(n17093), .A2(n1446), .ZN(n1442) );
  AOI221_X1 U1104 ( .B1(n1314), .B2(n210), .C1(n1451), .C2(n1452), .A(n1317), 
        .ZN(n1450) );
  INV_X1 U1105 ( .A(irq_i[1]), .ZN(n1449) );
  NAND2_X1 U1106 ( .A1(n17093), .A2(n1453), .ZN(n1448) );
  AND3_X1 U1107 ( .A1(irq_i[14]), .A2(n1454), .A3(n1455), .ZN(n13747) );
  OAI21_X1 U1108 ( .B1(n200), .B2(n1456), .A(n5619), .ZN(n1455) );
  INV_X1 U1109 ( .A(n1457), .ZN(n1454) );
  AOI211_X1 U1110 ( .C1(n1314), .C2(n245), .A(n1317), .B(n1458), .ZN(n1457) );
  AOI21_X1 U1111 ( .B1(hwdata_o[14]), .B2(n1124), .A(n1459), .ZN(n1458) );
  AOI22_X1 U1113 ( .A1(n1460), .A2(n1461), .B1(n4950), .B2(n17126), .ZN(n11746) );
  NOR3_X1 U1114 ( .A1(n1462), .A2(n1463), .A3(n1464), .ZN(n1461) );
  OAI33_X1 U1115 ( .A1(n1465), .A2(n5165), .A3(n16847), .B1(n1254), .B2(n1218), 
        .B3(n617), .ZN(n1464) );
  OAI33_X1 U1116 ( .A1(n569), .A2(n16802), .A3(n723), .B1(n1466), .B2(n1467), 
        .B3(n640), .ZN(n1463) );
  NAND2_X1 U1117 ( .A1(n16856), .A2(n16864), .ZN(n1466) );
  NAND3_X1 U1118 ( .A1(n1468), .A2(n632), .A3(n1469), .ZN(n569) );
  OR4_X1 U1119 ( .A1(n1470), .A2(n1471), .A3(n1472), .A4(n1473), .ZN(n1462) );
  NOR2_X1 U1120 ( .A1(n1474), .A2(n1475), .ZN(n1460) );
  OAI211_X1 U1121 ( .C1(n605), .C2(n694), .A(n1476), .B(n1477), .ZN(n1475) );
  INV_X1 U1122 ( .A(n1271), .ZN(n1477) );
  NAND3_X1 U1123 ( .A1(n988), .A2(n619), .A3(n17123), .ZN(n1271) );
  NAND2_X1 U1124 ( .A1(n1478), .A2(n16826), .ZN(n988) );
  OAI221_X1 U1125 ( .B1(n1479), .B2(n624), .C1(n1480), .C2(n16808), .A(n1481), 
        .ZN(n1474) );
  AOI22_X1 U1126 ( .A1(n526), .A2(n1482), .B1(n540), .B2(n1483), .ZN(n1481) );
  OAI211_X1 U1127 ( .C1(n1484), .C2(n1485), .A(n1486), .B(n941), .ZN(n1483) );
  NAND3_X1 U1128 ( .A1(n833), .A2(n473), .A3(n834), .ZN(n1485) );
  XOR2_X1 U1129 ( .A(n659), .B(n16801), .Z(n834) );
  NAND3_X1 U1130 ( .A1(n16814), .A2(n16802), .A3(n505), .ZN(n1484) );
  INV_X1 U1131 ( .A(n677), .ZN(n540) );
  NAND2_X1 U1132 ( .A1(n16680), .A2(n16659), .ZN(n677) );
  OAI22_X1 U1133 ( .A1(n16820), .A2(n745), .B1(n1205), .B2(n640), .ZN(n1482)
         );
  INV_X1 U1134 ( .A(n1487), .ZN(n1205) );
  NOR4_X1 U1135 ( .A1(n1488), .A2(n1489), .A3(n1490), .A4(n1491), .ZN(n1480)
         );
  AND3_X1 U1136 ( .A1(n697), .A2(n4974), .A3(n465), .ZN(n1489) );
  INV_X1 U1137 ( .A(n478), .ZN(n465) );
  NOR2_X1 U1138 ( .A1(n16803), .A2(n16812), .ZN(n697) );
  OAI22_X1 U1139 ( .A1(n860), .A2(n818), .B1(n846), .B2(n499), .ZN(n1488) );
  AOI222_X1 U1140 ( .A1(n1492), .A2(n1493), .B1(n475), .B2(n1494), .C1(n1495), 
        .C2(n16659), .ZN(n1479) );
  OAI22_X1 U1141 ( .A1(n1496), .A2(n16802), .B1(n1497), .B2(n1498), .ZN(n1495)
         );
  NAND2_X1 U1142 ( .A1(n16807), .A2(n444), .ZN(n1498) );
  NAND2_X1 U1143 ( .A1(n731), .A2(n16733), .ZN(n444) );
  INV_X1 U1144 ( .A(n674), .ZN(n1497) );
  XOR2_X1 U1145 ( .A(n1499), .B(n17099), .Z(n674) );
  OAI211_X1 U1146 ( .C1(n1500), .C2(n1501), .A(n1502), .B(n1503), .ZN(n1499)
         );
  XOR2_X1 U1147 ( .A(n1504), .B(n1505), .Z(n1503) );
  AND3_X1 U1148 ( .A1(n1506), .A2(n843), .A3(n680), .ZN(n1505) );
  AOI22_X1 U1149 ( .A1(vis_apsr_o[3]), .A2(n1508), .B1(n1509), .B2(n1510), 
        .ZN(n1506) );
  OAI211_X1 U1150 ( .C1(n731), .C2(n16733), .A(n843), .B(n1511), .ZN(n1504) );
  OAI22_X1 U1151 ( .A1(vis_apsr_o[0]), .A2(n92), .B1(n85), .B2(n1512), .ZN(
        n1511) );
  AOI222_X1 U1152 ( .A1(n16688), .A2(U186_Z_0), .B1(n4949), .B2(n94), .C1(n93), 
        .C2(n27), .ZN(n1512) );
  INV_X1 U1153 ( .A(n93), .ZN(n4949) );
  NAND2_X1 U1154 ( .A1(n1513), .A2(n1514), .ZN(n93) );
  INV_X1 U1155 ( .A(n85), .ZN(n92) );
  NOR2_X1 U1156 ( .A1(n1515), .A2(n1516), .ZN(n85) );
  OAI33_X1 U1157 ( .A1(n1517), .A2(n16868), .A3(n653), .B1(n1518), .B2(n16823), 
        .B3(n1519), .ZN(n1516) );
  OAI211_X1 U1158 ( .C1(n16796), .C2(n16814), .A(n16816), .B(n1520), .ZN(n1502) );
  AOI221_X1 U1159 ( .B1(n1521), .B2(vis_apsr_o[1]), .C1(n1524), .C2(n1525), 
        .A(n736), .ZN(n1520) );
  AOI21_X1 U1160 ( .B1(n16796), .B2(n16733), .A(n720), .ZN(n1501) );
  AOI22_X1 U1161 ( .A1(n1526), .A2(n1509), .B1(n1527), .B2(n1508), .ZN(n1500)
         );
  XOR2_X1 U1162 ( .A(n931), .B(n4954), .Z(n1527) );
  INV_X1 U1163 ( .A(n1508), .ZN(n1509) );
  XOR2_X1 U1164 ( .A(n679), .B(n1528), .Z(n1526) );
  INV_X1 U1165 ( .A(n931), .ZN(n679) );
  NAND2_X1 U1166 ( .A1(n16816), .A2(n16812), .ZN(n931) );
  AOI221_X1 U1167 ( .B1(n1529), .B2(n1530), .C1(n736), .C2(n17099), .A(n1531), 
        .ZN(n1496) );
  NAND2_X1 U1168 ( .A1(n582), .A2(n16683), .ZN(n1531) );
  NOR2_X1 U1169 ( .A1(n16657), .A2(n16733), .ZN(n736) );
  NOR3_X1 U1170 ( .A1(n923), .A2(n16815), .A3(n16814), .ZN(n1530) );
  NOR3_X1 U1171 ( .A1(n781), .A2(n712), .A3(n659), .ZN(n1529) );
  NAND2_X1 U1172 ( .A1(n1532), .A2(n16799), .ZN(n712) );
  OAI21_X1 U1173 ( .B1(n16812), .B2(n16795), .A(n16807), .ZN(n1494) );
  NAND3_X1 U1174 ( .A1(n720), .A2(n16795), .A3(n1533), .ZN(n1493) );
  AOI221_X1 U1175 ( .B1(n16797), .B2(n16800), .C1(n721), .C2(n17098), .A(n1238), .ZN(n1533) );
  INV_X1 U1176 ( .A(n669), .ZN(n1238) );
  AOI21_X1 U1177 ( .B1(n16866), .B2(n17127), .A(n1534), .ZN(n10553) );
  NOR4_X1 U1178 ( .A1(n1535), .A2(n1536), .A3(n1537), .A4(n1538), .ZN(n1534)
         );
  OAI221_X1 U1179 ( .B1(n16859), .B2(n762), .C1(n715), .C2(n813), .A(n1539), 
        .ZN(n1538) );
  AOI21_X1 U1180 ( .B1(n1540), .B2(n16686), .A(n1201), .ZN(n1539) );
  OAI211_X1 U1181 ( .C1(n585), .C2(n1541), .A(n17123), .B(n1542), .ZN(n1201)
         );
  NOR3_X1 U1182 ( .A1(n1543), .A2(n1471), .A3(n484), .ZN(n1542) );
  INV_X1 U1183 ( .A(n512), .ZN(n484) );
  NOR3_X1 U1184 ( .A1(n16856), .A2(n16823), .A3(n16680), .ZN(n1543) );
  OAI221_X1 U1185 ( .B1(n649), .B2(n818), .C1(n606), .C2(n1465), .A(n1544), 
        .ZN(n1537) );
  AOI222_X1 U1186 ( .A1(n1172), .A2(n16866), .B1(n822), .B2(n1545), .C1(n708), 
        .C2(n1546), .ZN(n1544) );
  NAND4_X1 U1187 ( .A1(n731), .A2(n16799), .A3(n1547), .A4(n1548), .ZN(n1546)
         );
  AOI211_X1 U1188 ( .C1(n1549), .C2(n16733), .A(n5244), .B(n718), .ZN(n1548)
         );
  INV_X1 U1189 ( .A(n1550), .ZN(n718) );
  NAND3_X1 U1190 ( .A1(n709), .A2(n16801), .A3(n5243), .ZN(n1549) );
  INV_X1 U1191 ( .A(n923), .ZN(n709) );
  NAND4_X1 U1192 ( .A1(n4967), .A2(n5026), .A3(n5241), .A4(n16794), .ZN(n923)
         );
  OAI211_X1 U1193 ( .C1(n16804), .C2(n1551), .A(n1552), .B(n16811), .ZN(n1545)
         );
  NOR3_X1 U1194 ( .A1(n1553), .A2(n16733), .A3(n722), .ZN(n1551) );
  OAI21_X1 U1195 ( .B1(n16686), .B2(n832), .A(n1554), .ZN(n722) );
  OAI21_X1 U1196 ( .B1(n551), .B2(n16686), .A(n16817), .ZN(n1554) );
  INV_X1 U1197 ( .A(n668), .ZN(n551) );
  NAND3_X1 U1198 ( .A1(n16798), .A2(n454), .A3(n1555), .ZN(n668) );
  NAND2_X1 U1199 ( .A1(n16657), .A2(n16798), .ZN(n832) );
  OAI211_X1 U1200 ( .C1(n1550), .C2(n1556), .A(n548), .B(n1557), .ZN(n1553) );
  NAND3_X1 U1201 ( .A1(n16796), .A2(n16686), .A3(n721), .ZN(n1557) );
  NAND2_X1 U1202 ( .A1(n939), .A2(n16657), .ZN(n548) );
  NAND2_X1 U1203 ( .A1(n720), .A2(n16800), .ZN(n1556) );
  NAND2_X1 U1204 ( .A1(n16801), .A2(n17099), .ZN(n1550) );
  OAI221_X1 U1205 ( .B1(n16866), .B2(n1558), .C1(n16803), .C2(n1559), .A(n1560), .ZN(n1536) );
  AOI22_X1 U1206 ( .A1(n543), .A2(n1561), .B1(n884), .B2(n1094), .ZN(n1560) );
  AOI222_X1 U1207 ( .A1(n731), .A2(n791), .B1(n1216), .B2(n16871), .C1(n720), 
        .C2(n732), .ZN(n1559) );
  INV_X1 U1208 ( .A(n843), .ZN(n720) );
  NAND2_X1 U1209 ( .A1(n16796), .A2(n16815), .ZN(n843) );
  INV_X1 U1210 ( .A(n1562), .ZN(n1216) );
  AOI221_X1 U1211 ( .B1(n1563), .B2(n563), .C1(n1564), .C2(n16868), .A(n1565), 
        .ZN(n1558) );
  OAI22_X1 U1212 ( .A1(n1467), .A2(n859), .B1(n5165), .B2(n995), .ZN(n1565) );
  NAND4_X1 U1213 ( .A1(n1566), .A2(n1308), .A3(n1567), .A4(n1568), .ZN(n1535)
         );
  AOI22_X1 U1214 ( .A1(n936), .A2(n16813), .B1(n746), .B2(n1487), .ZN(n1568)
         );
  NAND2_X1 U1215 ( .A1(n5230), .A2(n16820), .ZN(n1487) );
  OAI21_X1 U1216 ( .B1(n1172), .B2(n527), .A(n16855), .ZN(n1567) );
  INV_X1 U1217 ( .A(n699), .ZN(n1172) );
  OAI21_X1 U1218 ( .B1(n1569), .B2(n483), .A(n16834), .ZN(n1566) );
  OAI211_X1 U1219 ( .C1(n1570), .C2(n17126), .A(n1571), .B(n1572), .ZN(n10055)
         );
  AOI22_X1 U1220 ( .A1(n1573), .A2(n16862), .B1(n17126), .B2(n16841), .ZN(
        n1572) );
  NAND3_X1 U1221 ( .A1(n1574), .A2(n16856), .A3(n687), .ZN(n1571) );
  NOR4_X1 U1222 ( .A1(n1575), .A2(n1576), .A3(n1577), .A4(n1578), .ZN(n1570)
         );
  NOR4_X1 U1223 ( .A1(n714), .A2(n1579), .A3(n1580), .A4(n1035), .ZN(n1578) );
  INV_X1 U1224 ( .A(n660), .ZN(n1035) );
  INV_X1 U1225 ( .A(n610), .ZN(n714) );
  NOR4_X1 U1226 ( .A1(n16866), .A2(n994), .A3(n610), .A4(n995), .ZN(n1577) );
  OAI22_X1 U1227 ( .A1(n1581), .A2(n1086), .B1(n1254), .B2(n1582), .ZN(n1576)
         );
  NAND2_X1 U1228 ( .A1(n592), .A2(n632), .ZN(n1582) );
  NAND3_X1 U1229 ( .A1(n483), .A2(n16802), .A3(n630), .ZN(n1254) );
  AOI22_X1 U1230 ( .A1(n1090), .A2(n590), .B1(n1583), .B2(n16866), .ZN(n1581)
         );
  NOR2_X1 U1231 ( .A1(n606), .A2(n16830), .ZN(n1090) );
  OAI221_X1 U1232 ( .B1(n1584), .B2(n16821), .C1(n1585), .C2(n616), .A(n1586), 
        .ZN(n1575) );
  AOI21_X1 U1233 ( .B1(n16680), .B2(n1587), .A(n1588), .ZN(n1586) );
  AOI21_X1 U1234 ( .B1(n618), .B2(n1589), .A(n16831), .ZN(n1588) );
  NAND3_X1 U1235 ( .A1(n827), .A2(n16854), .A3(n612), .ZN(n1589) );
  INV_X1 U1236 ( .A(n644), .ZN(n612) );
  NAND2_X1 U1237 ( .A1(n897), .A2(n597), .ZN(n644) );
  NAND2_X1 U1238 ( .A1(n483), .A2(n897), .ZN(n618) );
  OAI221_X1 U1239 ( .B1(n443), .B2(n1562), .C1(n16814), .C2(n892), .A(n1590), 
        .ZN(n1587) );
  OR3_X1 U1240 ( .A1(n863), .A2(n650), .A3(n662), .ZN(n1590) );
  NOR4_X1 U1241 ( .A1(n1591), .A2(n1592), .A3(n730), .A4(n1593), .ZN(n1585) );
  NOR3_X1 U1242 ( .A1(n1594), .A2(n1595), .A3(n603), .ZN(n1593) );
  AOI211_X1 U1243 ( .C1(n1596), .C2(n17098), .A(n625), .B(n1597), .ZN(n1595)
         );
  NOR3_X1 U1244 ( .A1(n469), .A2(n16799), .A3(n1532), .ZN(n1597) );
  INV_X1 U1245 ( .A(n1022), .ZN(n1532) );
  NAND2_X1 U1246 ( .A1(n16801), .A2(n16686), .ZN(n1022) );
  NAND3_X1 U1247 ( .A1(n582), .A2(n669), .A3(n1598), .ZN(n1596) );
  AOI22_X1 U1248 ( .A1(n16800), .A2(n16817), .B1(n16801), .B2(n16796), .ZN(
        n1598) );
  OAI21_X1 U1249 ( .B1(n16812), .B2(n1599), .A(n1600), .ZN(n1592) );
  NAND3_X1 U1250 ( .A1(n708), .A2(n16807), .A3(n16797), .ZN(n1600) );
  AOI221_X1 U1251 ( .B1(n629), .B2(n16683), .C1(n708), .C2(n16815), .A(n1601), 
        .ZN(n1599) );
  OAI33_X1 U1252 ( .A1(n329), .A2(n503), .A3(n16657), .B1(n711), .B2(n16868), 
        .B3(n16815), .ZN(n1601) );
  OAI222_X1 U1253 ( .A1(n725), .A2(n329), .B1(n16802), .B2(n512), .C1(n821), 
        .C2(n580), .ZN(n1591) );
  NAND2_X1 U1254 ( .A1(n16871), .A2(n503), .ZN(n512) );
  NOR4_X1 U1255 ( .A1(n1602), .A2(n546), .A3(n848), .A4(n1200), .ZN(n1584) );
  NOR3_X1 U1256 ( .A1(n713), .A2(n649), .A3(n1603), .ZN(n848) );
  OAI211_X1 U1257 ( .C1(n556), .C2(n1217), .A(n1604), .B(n1177), .ZN(n1602) );
  OAI21_X1 U1258 ( .B1(n1605), .B2(n1606), .A(n543), .ZN(n1604) );
  INV_X1 U1261 ( .A(hprot_o[3]), .ZN(n1609) );
  OAI21_X1 U1262 ( .B1(haddr_o[28]), .B2(n1610), .A(n999), .ZN(n1608) );
  OR2_X1 U1263 ( .A1(n1611), .A2(hprot_o[0]), .ZN(n999) );
  AOI21_X1 U1268 ( .B1(n1618), .B2(haddr_o[29]), .A(n1619), .ZN(n1616) );
  INV_X1 U1269 ( .A(n1620), .ZN(n1619) );
  AOI22_X1 U1272 ( .A1(n17088), .A2(n16727), .B1(add_2072_SUM_7_), .B2(n17090), 
        .ZN(n1623) );
  AOI22_X1 U1274 ( .A1(add_2072_SUM_6_), .A2(n17091), .B1(n17088), .B2(n16722), 
        .ZN(n1626) );
  AOI221_X1 U1276 ( .B1(n1627), .B2(n1628), .C1(n16726), .C2(n17087), .A(n1629), .ZN(n1147) );
  AND2_X1 U1277 ( .A1(add_2072_SUM_5_), .A2(n17091), .ZN(n1629) );
  NAND2_X1 U1279 ( .A1(add_2072_SUM_4_), .A2(n17091), .ZN(n1633) );
  AND2_X1 U1282 ( .A1(add_2072_SUM_3_), .A2(n17091), .ZN(n1635) );
  AND2_X1 U1285 ( .A1(add_2072_SUM_2_), .A2(n17091), .ZN(n1637) );
  AOI22_X1 U1287 ( .A1(n17088), .A2(n16682), .B1(add_2072_SUM_1_), .B2(n17090), 
        .ZN(n1639) );
  AND3_X1 U1290 ( .A1(n1642), .A2(n1004), .A3(n17090), .ZN(n1641) );
  OR3_X1 U1291 ( .A1(n1106), .A2(n4973), .A3(n1643), .ZN(n1004) );
  OAI21_X1 U1292 ( .B1(n4973), .B2(n1106), .A(n1643), .ZN(n1642) );
  XOR2_X1 U1293 ( .A(n1003), .B(vis_pc_o[1]), .Z(n1643) );
  AOI222_X1 U1295 ( .A1(add_2072_SUM_25_), .A2(n17089), .B1(n1628), .B2(n1644), 
        .C1(n17086), .C2(n16698), .ZN(n1148) );
  AND2_X1 U1298 ( .A1(add_2072_SUM_24_), .A2(n17090), .ZN(n1646) );
  AOI222_X1 U1300 ( .A1(add_2072_SUM_23_), .A2(n17089), .B1(n1628), .B2(n1647), 
        .C1(n17086), .C2(n16655), .ZN(n1150) );
  AOI222_X1 U1302 ( .A1(add_2072_SUM_22_), .A2(n17089), .B1(n1628), .B2(n1648), 
        .C1(n17086), .C2(n16701), .ZN(n317) );
  AOI222_X1 U1304 ( .A1(add_2072_SUM_21_), .A2(n17089), .B1(n1628), .B2(n1649), 
        .C1(n17086), .C2(n16705), .ZN(n973) );
  AOI222_X1 U1306 ( .A1(add_2072_SUM_20_), .A2(n17089), .B1(n1628), .B2(n1650), 
        .C1(n17086), .C2(n16702), .ZN(n1153) );
  AND2_X1 U1309 ( .A1(add_2072_SUM_19_), .A2(n17090), .ZN(n1652) );
  AOI222_X1 U1311 ( .A1(add_2072_SUM_18_), .A2(n17089), .B1(n1628), .B2(n1653), 
        .C1(n17086), .C2(n16706), .ZN(n1155) );
  NAND2_X1 U1314 ( .A1(add_2072_SUM_17_), .A2(n17091), .ZN(n1656) );
  AOI222_X1 U1316 ( .A1(add_2072_SUM_16_), .A2(n17089), .B1(n1628), .B2(n1657), 
        .C1(n17086), .C2(n16672), .ZN(n1157) );
  AND2_X1 U1319 ( .A1(add_2072_SUM_15_), .A2(n17090), .ZN(n1659) );
  AOI222_X1 U1321 ( .A1(add_2072_SUM_14_), .A2(n17089), .B1(n1628), .B2(n1660), 
        .C1(n17086), .C2(n16711), .ZN(n1159) );
  AOI22_X1 U1323 ( .A1(add_2072_SUM_13_), .A2(n17091), .B1(n17087), .B2(n16715), .ZN(n1662) );
  AOI222_X1 U1325 ( .A1(add_2072_SUM_12_), .A2(n17089), .B1(n1628), .B2(n1663), 
        .C1(n17086), .C2(n16658), .ZN(n956) );
  AOI222_X1 U1327 ( .A1(add_2072_SUM_11_), .A2(n17089), .B1(n1628), .B2(n1664), 
        .C1(n17086), .C2(n16679), .ZN(n957) );
  AND2_X1 U1330 ( .A1(add_2072_SUM_10_), .A2(n17090), .ZN(n1666) );
  AND2_X1 U1333 ( .A1(add_2072_SUM_8_), .A2(n17090), .ZN(n1668) );
  NOR2_X1 U1335 ( .A1(n17084), .A2(n1625), .ZN(add_2082_A_9_) );
  NOR2_X1 U1336 ( .A1(n17083), .A2(n1672), .ZN(add_2082_A_8_) );
  NOR2_X1 U1337 ( .A1(n17083), .A2(n1630), .ZN(add_2082_A_7_) );
  NOR2_X1 U1338 ( .A1(n17083), .A2(n1673), .ZN(add_2082_A_6_) );
  NOR2_X1 U1339 ( .A1(n17083), .A2(n1674), .ZN(add_2082_A_5_) );
  NOR2_X1 U1340 ( .A1(n17083), .A2(n1638), .ZN(add_2082_A_4_) );
  NOR3_X1 U1341 ( .A1(n1675), .A2(n17083), .A3(n1676), .ZN(add_2082_A_3_) );
  NOR3_X1 U1342 ( .A1(n890), .A2(n4950), .A3(n16847), .ZN(n1675) );
  NOR2_X1 U1343 ( .A1(n17083), .A2(n1677), .ZN(add_2082_A_31_) );
  NOR2_X1 U1344 ( .A1(n17083), .A2(n1678), .ZN(add_2082_A_30_) );
  NOR2_X1 U1345 ( .A1(n17083), .A2(n1679), .ZN(add_2082_A_2_) );
  NOR2_X1 U1346 ( .A1(n17083), .A2(n1680), .ZN(add_2082_A_29_) );
  NOR2_X1 U1347 ( .A1(n17083), .A2(n1681), .ZN(add_2082_A_28_) );
  NOR2_X1 U1348 ( .A1(n17084), .A2(n1682), .ZN(add_2082_A_27_) );
  NOR2_X1 U1349 ( .A1(n1683), .A2(n17085), .ZN(add_2082_A_26_) );
  NOR2_X1 U1350 ( .A1(n17084), .A2(n1684), .ZN(add_2082_A_25_) );
  NOR2_X1 U1351 ( .A1(n17084), .A2(n1685), .ZN(add_2082_A_24_) );
  NOR2_X1 U1352 ( .A1(n17084), .A2(n1686), .ZN(add_2082_A_23_) );
  NOR2_X1 U1353 ( .A1(n17084), .A2(n1687), .ZN(add_2082_A_22_) );
  NOR2_X1 U1354 ( .A1(n17084), .A2(n1688), .ZN(add_2082_A_21_) );
  NOR2_X1 U1355 ( .A1(n17084), .A2(n1654), .ZN(add_2082_A_20_) );
  NOR2_X1 U1356 ( .A1(n17084), .A2(n1689), .ZN(add_2082_A_1_) );
  NOR2_X1 U1357 ( .A1(n17084), .A2(n1690), .ZN(add_2082_A_19_) );
  NOR2_X1 U1358 ( .A1(n17084), .A2(n1691), .ZN(add_2082_A_18_) );
  NOR2_X1 U1359 ( .A1(n17084), .A2(n1692), .ZN(add_2082_A_17_) );
  NOR2_X1 U1360 ( .A1(n17085), .A2(n1661), .ZN(add_2082_A_16_) );
  NOR2_X1 U1361 ( .A1(n1693), .A2(n17085), .ZN(add_2082_A_15_) );
  AND2_X1 U1362 ( .A1(n1664), .A2(n1514), .ZN(add_2082_A_14_) );
  NOR2_X1 U1363 ( .A1(n17085), .A2(n1694), .ZN(add_2082_A_13_) );
  NOR2_X1 U1364 ( .A1(n17085), .A2(n1695), .ZN(add_2082_A_12_) );
  NOR2_X1 U1365 ( .A1(n17085), .A2(n1696), .ZN(add_2082_A_11_) );
  NOR2_X1 U1366 ( .A1(n17083), .A2(n1621), .ZN(add_2082_A_10_) );
  NAND4_X1 U1368 ( .A1(n662), .A2(n1697), .A3(n1698), .A4(n1699), .ZN(n1514)
         );
  AOI221_X1 U1369 ( .B1(n827), .B2(n16828), .C1(n1095), .C2(n16858), .A(n1700), 
        .ZN(n1699) );
  OAI22_X1 U1370 ( .A1(n16859), .A2(n696), .B1(n585), .B2(n16805), .ZN(n1700)
         );
  AOI22_X1 U1371 ( .A1(n1701), .A2(n1702), .B1(n1097), .B2(n1574), .ZN(n1698)
         );
  OAI211_X1 U1372 ( .C1(n16853), .C2(n16805), .A(n1303), .B(n998), .ZN(n1702)
         );
  OAI21_X1 U1373 ( .B1(n532), .B2(n617), .A(n16690), .ZN(n1701) );
  NAND2_X1 U1374 ( .A1(n526), .A2(n16839), .ZN(n662) );
  NOR2_X1 U1375 ( .A1(n4950), .A2(n1703), .ZN(add_2073_B_1_) );
  AOI211_X1 U1376 ( .C1(n589), .C2(n565), .A(n1704), .B(n1705), .ZN(n1703) );
  OAI221_X1 U1377 ( .B1(n1706), .B2(n1707), .C1(n16869), .C2(n1708), .A(n1709), 
        .ZN(n1704) );
  OR4_X1 U1378 ( .A1(n1278), .A2(n653), .A3(n16844), .A4(n16865), .ZN(n1709)
         );
  INV_X1 U1379 ( .A(n1710), .ZN(n1708) );
  OAI22_X1 U1380 ( .A1(n863), .A2(n16837), .B1(n1711), .B2(n4953), .ZN(n1710)
         );
  AOI22_X1 U1381 ( .A1(n16829), .A2(n16851), .B1(n16866), .B2(n1712), .ZN(
        n1711) );
  NAND2_X1 U1382 ( .A1(n1564), .A2(n16825), .ZN(n1707) );
  OAI22_X1 U1383 ( .A1(n5259), .A2(n1713), .B1(n1714), .B2(n1715), .ZN(U98_Z_0) );
  AOI211_X1 U1384 ( .C1(n1716), .C2(n659), .A(n1717), .B(n1718), .ZN(n1714) );
  OAI22_X1 U1385 ( .A1(n5253), .A2(n532), .B1(n5241), .B2(n1719), .ZN(n1718)
         );
  OAI221_X1 U1386 ( .B1(n776), .B2(n1307), .C1(n17099), .C2(n819), .A(n1720), 
        .ZN(n1717) );
  INV_X1 U1387 ( .A(n1721), .ZN(n1716) );
  OAI22_X1 U1388 ( .A1(n5544), .A2(n1713), .B1(n1722), .B2(n1715), .ZN(U97_Z_0) );
  AOI211_X1 U1389 ( .C1(n597), .C2(n1723), .A(n1724), .B(n1725), .ZN(n1722) );
  INV_X1 U1390 ( .A(n1720), .ZN(n1725) );
  OAI211_X1 U1391 ( .C1(n16794), .C2(n1719), .A(n1726), .B(n1727), .ZN(n1724)
         );
  NAND3_X1 U1392 ( .A1(n16817), .A2(n16674), .A3(n1728), .ZN(n1727) );
  OAI21_X1 U1393 ( .B1(n1729), .B2(n1730), .A(n614), .ZN(n1726) );
  INV_X1 U1394 ( .A(n664), .ZN(n1730) );
  NOR3_X1 U1395 ( .A1(n776), .A2(n16810), .A3(n16806), .ZN(n1729) );
  AOI22_X1 U1397 ( .A1(n17088), .A2(n16719), .B1(add_2072_SUM_9_), .B2(n17090), 
        .ZN(n1731) );
  OAI21_X1 U1398 ( .B1(n5120), .B2(n1732), .A(n1733), .ZN(U811_Z_0) );
  OAI21_X1 U1399 ( .B1(n1734), .B2(n1735), .A(n1732), .ZN(n1733) );
  OAI221_X1 U1400 ( .B1(n4967), .B2(n1736), .C1(n16856), .C2(n650), .A(n1737), 
        .ZN(n1735) );
  AOI222_X1 U1401 ( .A1(n1738), .A2(n413), .B1(n1739), .B2(n16674), .C1(n5120), 
        .C2(n1740), .ZN(n1737) );
  INV_X1 U1403 ( .A(n1741), .ZN(n1736) );
  NAND4_X1 U1404 ( .A1(n890), .A2(n857), .A3(n1742), .A4(n1743), .ZN(n1734) );
  AOI21_X1 U1405 ( .B1(n1744), .B2(n1745), .A(n1746), .ZN(n1743) );
  OAI33_X1 U1406 ( .A1(n514), .A2(n16845), .A3(n16858), .B1(n941), .B2(n16683), 
        .B3(n1184), .ZN(n1746) );
  XOR2_X1 U1407 ( .A(n1747), .B(n1748), .Z(n1744) );
  NAND2_X1 U1408 ( .A1(n543), .A2(n897), .ZN(n857) );
  OAI22_X1 U1409 ( .A1(n4987), .A2(n17080), .B1(n1750), .B2(n17081), .ZN(
        U810_Z_0) );
  OAI22_X1 U1410 ( .A1(n1752), .A2(n17126), .B1(n4953), .B2(n1753), .ZN(
        U809_Z_0) );
  AOI21_X1 U1411 ( .B1(n1521), .B2(n84), .A(n17127), .ZN(n1753) );
  INV_X1 U1412 ( .A(n1525), .ZN(n1521) );
  AOI221_X1 U1413 ( .B1(n86), .B2(n1754), .C1(n88), .C2(n1755), .A(n1756), 
        .ZN(n1752) );
  AND3_X1 U1414 ( .A1(n84), .A2(n1525), .A3(n1524), .ZN(n1756) );
  INV_X1 U1415 ( .A(n1757), .ZN(n1524) );
  AOI22_X1 U1416 ( .A1(n1758), .A2(n1759), .B1(U4_DATA1_0), .B2(n4947), .ZN(
        n1757) );
  OAI22_X1 U1417 ( .A1(n1760), .A2(n1761), .B1(n4953), .B2(n1762), .ZN(n1758)
         );
  INV_X1 U1418 ( .A(n1762), .ZN(n1761) );
  NAND2_X1 U1419 ( .A1(n1763), .A2(n1764), .ZN(n1762) );
  AOI21_X1 U1420 ( .B1(n1765), .B2(n1766), .A(n1767), .ZN(n1760) );
  AOI211_X1 U1421 ( .C1(n1768), .C2(n16833), .A(n1765), .B(n1769), .ZN(n1767)
         );
  NOR3_X1 U1422 ( .A1(n1770), .A2(n16833), .A3(n1771), .ZN(n1769) );
  NOR3_X1 U1423 ( .A1(n1772), .A2(n1773), .A3(n1774), .ZN(n1771) );
  INV_X1 U1424 ( .A(n1775), .ZN(n1770) );
  AOI22_X1 U1425 ( .A1(n1776), .A2(n1777), .B1(n1774), .B2(n1778), .ZN(n1775)
         );
  OAI22_X1 U1426 ( .A1(n1779), .A2(n1780), .B1(n1781), .B2(n1773), .ZN(n1778)
         );
  INV_X1 U1427 ( .A(n1782), .ZN(n1776) );
  OAI22_X1 U1428 ( .A1(n1783), .A2(n1784), .B1(n1768), .B2(n16848), .ZN(n1766)
         );
  AOI221_X1 U1429 ( .B1(n1785), .B2(n1786), .C1(n1777), .C2(n1787), .A(n1788), 
        .ZN(n1768) );
  OAI33_X1 U1430 ( .A1(n1774), .A2(n1773), .A3(n1789), .B1(n1780), .B2(n1790), 
        .B3(n1791), .ZN(n1788) );
  NOR2_X1 U1431 ( .A1(n1790), .A2(n1773), .ZN(n1785) );
  AOI21_X1 U1432 ( .B1(n1792), .B2(n1763), .A(n1764), .ZN(n1765) );
  INV_X1 U1433 ( .A(n1793), .ZN(n1764) );
  OAI21_X1 U1434 ( .B1(n1794), .B2(n1795), .A(n529), .ZN(n1792) );
  OAI221_X1 U1435 ( .B1(n1796), .B2(n16869), .C1(n1797), .C2(n16824), .A(n1798), .ZN(n1525) );
  INV_X1 U1436 ( .A(n1515), .ZN(n1798) );
  OAI221_X1 U1437 ( .B1(n606), .B2(n849), .C1(n1519), .C2(n1580), .A(n1799), 
        .ZN(n1515) );
  OAI21_X1 U1438 ( .B1(n1800), .B2(n1801), .A(n16871), .ZN(n1799) );
  NOR3_X1 U1439 ( .A1(n16826), .A2(n1104), .A3(n16864), .ZN(n1800) );
  AOI211_X1 U1440 ( .C1(n1802), .C2(n529), .A(n1803), .B(n1804), .ZN(n1797) );
  AOI21_X1 U1441 ( .B1(n1234), .B2(n16848), .A(n849), .ZN(n1804) );
  INV_X1 U1442 ( .A(n1210), .ZN(n1802) );
  AOI21_X1 U1443 ( .B1(n16866), .B2(n1805), .A(n1806), .ZN(n1796) );
  OAI22_X1 U1444 ( .A1(n4998), .A2(n17080), .B1(n1807), .B2(n17081), .ZN(
        U806_Z_0) );
  OAI22_X1 U1445 ( .A1(n4963), .A2(n17080), .B1(n1808), .B2(n17081), .ZN(
        U805_Z_0) );
  OAI22_X1 U1446 ( .A1(n5022), .A2(n17080), .B1(n1809), .B2(n17081), .ZN(
        U804_Z_0) );
  OAI22_X1 U1447 ( .A1(n5040), .A2(n17080), .B1(n1810), .B2(n17082), .ZN(
        U803_Z_0) );
  OAI22_X1 U1448 ( .A1(n5227), .A2(n980), .B1(n1669), .B2(n1811), .ZN(U802_Z_0) );
  OAI22_X1 U1449 ( .A1(n4981), .A2(n17075), .B1(n1808), .B2(n17076), .ZN(
        U801_Z_0) );
  OAI22_X1 U1450 ( .A1(n4997), .A2(n17075), .B1(n1807), .B2(n17076), .ZN(
        U800_Z_0) );
  OAI22_X1 U1451 ( .A1(n5021), .A2(n17075), .B1(n1809), .B2(n17076), .ZN(
        U799_Z_0) );
  OAI22_X1 U1452 ( .A1(n4986), .A2(n17075), .B1(n1750), .B2(n17076), .ZN(
        U798_Z_0) );
  OAI22_X1 U1453 ( .A1(n5039), .A2(n17075), .B1(n1810), .B2(n17077), .ZN(
        U797_Z_0) );
  OAI22_X1 U1454 ( .A1(n5027), .A2(n1732), .B1(n1814), .B2(n1815), .ZN(
        U795_Z_0) );
  NOR4_X1 U1455 ( .A1(n1816), .A2(n1817), .A3(n1818), .A4(n1819), .ZN(n1815)
         );
  AOI21_X1 U1456 ( .B1(n1820), .B2(n1821), .A(n788), .ZN(n1819) );
  OAI21_X1 U1457 ( .B1(n16800), .B2(n1822), .A(n1823), .ZN(n1817) );
  OAI211_X1 U1458 ( .C1(n1824), .C2(n1825), .A(n1745), .B(n1826), .ZN(n1823)
         );
  OAI221_X1 U1459 ( .B1(n4967), .B2(n1827), .C1(n5025), .C2(n1828), .A(n1829), 
        .ZN(n1816) );
  AOI22_X1 U1460 ( .A1(n1741), .A2(n461), .B1(n1830), .B2(n16674), .ZN(n1829)
         );
  OAI21_X1 U1461 ( .B1(n1113), .B2(n946), .A(n1831), .ZN(U792_Z_0) );
  NAND4_X1 U1462 ( .A1(n1111), .A2(n5149), .A3(n946), .A4(n253), .ZN(n1831) );
  INV_X1 U1463 ( .A(n256), .ZN(n946) );
  NOR4_X1 U1464 ( .A1(n1610), .A2(n1811), .A3(n1607), .A4(haddr_o[28]), .ZN(
        n256) );
  AND2_X1 U1467 ( .A1(add_2072_SUM_26_), .A2(n17090), .ZN(n1833) );
  OR4_X1 U1468 ( .A1(n978), .A2(n1834), .A3(n17089), .A4(n909), .ZN(n1607) );
  OAI21_X1 U1469 ( .B1(n1669), .B2(n1614), .A(n1835), .ZN(n978) );
  OAI22_X1 U1470 ( .A1(n1613), .A2(n1612), .B1(n327), .B2(n1836), .ZN(n1835)
         );
  INV_X1 U1471 ( .A(n683), .ZN(n1836) );
  INV_X1 U1472 ( .A(n1611), .ZN(n1613) );
  NAND3_X1 U1473 ( .A1(n1837), .A2(n1838), .A3(n1325), .ZN(n1611) );
  NOR3_X1 U1474 ( .A1(n1839), .A2(lockup_o), .A3(n1834), .ZN(n1325) );
  NAND3_X1 U1475 ( .A1(n1840), .A2(n1841), .A3(n1842), .ZN(n1834) );
  AOI221_X1 U1476 ( .B1(n1843), .B2(n746), .C1(n1094), .C2(n1844), .A(n1845), 
        .ZN(n1842) );
  NAND3_X1 U1477 ( .A1(n1177), .A2(n1846), .A3(n1092), .ZN(n1845) );
  OAI21_X1 U1478 ( .B1(n16680), .B2(n1847), .A(n522), .ZN(n1844) );
  INV_X1 U1479 ( .A(n1848), .ZN(n1847) );
  NOR2_X1 U1480 ( .A1(n860), .A2(n911), .ZN(n1843) );
  AOI222_X1 U1481 ( .A1(n16823), .A2(n1848), .B1(n799), .B2(n1849), .C1(n1850), 
        .C2(n16821), .ZN(n1841) );
  OAI211_X1 U1482 ( .C1(n860), .C2(n1851), .A(n1852), .B(n1853), .ZN(n1850) );
  AOI221_X1 U1483 ( .B1(n543), .B2(n1854), .C1(n1855), .C2(n16868), .A(n1200), 
        .ZN(n1853) );
  NOR3_X1 U1484 ( .A1(n16823), .A2(n16853), .A3(n813), .ZN(n1200) );
  NOR2_X1 U1485 ( .A1(n16859), .A2(n1784), .ZN(n1855) );
  OAI21_X1 U1486 ( .B1(n649), .B2(n16839), .A(n1856), .ZN(n1854) );
  INV_X1 U1487 ( .A(n753), .ZN(n649) );
  OAI21_X1 U1488 ( .B1(n1213), .B2(n16824), .A(n1569), .ZN(n1852) );
  INV_X1 U1489 ( .A(n818), .ZN(n1569) );
  INV_X1 U1490 ( .A(n556), .ZN(n1213) );
  INV_X1 U1491 ( .A(n746), .ZN(n1851) );
  NOR2_X1 U1492 ( .A1(n859), .A2(n16848), .ZN(n746) );
  NAND2_X1 U1493 ( .A1(n527), .A2(n610), .ZN(n859) );
  OAI22_X1 U1494 ( .A1(n16833), .A2(n715), .B1(n585), .B2(n1307), .ZN(n1849)
         );
  OAI211_X1 U1495 ( .C1(n585), .C2(n1857), .A(n1858), .B(n1859), .ZN(n1848) );
  AOI21_X1 U1496 ( .B1(n798), .B2(n527), .A(n16826), .ZN(n1859) );
  NAND3_X1 U1497 ( .A1(n728), .A2(n808), .A3(n608), .ZN(n1858) );
  AOI21_X1 U1498 ( .B1(n565), .B2(n608), .A(n701), .ZN(n1840) );
  OAI21_X1 U1499 ( .B1(n673), .B2(n522), .A(n1860), .ZN(n701) );
  OAI33_X1 U1502 ( .A1(n524), .A2(n16680), .A3(n1023), .B1(n532), .B2(n1863), 
        .B3(n16828), .ZN(n1862) );
  AOI21_X1 U1503 ( .B1(n998), .B2(n502), .A(n1864), .ZN(n1863) );
  NOR4_X1 U1504 ( .A1(n5228), .A2(n579), .A3(n617), .A4(n918), .ZN(n1864) );
  AOI21_X1 U1505 ( .B1(n1865), .B2(n1846), .A(n5228), .ZN(n1861) );
  NAND4_X1 U1506 ( .A1(n997), .A2(n991), .A3(n1574), .A4(n16853), .ZN(n1846)
         );
  INV_X1 U1507 ( .A(n1866), .ZN(n1865) );
  OAI22_X1 U1508 ( .A1(n1867), .A2(n1326), .B1(n16869), .B2(n375), .ZN(n1838)
         );
  NOR2_X1 U1510 ( .A1(n4973), .A2(n1003), .ZN(n1867) );
  OAI21_X1 U1511 ( .B1(n1007), .B2(n187), .A(n1009), .ZN(n1003) );
  OAI21_X1 U1513 ( .B1(n1326), .B2(n1001), .A(n4973), .ZN(n1837) );
  INV_X1 U1514 ( .A(n1106), .ZN(n1001) );
  NOR2_X1 U1515 ( .A1(n188), .A2(n1007), .ZN(n1326) );
  AOI21_X1 U1516 ( .B1(n16856), .B2(n1868), .A(n727), .ZN(n188) );
  INV_X1 U1517 ( .A(n327), .ZN(n1669) );
  OAI22_X1 U1518 ( .A1(n1632), .A2(n16785), .B1(n1689), .B2(n1622), .ZN(n327)
         );
  NAND3_X1 U1520 ( .A1(haddr_o[30]), .A2(haddr_o[31]), .A3(haddr_o[29]), .ZN(
        n1610) );
  NAND2_X1 U1522 ( .A1(add_2072_SUM_27_), .A2(n17091), .ZN(n1869) );
  AOI22_X1 U1523 ( .A1(n16693), .A2(n17088), .B1(n1870), .B2(n1628), .ZN(n1620) );
  INV_X1 U1525 ( .A(n1617), .ZN(n1871) );
  OAI22_X1 U1526 ( .A1(n27), .A2(n1632), .B1(n1872), .B2(n1622), .ZN(n1617) );
  INV_X1 U1527 ( .A(n16688), .ZN(n27) );
  XOR2_X1 U1528 ( .A(n5006), .B(add_2072_carry[29]), .Z(n1618) );
  NAND2_X1 U1530 ( .A1(add_2072_SUM_28_), .A2(n17091), .ZN(n1874) );
  INV_X1 U1532 ( .A(hwrite_o), .ZN(n1113) );
  OAI21_X1 U1534 ( .B1(n1879), .B2(n1880), .A(n195), .ZN(n1878) );
  NOR3_X1 U1535 ( .A1(n860), .A2(n616), .A3(n918), .ZN(n1879) );
  NOR2_X1 U1536 ( .A1(n742), .A2(n1881), .ZN(n1877) );
  NOR4_X1 U1537 ( .A1(n16808), .A2(n1882), .A3(n653), .A4(n1303), .ZN(n1881)
         );
  NOR2_X1 U1538 ( .A1(n995), .A2(n1303), .ZN(n742) );
  NAND2_X1 U1539 ( .A1(n608), .A2(n16825), .ZN(n995) );
  INV_X1 U1540 ( .A(n1883), .ZN(n1875) );
  OAI22_X1 U1541 ( .A1(n1884), .A2(n1885), .B1(n226), .B2(n1886), .ZN(U791_Z_0) );
  OAI22_X1 U1542 ( .A1(n5521), .A2(n1884), .B1(n229), .B2(n1886), .ZN(U790_Z_0) );
  OAI22_X1 U1543 ( .A1(n5151), .A2(n1884), .B1(n245), .B2(n1886), .ZN(U789_Z_0) );
  OAI22_X1 U1544 ( .A1(n5150), .A2(n1884), .B1(n247), .B2(n1886), .ZN(U788_Z_0) );
  OAI22_X1 U1545 ( .A1(n5152), .A2(n1884), .B1(n19), .B2(n1886), .ZN(U787_Z_0)
         );
  OAI22_X1 U1547 ( .A1(n5153), .A2(n1884), .B1(n1190), .B2(n1886), .ZN(
        U786_Z_0) );
  OAI22_X1 U1548 ( .A1(n5154), .A2(n1884), .B1(n1077), .B2(n1886), .ZN(
        U785_Z_0) );
  OAI22_X1 U1549 ( .A1(n5155), .A2(n1884), .B1(n1187), .B2(n1886), .ZN(
        U784_Z_0) );
  INV_X1 U1550 ( .A(n1886), .ZN(n1884) );
  OAI22_X1 U1552 ( .A1(n5518), .A2(n1888), .B1(n226), .B2(n1889), .ZN(U783_Z_0) );
  OAI22_X1 U1553 ( .A1(n5522), .A2(n1888), .B1(n229), .B2(n1889), .ZN(U782_Z_0) );
  OAI22_X1 U1554 ( .A1(n5157), .A2(n1888), .B1(n245), .B2(n1889), .ZN(U781_Z_0) );
  OAI22_X1 U1555 ( .A1(n5156), .A2(n1888), .B1(n247), .B2(n1889), .ZN(U780_Z_0) );
  OAI22_X1 U1556 ( .A1(n5158), .A2(n1888), .B1(n19), .B2(n1889), .ZN(U779_Z_0)
         );
  OAI22_X1 U1557 ( .A1(n5159), .A2(n1888), .B1(n1190), .B2(n1889), .ZN(
        U778_Z_0) );
  OAI22_X1 U1558 ( .A1(n5160), .A2(n1888), .B1(n1077), .B2(n1889), .ZN(
        U777_Z_0) );
  OAI22_X1 U1559 ( .A1(n5161), .A2(n1888), .B1(n1187), .B2(n1889), .ZN(
        U776_Z_0) );
  INV_X1 U1560 ( .A(n1889), .ZN(n1888) );
  OAI22_X1 U1562 ( .A1(n5519), .A2(n1891), .B1(n226), .B2(n1892), .ZN(U775_Z_0) );
  OAI22_X1 U1563 ( .A1(n5523), .A2(n1891), .B1(n229), .B2(n1892), .ZN(U774_Z_0) );
  OAI22_X1 U1564 ( .A1(n5046), .A2(n1891), .B1(n245), .B2(n1892), .ZN(U773_Z_0) );
  OAI22_X1 U1565 ( .A1(n5023), .A2(n1891), .B1(n247), .B2(n1892), .ZN(U772_Z_0) );
  OAI22_X1 U1566 ( .A1(n5053), .A2(n1891), .B1(n19), .B2(n1892), .ZN(U771_Z_0)
         );
  OAI22_X1 U1567 ( .A1(n5008), .A2(n1891), .B1(n1190), .B2(n1892), .ZN(
        U770_Z_0) );
  OAI22_X1 U1568 ( .A1(n5009), .A2(n1891), .B1(n1077), .B2(n1892), .ZN(
        U769_Z_0) );
  OAI22_X1 U1569 ( .A1(n5010), .A2(n1891), .B1(n1187), .B2(n1892), .ZN(
        U768_Z_0) );
  INV_X1 U1570 ( .A(n1892), .ZN(n1891) );
  OAI22_X1 U1572 ( .A1(n5548), .A2(n1894), .B1(n226), .B2(n1895), .ZN(U767_Z_0) );
  OAI22_X1 U1573 ( .A1(n5549), .A2(n1894), .B1(n229), .B2(n1895), .ZN(U766_Z_0) );
  OAI22_X1 U1574 ( .A1(n5550), .A2(n1894), .B1(n245), .B2(n1895), .ZN(U765_Z_0) );
  OAI22_X1 U1575 ( .A1(n5547), .A2(n1894), .B1(n247), .B2(n1895), .ZN(U764_Z_0) );
  OAI22_X1 U1576 ( .A1(n1894), .A2(n1896), .B1(n19), .B2(n1895), .ZN(U763_Z_0)
         );
  OAI22_X1 U1577 ( .A1(n5551), .A2(n1894), .B1(n1190), .B2(n1895), .ZN(
        U762_Z_0) );
  OAI22_X1 U1578 ( .A1(n5552), .A2(n1894), .B1(n1077), .B2(n1895), .ZN(
        U761_Z_0) );
  OAI22_X1 U1579 ( .A1(n5553), .A2(n1894), .B1(n1187), .B2(n1895), .ZN(
        U760_Z_0) );
  INV_X1 U1580 ( .A(n1895), .ZN(n1894) );
  OAI22_X1 U1582 ( .A1(n1814), .A2(n1898), .B1(n16809), .B2(n1899), .ZN(
        U756_Z_0) );
  AOI21_X1 U1583 ( .B1(n1740), .B2(n1900), .A(n1814), .ZN(n1899) );
  NOR4_X1 U1584 ( .A1(n1901), .A2(n1902), .A3(n1818), .A4(n1903), .ZN(n1898)
         );
  NOR3_X1 U1585 ( .A1(n1900), .A2(n788), .A3(n16656), .ZN(n1903) );
  INV_X1 U1586 ( .A(n1740), .ZN(n788) );
  INV_X1 U1587 ( .A(n1742), .ZN(n1818) );
  NAND2_X1 U1588 ( .A1(n527), .A2(n1904), .ZN(n1742) );
  OAI21_X1 U1589 ( .B1(n5241), .B2(n16856), .A(n605), .ZN(n1904) );
  OAI22_X1 U1590 ( .A1(n17099), .A2(n1822), .B1(n1905), .B2(n1906), .ZN(n1902)
         );
  XNOR2_X1 U1591 ( .A(n1826), .B(n1907), .ZN(n1906) );
  INV_X1 U1592 ( .A(n1745), .ZN(n1905) );
  INV_X1 U1593 ( .A(n1739), .ZN(n1822) );
  NAND2_X1 U1594 ( .A1(n1908), .A2(n1909), .ZN(n1739) );
  OAI221_X1 U1595 ( .B1(n5026), .B2(n1827), .C1(n175), .C2(n1828), .A(n1910), 
        .ZN(n1901) );
  AOI22_X1 U1596 ( .A1(n1741), .A2(n454), .B1(n1830), .B2(n16798), .ZN(n1910)
         );
  INV_X1 U1597 ( .A(n772), .ZN(n1830) );
  INV_X1 U1599 ( .A(n1732), .ZN(n1814) );
  OAI21_X1 U1600 ( .B1(n5100), .B2(n1732), .A(n1911), .ZN(U755_Z_0) );
  OAI21_X1 U1601 ( .B1(n1912), .B2(n1913), .A(n1732), .ZN(n1911) );
  OAI221_X1 U1602 ( .B1(n17099), .B2(n772), .C1(n16859), .C2(n524), .A(n1914), 
        .ZN(n1913) );
  AOI222_X1 U1603 ( .A1(n1741), .A2(n16734), .B1(n1915), .B2(n16657), .C1(
        n1738), .C2(n415), .ZN(n1914) );
  INV_X1 U1605 ( .A(n1828), .ZN(n1738) );
  OAI21_X1 U1606 ( .B1(n807), .B2(n1916), .A(n194), .ZN(n1828) );
  NOR2_X1 U1608 ( .A1(n998), .A2(n745), .ZN(n1916) );
  INV_X1 U1609 ( .A(n1909), .ZN(n1915) );
  OAI21_X1 U1610 ( .B1(n1917), .B2(n792), .A(n16811), .ZN(n1909) );
  AND2_X1 U1611 ( .A1(n936), .A2(n16820), .ZN(n792) );
  NOR2_X1 U1612 ( .A1(n1552), .A2(n16869), .ZN(n936) );
  NOR2_X1 U1613 ( .A1(n579), .A2(n478), .ZN(n1917) );
  OAI211_X1 U1614 ( .C1(n851), .C2(n945), .A(n1291), .B(n1918), .ZN(n1741) );
  AOI21_X1 U1615 ( .B1(n476), .B2(n16816), .A(n1919), .ZN(n1918) );
  NOR4_X1 U1616 ( .A1(n16814), .A2(n16659), .A3(n1261), .A4(n1184), .ZN(n1919)
         );
  AOI22_X1 U1617 ( .A1(n1920), .A2(n476), .B1(n466), .B2(n482), .ZN(n1291) );
  NOR2_X1 U1618 ( .A1(n819), .A2(n16811), .ZN(n482) );
  NAND2_X1 U1619 ( .A1(n1220), .A2(n466), .ZN(n772) );
  OAI221_X1 U1620 ( .B1(n680), .B2(n1908), .C1(n5241), .C2(n1827), .A(n1921), 
        .ZN(n1912) );
  AOI221_X1 U1621 ( .B1(n1922), .B2(n1740), .C1(n1923), .C2(n1745), .A(n799), 
        .ZN(n1921) );
  OAI33_X1 U1622 ( .A1(n1920), .A2(n16815), .A3(n443), .B1(n940), .B2(n16811), 
        .B3(n1184), .ZN(n1745) );
  NAND2_X1 U1623 ( .A1(n822), .A2(n16733), .ZN(n940) );
  OAI22_X1 U1624 ( .A1(n1924), .A2(n1925), .B1(n1907), .B2(n1826), .ZN(n1923)
         );
  NAND2_X1 U1625 ( .A1(n1824), .A2(n1825), .ZN(n1826) );
  XOR2_X1 U1626 ( .A(n1926), .B(n1927), .Z(n1825) );
  AND2_X1 U1627 ( .A1(n1748), .A2(n1747), .ZN(n1824) );
  INV_X1 U1628 ( .A(n1928), .ZN(n1747) );
  AOI21_X1 U1629 ( .B1(n1929), .B2(n16800), .A(n1927), .ZN(n1748) );
  XNOR2_X1 U1630 ( .A(n1925), .B(n1924), .ZN(n1907) );
  NAND2_X1 U1631 ( .A1(n1927), .A2(n1926), .ZN(n1925) );
  XOR2_X1 U1632 ( .A(n1930), .B(n1931), .Z(n1926) );
  NOR2_X1 U1633 ( .A1(n1929), .A2(n16799), .ZN(n1927) );
  OAI21_X1 U1634 ( .B1(n1932), .B2(n16674), .A(n1933), .ZN(n1929) );
  XOR2_X1 U1635 ( .A(n1934), .B(n1935), .Z(n1924) );
  AOI22_X1 U1636 ( .A1(n1930), .A2(n1931), .B1(n1936), .B2(n1937), .ZN(n1935)
         );
  XOR2_X1 U1637 ( .A(n1937), .B(n1936), .Z(n1931) );
  XOR2_X1 U1638 ( .A(n1938), .B(n1939), .Z(n1937) );
  INV_X1 U1639 ( .A(n1933), .ZN(n1930) );
  NAND2_X1 U1640 ( .A1(n1932), .A2(n16674), .ZN(n1933) );
  AOI21_X1 U1641 ( .B1(n1940), .B2(n5244), .A(n1936), .ZN(n1932) );
  NOR2_X1 U1642 ( .A1(n1940), .A2(n5244), .ZN(n1936) );
  OAI21_X1 U1643 ( .B1(n781), .B2(n1941), .A(n1938), .ZN(n1940) );
  OAI22_X1 U1644 ( .A1(n1939), .A2(n1938), .B1(n1942), .B2(n1943), .ZN(n1934)
         );
  NAND2_X1 U1645 ( .A1(n1941), .A2(n781), .ZN(n1938) );
  XOR2_X1 U1646 ( .A(n16794), .B(n1944), .Z(n1941) );
  XNOR2_X1 U1647 ( .A(n1943), .B(n1942), .ZN(n1939) );
  AOI21_X1 U1648 ( .B1(n454), .B2(n1945), .A(n1555), .ZN(n1942) );
  NOR2_X1 U1649 ( .A1(n4967), .A2(n5026), .ZN(n1555) );
  OR2_X1 U1650 ( .A1(n1944), .A2(n16794), .ZN(n1943) );
  XOR2_X1 U1651 ( .A(n5241), .B(n1945), .Z(n1944) );
  XNOR2_X1 U1652 ( .A(n461), .B(n4967), .ZN(n1945) );
  OAI221_X1 U1653 ( .B1(n860), .B2(n514), .C1(n16854), .C2(n1093), .A(n1309), 
        .ZN(n1740) );
  AOI22_X1 U1654 ( .A1(n16862), .A2(n1573), .B1(n589), .B2(n1946), .ZN(n1309)
         );
  INV_X1 U1655 ( .A(n1583), .ZN(n1093) );
  XOR2_X1 U1656 ( .A(n794), .B(n795), .Z(n1922) );
  NOR2_X1 U1657 ( .A1(n1900), .A2(n16809), .ZN(n794) );
  OAI21_X1 U1658 ( .B1(n1540), .B2(n732), .A(n631), .ZN(n1827) );
  INV_X1 U1659 ( .A(n1184), .ZN(n631) );
  NAND2_X1 U1660 ( .A1(n16820), .A2(n16802), .ZN(n1184) );
  NAND2_X1 U1661 ( .A1(n16812), .A2(n16657), .ZN(n680) );
  OAI21_X1 U1662 ( .B1(n1947), .B2(n17126), .A(n1948), .ZN(n1732) );
  NAND3_X1 U1663 ( .A1(n827), .A2(n911), .A3(n687), .ZN(n1948) );
  INV_X1 U1664 ( .A(n1059), .ZN(n687) );
  NAND2_X1 U1665 ( .A1(n17124), .A2(n16805), .ZN(n1059) );
  NOR4_X1 U1666 ( .A1(n1949), .A2(n1950), .A3(n1951), .A4(n1299), .ZN(n1947)
         );
  NAND4_X1 U1667 ( .A1(n1952), .A2(n1953), .A3(n1954), .A4(n1955), .ZN(n1299)
         );
  NOR4_X1 U1668 ( .A1(n1956), .A2(n1470), .A3(n1573), .A4(n1490), .ZN(n1955)
         );
  NOR4_X1 U1669 ( .A1(n1579), .A2(n16689), .A3(n585), .A4(n16853), .ZN(n1490)
         );
  INV_X1 U1670 ( .A(n1957), .ZN(n1573) );
  NOR2_X1 U1671 ( .A1(n1465), .A2(n16859), .ZN(n1470) );
  OAI22_X1 U1672 ( .A1(n1958), .A2(n503), .B1(n497), .B2(n16657), .ZN(n1956)
         );
  AOI221_X1 U1673 ( .B1(n333), .B2(n16804), .C1(n934), .C2(n1959), .A(n541), 
        .ZN(n1958) );
  NOR2_X1 U1674 ( .A1(n478), .A2(n16812), .ZN(n541) );
  INV_X1 U1675 ( .A(n1960), .ZN(n1959) );
  AOI22_X1 U1676 ( .A1(n939), .A2(n505), .B1(n731), .B2(n833), .ZN(n1960) );
  NOR2_X1 U1677 ( .A1(n16799), .A2(n16797), .ZN(n833) );
  NOR2_X1 U1678 ( .A1(n669), .A2(n17099), .ZN(n939) );
  INV_X1 U1679 ( .A(n941), .ZN(n934) );
  AOI222_X1 U1680 ( .A1(n1540), .A2(n16802), .B1(n16794), .B2(n1472), .C1(n473), .C2(n475), .ZN(n1954) );
  INV_X1 U1681 ( .A(n510), .ZN(n1952) );
  OAI211_X1 U1682 ( .C1(n1580), .C2(n1214), .A(n1961), .B(n1962), .ZN(n510) );
  AOI22_X1 U1683 ( .A1(n1472), .A2(n16837), .B1(n629), .B2(n16659), .ZN(n1962)
         );
  NAND3_X1 U1684 ( .A1(n16807), .A2(n1963), .A3(n708), .ZN(n1961) );
  NAND2_X1 U1685 ( .A1(n565), .A2(n16870), .ZN(n1214) );
  NOR2_X1 U1686 ( .A1(n1519), .A2(n696), .ZN(n1951) );
  OAI22_X1 U1687 ( .A1(n16820), .A2(n673), .B1(n1964), .B2(n692), .ZN(n1950)
         );
  OAI221_X1 U1688 ( .B1(n762), .B2(n607), .C1(n610), .C2(n699), .A(n1965), 
        .ZN(n1949) );
  NOR3_X1 U1689 ( .A1(n1966), .A2(n1491), .A3(n1967), .ZN(n1965) );
  NOR3_X1 U1690 ( .A1(n1267), .A2(n16815), .A3(n1261), .ZN(n1967) );
  NOR4_X1 U1691 ( .A1(n1307), .A2(n797), .A3(n16862), .A4(n16866), .ZN(n1491)
         );
  AND3_X1 U1692 ( .A1(n807), .A2(n808), .A3(n16837), .ZN(n1966) );
  NOR2_X1 U1693 ( .A1(n641), .A2(n17097), .ZN(n807) );
  NAND2_X1 U1694 ( .A1(n195), .A2(n16694), .ZN(n607) );
  OAI22_X1 U1695 ( .A1(n5545), .A2(n1713), .B1(n1968), .B2(n1715), .ZN(
        U754_Z_0) );
  NOR2_X1 U1696 ( .A1(n1969), .A2(n1970), .ZN(n1968) );
  OAI221_X1 U1697 ( .B1(n5243), .B2(n1721), .C1(n16800), .C2(n819), .A(n1170), 
        .ZN(n1970) );
  OAI221_X1 U1698 ( .B1(n1971), .B2(n1307), .C1(n5003), .C2(n532), .A(n1972), 
        .ZN(n1969) );
  INV_X1 U1699 ( .A(n1973), .ZN(n1972) );
  OAI21_X1 U1700 ( .B1(n1719), .B2(n5026), .A(n694), .ZN(n1973) );
  AOI221_X1 U1701 ( .B1(n1974), .B2(n776), .C1(n1975), .C2(n437), .A(n1976), 
        .ZN(n1971) );
  OAI22_X1 U1702 ( .A1(n5450), .A2(n17070), .B1(n1808), .B2(n17071), .ZN(
        U752_Z_0) );
  OAI22_X1 U1703 ( .A1(n5451), .A2(n17070), .B1(n1807), .B2(n17071), .ZN(
        U751_Z_0) );
  OAI22_X1 U1704 ( .A1(n5452), .A2(n17070), .B1(n1809), .B2(n17071), .ZN(
        U750_Z_0) );
  OAI22_X1 U1705 ( .A1(n5453), .A2(n17070), .B1(n1750), .B2(n17071), .ZN(
        U749_Z_0) );
  OAI22_X1 U1706 ( .A1(n5454), .A2(n17070), .B1(n1810), .B2(n17072), .ZN(
        U748_Z_0) );
  OAI22_X1 U1707 ( .A1(n5421), .A2(n17065), .B1(n1808), .B2(n17066), .ZN(
        U747_Z_0) );
  OAI22_X1 U1708 ( .A1(n5422), .A2(n17065), .B1(n1807), .B2(n17066), .ZN(
        U746_Z_0) );
  OAI22_X1 U1709 ( .A1(n5423), .A2(n17065), .B1(n1809), .B2(n17066), .ZN(
        U745_Z_0) );
  OAI22_X1 U1710 ( .A1(n5424), .A2(n17065), .B1(n1750), .B2(n17066), .ZN(
        U744_Z_0) );
  OAI22_X1 U1711 ( .A1(n5425), .A2(n17065), .B1(n1810), .B2(n17067), .ZN(
        U743_Z_0) );
  OAI22_X1 U1712 ( .A1(n5392), .A2(n17060), .B1(n1808), .B2(n17061), .ZN(
        U742_Z_0) );
  OAI22_X1 U1713 ( .A1(n5393), .A2(n17060), .B1(n1807), .B2(n17061), .ZN(
        U741_Z_0) );
  OAI22_X1 U1714 ( .A1(n5394), .A2(n17060), .B1(n1809), .B2(n17061), .ZN(
        U740_Z_0) );
  OAI22_X1 U1715 ( .A1(n5395), .A2(n17060), .B1(n1750), .B2(n17061), .ZN(
        U739_Z_0) );
  OAI22_X1 U1716 ( .A1(n5396), .A2(n17060), .B1(n1810), .B2(n17062), .ZN(
        U738_Z_0) );
  OAI22_X1 U1717 ( .A1(n5363), .A2(n17055), .B1(n1808), .B2(n17056), .ZN(
        U737_Z_0) );
  OAI22_X1 U1718 ( .A1(n5364), .A2(n17055), .B1(n1807), .B2(n17056), .ZN(
        U736_Z_0) );
  OAI22_X1 U1719 ( .A1(n5365), .A2(n17055), .B1(n1809), .B2(n17056), .ZN(
        U735_Z_0) );
  OAI22_X1 U1720 ( .A1(n5366), .A2(n17055), .B1(n1750), .B2(n17056), .ZN(
        U734_Z_0) );
  OAI22_X1 U1721 ( .A1(n5367), .A2(n17055), .B1(n1810), .B2(n17057), .ZN(
        U733_Z_0) );
  OAI22_X1 U1722 ( .A1(n5334), .A2(n17050), .B1(n1808), .B2(n17051), .ZN(
        U732_Z_0) );
  OAI22_X1 U1723 ( .A1(n5335), .A2(n17050), .B1(n1807), .B2(n17051), .ZN(
        U731_Z_0) );
  OAI22_X1 U1724 ( .A1(n5336), .A2(n17050), .B1(n1809), .B2(n17051), .ZN(
        U730_Z_0) );
  OAI22_X1 U1725 ( .A1(n5337), .A2(n17050), .B1(n1750), .B2(n17051), .ZN(
        U729_Z_0) );
  OAI22_X1 U1726 ( .A1(n5338), .A2(n17050), .B1(n1810), .B2(n17052), .ZN(
        U728_Z_0) );
  OAI22_X1 U1727 ( .A1(n5305), .A2(n17045), .B1(n1808), .B2(n17046), .ZN(
        U727_Z_0) );
  OAI22_X1 U1728 ( .A1(n5306), .A2(n17045), .B1(n1807), .B2(n17046), .ZN(
        U726_Z_0) );
  OAI22_X1 U1729 ( .A1(n5307), .A2(n17045), .B1(n1809), .B2(n17046), .ZN(
        U725_Z_0) );
  OAI22_X1 U1730 ( .A1(n5308), .A2(n17045), .B1(n1750), .B2(n17046), .ZN(
        U724_Z_0) );
  OAI22_X1 U1731 ( .A1(n5309), .A2(n17045), .B1(n1810), .B2(n17047), .ZN(
        U723_Z_0) );
  OAI22_X1 U1732 ( .A1(n5284), .A2(n17040), .B1(n1808), .B2(n17041), .ZN(
        U722_Z_0) );
  OAI22_X1 U1733 ( .A1(n5285), .A2(n17040), .B1(n1807), .B2(n17041), .ZN(
        U721_Z_0) );
  OAI22_X1 U1734 ( .A1(n5286), .A2(n17040), .B1(n1809), .B2(n17041), .ZN(
        U720_Z_0) );
  OAI22_X1 U1735 ( .A1(n5287), .A2(n17040), .B1(n1750), .B2(n17041), .ZN(
        U719_Z_0) );
  OAI22_X1 U1736 ( .A1(n5288), .A2(n17040), .B1(n1810), .B2(n17042), .ZN(
        U718_Z_0) );
  OAI22_X1 U1737 ( .A1(n5263), .A2(n17035), .B1(n1808), .B2(n17036), .ZN(
        U717_Z_0) );
  OAI22_X1 U1738 ( .A1(n5264), .A2(n17035), .B1(n1807), .B2(n17036), .ZN(
        U716_Z_0) );
  OAI22_X1 U1739 ( .A1(n5265), .A2(n17035), .B1(n1809), .B2(n17036), .ZN(
        U715_Z_0) );
  OAI22_X1 U1740 ( .A1(n5266), .A2(n17035), .B1(n1750), .B2(n17036), .ZN(
        U714_Z_0) );
  OAI22_X1 U1741 ( .A1(n5267), .A2(n17035), .B1(n1810), .B2(n17037), .ZN(
        U713_Z_0) );
  OAI22_X1 U1742 ( .A1(n4962), .A2(n17030), .B1(n1808), .B2(n17031), .ZN(
        U712_Z_0) );
  OAI22_X1 U1743 ( .A1(n4996), .A2(n17030), .B1(n1807), .B2(n17031), .ZN(
        U711_Z_0) );
  OAI22_X1 U1744 ( .A1(n5020), .A2(n17030), .B1(n1809), .B2(n17031), .ZN(
        U710_Z_0) );
  OAI22_X1 U1745 ( .A1(n4985), .A2(n17030), .B1(n1750), .B2(n17031), .ZN(
        U709_Z_0) );
  OAI22_X1 U1746 ( .A1(n5038), .A2(n17030), .B1(n1810), .B2(n17032), .ZN(
        U708_Z_0) );
  OAI22_X1 U1747 ( .A1(n5169), .A2(n17025), .B1(n1808), .B2(n17026), .ZN(
        U707_Z_0) );
  OAI22_X1 U1748 ( .A1(n5170), .A2(n17025), .B1(n1807), .B2(n17026), .ZN(
        U706_Z_0) );
  OAI22_X1 U1749 ( .A1(n5171), .A2(n17025), .B1(n1809), .B2(n17026), .ZN(
        U705_Z_0) );
  OAI22_X1 U1750 ( .A1(n5172), .A2(n17025), .B1(n1750), .B2(n17026), .ZN(
        U704_Z_0) );
  OAI22_X1 U1751 ( .A1(n5173), .A2(n17025), .B1(n1810), .B2(n17027), .ZN(
        U703_Z_0) );
  OAI22_X1 U1752 ( .A1(n4979), .A2(n17020), .B1(n1808), .B2(n17021), .ZN(
        U702_Z_0) );
  OAI22_X1 U1753 ( .A1(n4995), .A2(n17020), .B1(n1807), .B2(n17021), .ZN(
        U701_Z_0) );
  OAI22_X1 U1754 ( .A1(n5019), .A2(n17020), .B1(n1809), .B2(n17021), .ZN(
        U700_Z_0) );
  OAI22_X1 U1755 ( .A1(n4984), .A2(n17020), .B1(n1750), .B2(n17021), .ZN(
        U699_Z_0) );
  OAI22_X1 U1756 ( .A1(n5037), .A2(n17020), .B1(n1810), .B2(n17022), .ZN(
        U698_Z_0) );
  OAI22_X1 U1757 ( .A1(n5198), .A2(n17015), .B1(n1808), .B2(n17016), .ZN(
        U697_Z_0) );
  OAI22_X1 U1758 ( .A1(n5199), .A2(n17015), .B1(n1807), .B2(n17016), .ZN(
        U696_Z_0) );
  OAI22_X1 U1759 ( .A1(n5200), .A2(n17015), .B1(n1809), .B2(n17016), .ZN(
        U695_Z_0) );
  OAI22_X1 U1760 ( .A1(n5201), .A2(n17015), .B1(n1750), .B2(n17016), .ZN(
        U694_Z_0) );
  INV_X1 U1762 ( .A(n190), .ZN(n179) );
  AOI221_X1 U1763 ( .B1(n2002), .B2(n2003), .C1(n2004), .C2(n2005), .A(n2006), 
        .ZN(n190) );
  INV_X1 U1764 ( .A(n2007), .ZN(n2006) );
  AOI221_X1 U1765 ( .B1(n2008), .B2(n2009), .C1(n2010), .C2(n2011), .A(n2012), 
        .ZN(n2007) );
  OAI22_X1 U1766 ( .A1(n5202), .A2(n17015), .B1(n1810), .B2(n17017), .ZN(
        U693_Z_0) );
  AOI22_X1 U1768 ( .A1(add_2073_SUM_1_), .A2(n17011), .B1(n17008), .B2(n1354), 
        .ZN(n2014) );
  INV_X1 U1769 ( .A(n2017), .ZN(n2013) );
  AOI221_X1 U1770 ( .B1(n2004), .B2(n2018), .C1(n2002), .C2(n2019), .A(n2020), 
        .ZN(n192) );
  INV_X1 U1771 ( .A(n2021), .ZN(n2020) );
  AOI221_X1 U1772 ( .B1(n2008), .B2(n2022), .C1(n2023), .C2(n2011), .A(n2012), 
        .ZN(n2021) );
  OAI22_X1 U1773 ( .A1(n5055), .A2(n2024), .B1(n2025), .B2(n2026), .ZN(
        U692_Z_0) );
  AOI22_X1 U1774 ( .A1(n2027), .A2(n2028), .B1(vis_pc_o[1]), .B2(n2029), .ZN(
        n2025) );
  INV_X1 U1777 ( .A(n2026), .ZN(n2024) );
  NAND2_X1 U1778 ( .A1(n17124), .A2(n2030), .ZN(n2026) );
  NAND3_X1 U1779 ( .A1(n753), .A2(n200), .A3(n2031), .ZN(n2030) );
  NAND4_X1 U1780 ( .A1(n2032), .A2(n2027), .A3(n16671), .A4(n16656), .ZN(n2031) );
  OAI22_X1 U1781 ( .A1(n4968), .A2(n2033), .B1(n2034), .B2(n2035), .ZN(
        U691_Z_0) );
  AOI21_X1 U1782 ( .B1(n2036), .B2(n2037), .A(n2038), .ZN(n2034) );
  OAI33_X1 U1783 ( .A1(n851), .A2(n4967), .A3(n16847), .B1(n2039), .B2(n5026), 
        .B3(n16794), .ZN(n2038) );
  NAND2_X1 U1784 ( .A1(n4967), .A2(n855), .ZN(n2039) );
  INV_X1 U1785 ( .A(n1178), .ZN(n855) );
  NAND2_X1 U1786 ( .A1(n527), .A2(n16849), .ZN(n1178) );
  OAI21_X1 U1787 ( .B1(n5233), .B2(n753), .A(n5055), .ZN(n2037) );
  OAI221_X1 U1788 ( .B1(n16847), .B2(n640), .C1(n16829), .C2(n16734), .A(n2040), .ZN(n2036) );
  NOR3_X1 U1789 ( .A1(n2041), .A2(n2042), .A3(n799), .ZN(n2040) );
  AOI21_X1 U1790 ( .B1(n451), .B2(n17096), .A(n16851), .ZN(n2041) );
  INV_X1 U1791 ( .A(n2035), .ZN(n2033) );
  OAI21_X1 U1792 ( .B1(n2043), .B2(n2044), .A(n17125), .ZN(n2035) );
  OAI221_X1 U1793 ( .B1(n1023), .B2(n522), .C1(n1857), .C2(n713), .A(n2045), 
        .ZN(n2044) );
  AOI22_X1 U1794 ( .A1(n785), .A2(n565), .B1(n534), .B2(n528), .ZN(n2045) );
  INV_X1 U1795 ( .A(n1230), .ZN(n534) );
  NAND2_X1 U1796 ( .A1(n528), .A2(n16849), .ZN(n522) );
  NAND4_X1 U1797 ( .A1(n2046), .A2(n738), .A3(n2047), .A4(n2048), .ZN(n2043)
         );
  AOI22_X1 U1798 ( .A1(n546), .A2(n17097), .B1(n1472), .B2(n16734), .ZN(n2048)
         );
  NOR2_X1 U1799 ( .A1(n594), .A2(n17096), .ZN(n1472) );
  NOR2_X1 U1800 ( .A1(n1217), .A2(n16859), .ZN(n546) );
  NAND3_X1 U1801 ( .A1(n527), .A2(n16824), .A3(n728), .ZN(n2047) );
  NAND3_X1 U1802 ( .A1(n1097), .A2(n1574), .A3(n2049), .ZN(n2046) );
  OAI22_X1 U1803 ( .A1(n5260), .A2(n17003), .B1(n1809), .B2(n17004), .ZN(
        U687_Z_0) );
  OAI22_X1 U1804 ( .A1(n5261), .A2(n17003), .B1(n1807), .B2(n17004), .ZN(
        U686_Z_0) );
  OAI22_X1 U1805 ( .A1(n5262), .A2(n17003), .B1(n1808), .B2(n17005), .ZN(
        U685_Z_0) );
  OAI22_X1 U1806 ( .A1(n5018), .A2(n16998), .B1(n1809), .B2(n16999), .ZN(
        U684_Z_0) );
  INV_X1 U1808 ( .A(n39), .ZN(n2056) );
  AOI221_X1 U1809 ( .B1(n2057), .B2(n2008), .C1(n2058), .C2(n2002), .A(n2059), 
        .ZN(n39) );
  INV_X1 U1810 ( .A(n2060), .ZN(n2059) );
  AOI221_X1 U1811 ( .B1(n2011), .B2(n2061), .C1(n2004), .C2(n2062), .A(n2012), 
        .ZN(n2060) );
  OAI22_X1 U1812 ( .A1(n4994), .A2(n16998), .B1(n1807), .B2(n16999), .ZN(
        U683_Z_0) );
  AOI221_X1 U1814 ( .B1(n2066), .B2(n2067), .C1(n2068), .C2(n2069), .A(n2070), 
        .ZN(n76) );
  INV_X1 U1815 ( .A(n2071), .ZN(n2070) );
  AOI221_X1 U1816 ( .B1(n2072), .B2(n2073), .C1(n2074), .C2(n2075), .A(n2076), 
        .ZN(n2071) );
  OAI22_X1 U1817 ( .A1(n4969), .A2(n16998), .B1(n1808), .B2(n17000), .ZN(
        U682_Z_0) );
  OAI22_X1 U1819 ( .A1(n5643), .A2(n17003), .B1(n2079), .B2(n17005), .ZN(
        U681_Z_0) );
  OAI22_X1 U1820 ( .A1(n5642), .A2(n16998), .B1(n2079), .B2(n17000), .ZN(
        U680_Z_0) );
  OAI22_X1 U1821 ( .A1(n5641), .A2(n17040), .B1(n2079), .B2(n17042), .ZN(
        U679_Z_0) );
  OAI22_X1 U1822 ( .A1(n5640), .A2(n17035), .B1(n2079), .B2(n17037), .ZN(
        U678_Z_0) );
  OAI22_X1 U1823 ( .A1(n5082), .A2(n17030), .B1(n2079), .B2(n17032), .ZN(
        U677_Z_0) );
  OAI22_X1 U1824 ( .A1(n5174), .A2(n17025), .B1(n2079), .B2(n17027), .ZN(
        U676_Z_0) );
  OAI22_X1 U1825 ( .A1(n5081), .A2(n17020), .B1(n2079), .B2(n17022), .ZN(
        U675_Z_0) );
  OAI22_X1 U1826 ( .A1(n5203), .A2(n17015), .B1(n2079), .B2(n17017), .ZN(
        U674_Z_0) );
  OAI22_X1 U1827 ( .A1(n5310), .A2(n17045), .B1(n2079), .B2(n17047), .ZN(
        U673_Z_0) );
  OAI22_X1 U1828 ( .A1(n5339), .A2(n17050), .B1(n2079), .B2(n17052), .ZN(
        U672_Z_0) );
  OAI22_X1 U1829 ( .A1(n5368), .A2(n17055), .B1(n2079), .B2(n17057), .ZN(
        U671_Z_0) );
  OAI22_X1 U1830 ( .A1(n5397), .A2(n17060), .B1(n2079), .B2(n17062), .ZN(
        U670_Z_0) );
  OAI22_X1 U1831 ( .A1(n5426), .A2(n17065), .B1(n2079), .B2(n17067), .ZN(
        U669_Z_0) );
  OAI22_X1 U1832 ( .A1(n5455), .A2(n17070), .B1(n2079), .B2(n17072), .ZN(
        U668_Z_0) );
  OAI22_X1 U1833 ( .A1(n5080), .A2(n17075), .B1(n2079), .B2(n17077), .ZN(
        U667_Z_0) );
  OAI22_X1 U1834 ( .A1(n5479), .A2(n17080), .B1(n2079), .B2(n17082), .ZN(
        U666_Z_0) );
  INV_X1 U1836 ( .A(n2082), .ZN(n2081) );
  AOI221_X1 U1837 ( .B1(n17006), .B2(n2083), .C1(add_2073_SUM_31_), .C2(n17010), .A(n2084), .ZN(n2082) );
  OAI22_X1 U1838 ( .A1(n4954), .A2(n2085), .B1(n2086), .B2(n2087), .ZN(
        U665_Z_0) );
  AOI222_X1 U1839 ( .A1(n88), .A2(n2083), .B1(n1528), .B2(n84), .C1(n86), .C2(
        n117), .ZN(n2086) );
  OAI221_X1 U1840 ( .B1(n2088), .B2(n2089), .C1(n2090), .C2(n2091), .A(n2092), 
        .ZN(n117) );
  AOI221_X1 U1841 ( .B1(n2074), .B2(n2093), .C1(n2067), .C2(n2094), .A(n2076), 
        .ZN(n2092) );
  INV_X1 U1842 ( .A(n2095), .ZN(n1528) );
  OAI22_X1 U1843 ( .A1(n4947), .A2(n2096), .B1(n2097), .B2(n1759), .ZN(n2095)
         );
  NOR4_X1 U1844 ( .A1(n2098), .A2(n2099), .A3(n2100), .A4(n2101), .ZN(n2097)
         );
  NAND4_X1 U1845 ( .A1(n2102), .A2(n2103), .A3(n2104), .A4(n2105), .ZN(n2101)
         );
  AND4_X1 U1846 ( .A1(n2106), .A2(n2107), .A3(n2108), .A4(n2109), .ZN(n2105)
         );
  INV_X1 U1847 ( .A(n2110), .ZN(n2108) );
  AND2_X1 U1848 ( .A1(n2111), .A2(n2112), .ZN(n2106) );
  AND3_X1 U1849 ( .A1(n2113), .A2(n2114), .A3(n2115), .ZN(n2104) );
  NAND4_X1 U1850 ( .A1(n2116), .A2(n2063), .A3(n2117), .A4(n2118), .ZN(n2100)
         );
  AOI211_X1 U1851 ( .C1(n16995), .C2(n2120), .A(n2121), .B(n2080), .ZN(n2118)
         );
  OAI221_X1 U1852 ( .B1(n1677), .B2(n2122), .C1(n4954), .C2(n2123), .A(n2124), 
        .ZN(n2080) );
  INV_X1 U1853 ( .A(n2125), .ZN(n2123) );
  AOI22_X1 U1854 ( .A1(U180_Z_0), .A2(n2126), .B1(n2127), .B2(n2128), .ZN(
        n2122) );
  INV_X1 U1855 ( .A(U180_Z_0), .ZN(n2128) );
  OAI221_X1 U1856 ( .B1(n16992), .B2(n2130), .C1(n2131), .C2(n2132), .A(n2133), 
        .ZN(n2121) );
  OAI21_X1 U1857 ( .B1(n2134), .B2(n2135), .A(n17011), .ZN(n2133) );
  NAND4_X1 U1858 ( .A1(n2136), .A2(n2137), .A3(n2138), .A4(n2139), .ZN(n2135)
         );
  NOR4_X1 U1859 ( .A1(n16658), .A2(n16679), .A3(n16653), .A4(n16719), .ZN(
        n2139) );
  NOR3_X1 U1860 ( .A1(n16710), .A2(add_2073_SUM_1_), .A3(n16672), .ZN(n2138)
         );
  INV_X1 U1861 ( .A(n16711), .ZN(n2137) );
  INV_X1 U1862 ( .A(n16715), .ZN(n2136) );
  NAND4_X1 U1863 ( .A1(n1655), .A2(n2140), .A3(n2141), .A4(n2142), .ZN(n2134)
         );
  NOR3_X1 U1864 ( .A1(n2143), .A2(add_2073_SUM_31_), .A3(n16663), .ZN(n2142)
         );
  OR3_X1 U1865 ( .A1(add_2073_SUM_7_), .A2(n16722), .A3(n16682), .ZN(n2143) );
  NOR3_X1 U1866 ( .A1(n16668), .A2(n16655), .A3(n16702), .ZN(n2141) );
  INV_X1 U1867 ( .A(n16706), .ZN(n2140) );
  INV_X1 U1868 ( .A(n16709), .ZN(n1655) );
  AOI211_X1 U1869 ( .C1(n5818), .C2(n2144), .A(n2145), .B(n2146), .ZN(n2132)
         );
  INV_X1 U1870 ( .A(n2147), .ZN(n2146) );
  AOI22_X1 U1871 ( .A1(n2148), .A2(n5819), .B1(n1665), .B2(n5807), .ZN(n2147)
         );
  OAI221_X1 U1872 ( .B1(n1654), .B2(n2149), .C1(n1691), .C2(n2150), .A(n2151), 
        .ZN(n2145) );
  AOI22_X1 U1873 ( .A1(n4952), .A2(n1645), .B1(n5815), .B2(n1651), .ZN(n2151)
         );
  AOI211_X1 U1874 ( .C1(n2152), .C2(n2144), .A(n2153), .B(n2154), .ZN(n2130)
         );
  OAI22_X1 U1875 ( .A1(n1625), .A2(n5819), .B1(n1694), .B2(n5807), .ZN(n2154)
         );
  OAI221_X1 U1876 ( .B1(n1682), .B2(n4952), .C1(n1687), .C2(n5815), .A(n2155), 
        .ZN(n2153) );
  AOI22_X1 U1877 ( .A1(n2149), .A2(n2156), .B1(n2150), .B2(n1658), .ZN(n2155)
         );
  INV_X1 U1878 ( .A(n5811), .ZN(n2150) );
  INV_X1 U1879 ( .A(n5813), .ZN(n2149) );
  INV_X1 U1880 ( .A(n5818), .ZN(n2152) );
  NAND4_X1 U1881 ( .A1(n2157), .A2(n2158), .A3(n2159), .A4(n2160), .ZN(n2120)
         );
  AOI222_X1 U1882 ( .A1(n1686), .A2(n5816), .B1(n1682), .B2(n4952), .C1(n1630), 
        .C2(n5817), .ZN(n2160) );
  INV_X1 U1883 ( .A(n2161), .ZN(n1630) );
  AOI222_X1 U1884 ( .A1(n1654), .A2(n5813), .B1(n1687), .B2(n5815), .C1(n1688), 
        .C2(n5814), .ZN(n2159) );
  AOI222_X1 U1885 ( .A1(n1692), .A2(n5810), .B1(n1690), .B2(n5812), .C1(n1691), 
        .C2(n5811), .ZN(n2158) );
  AOI222_X1 U1886 ( .A1(n1661), .A2(n5818), .B1(n1694), .B2(n5807), .C1(n1625), 
        .C2(n5819), .ZN(n2157) );
  NOR3_X1 U1887 ( .A1(n2001), .A2(n2054), .A3(n2017), .ZN(n2117) );
  OAI221_X1 U1888 ( .B1(n2162), .B2(n2163), .C1(n186), .C2(n2164), .A(n2165), 
        .ZN(n2017) );
  NOR3_X1 U1889 ( .A1(n2166), .A2(n2055), .A3(n2167), .ZN(n2165) );
  NOR4_X1 U1890 ( .A1(n16810), .A2(n16656), .A3(n1045), .A4(n2168), .ZN(n2167)
         );
  NOR3_X1 U1891 ( .A1(add_2082_B_1_), .A2(n16992), .A3(n1689), .ZN(n2166) );
  INV_X1 U1892 ( .A(add_2082_B_1_), .ZN(n2163) );
  XOR2_X1 U1893 ( .A(n2169), .B(n2170), .Z(add_2082_B_1_) );
  AOI22_X1 U1894 ( .A1(n16988), .A2(n1354), .B1(n2172), .B2(n2173), .ZN(n2170)
         );
  AOI22_X1 U1895 ( .A1(n1689), .A2(n16995), .B1(n2174), .B2(n2126), .ZN(n2162)
         );
  INV_X1 U1896 ( .A(n2174), .ZN(n1689) );
  NAND2_X1 U1897 ( .A1(n2175), .A2(n2176), .ZN(n2174) );
  AOI221_X1 U1898 ( .B1(n16985), .B2(vis_r11_o[0]), .C1(n16984), .C2(
        vis_r14_o[0]), .A(n2181), .ZN(n2176) );
  OAI22_X1 U1899 ( .A1(n5267), .A2(n2182), .B1(n2183), .B2(n2184), .ZN(n2181)
         );
  AOI221_X1 U1901 ( .B1(n16979), .B2(vis_r9_o[0]), .C1(n16976), .C2(n2188), 
        .A(n2189), .ZN(n2175) );
  OAI22_X1 U1902 ( .A1(n5396), .A2(n2190), .B1(n5338), .B2(n2191), .ZN(n2189)
         );
  OAI211_X1 U1903 ( .C1(n2192), .C2(n2193), .A(n2194), .B(n2195), .ZN(n2054)
         );
  AOI22_X1 U1904 ( .A1(n17008), .A2(n2196), .B1(n16726), .B2(n17011), .ZN(
        n2195) );
  NAND3_X1 U1905 ( .A1(n1627), .A2(n2127), .A3(n2193), .ZN(n2194) );
  INV_X1 U1906 ( .A(n5821), .ZN(n2193) );
  XOR2_X1 U1907 ( .A(n16990), .B(n2197), .Z(n5821) );
  AOI221_X1 U1908 ( .B1(n2198), .B2(n16674), .C1(n16988), .C2(n2196), .A(n2199), .ZN(n2197) );
  OAI22_X1 U1909 ( .A1(n5256), .A2(n2200), .B1(n5258), .B2(n2201), .ZN(n2199)
         );
  AOI22_X1 U1910 ( .A1(n1672), .A2(n16995), .B1(n1627), .B2(n2126), .ZN(n2192)
         );
  INV_X1 U1911 ( .A(n1627), .ZN(n1672) );
  NAND4_X1 U1912 ( .A1(n2202), .A2(n2203), .A3(n2204), .A4(n2205), .ZN(n1627)
         );
  AOI222_X1 U1913 ( .A1(n16973), .A2(vis_msp_o[5]), .B1(n16972), .B2(n2209), 
        .C1(n16968), .C2(vis_psp_o[5]), .ZN(n2205) );
  AOI222_X1 U1914 ( .A1(n16982), .A2(vis_r14_o[7]), .B1(n16964), .B2(
        vis_r12_o[7]), .C1(n16985), .C2(vis_r11_o[7]), .ZN(n2204) );
  AOI222_X1 U1915 ( .A1(n16979), .A2(vis_r9_o[7]), .B1(n16962), .B2(
        vis_r10_o[7]), .C1(n16959), .C2(vis_r8_o[7]), .ZN(n2203) );
  AOI22_X1 U1916 ( .A1(n16976), .A2(n2221), .B1(n16955), .B2(n1152), .ZN(n2202) );
  OAI211_X1 U1917 ( .C1(n2223), .C2(n2224), .A(n2225), .B(n2226), .ZN(n2001)
         );
  AOI222_X1 U1918 ( .A1(n16732), .A2(n17009), .B1(n2227), .B2(vis_ipsr_o[1]), 
        .C1(n17007), .C2(n2028), .ZN(n2226) );
  AOI21_X1 U1919 ( .B1(n2228), .B2(n2224), .A(n2229), .ZN(n2225) );
  NOR4_X1 U1920 ( .A1(n16809), .A2(n5055), .A3(n16810), .A4(n2168), .ZN(n2229)
         );
  NOR2_X1 U1921 ( .A1(n16992), .A2(n1679), .ZN(n2228) );
  INV_X1 U1922 ( .A(n5822), .ZN(n2224) );
  XOR2_X1 U1923 ( .A(n16990), .B(n2230), .Z(n5822) );
  AOI222_X1 U1924 ( .A1(n16988), .A2(n2028), .B1(n2198), .B2(n451), .C1(n2231), 
        .C2(n2173), .ZN(n2230) );
  AOI22_X1 U1925 ( .A1(n1679), .A2(n16994), .B1(n2232), .B2(n2126), .ZN(n2223)
         );
  INV_X1 U1926 ( .A(n2232), .ZN(n1679) );
  AOI221_X1 U1927 ( .B1(n89), .B2(n17006), .C1(vis_apsr_o[0]), .C2(n2125), .A(
        n2055), .ZN(n2063) );
  INV_X1 U1928 ( .A(n2233), .ZN(n2116) );
  NAND4_X1 U1929 ( .A1(n2234), .A2(n2235), .A3(n2236), .A4(n2237), .ZN(n2099)
         );
  NOR3_X1 U1930 ( .A1(n2238), .A2(n2239), .A3(n2240), .ZN(n2237) );
  AOI21_X1 U1931 ( .B1(n2241), .B2(n2242), .A(n2243), .ZN(n2240) );
  NOR4_X1 U1932 ( .A1(n2244), .A2(n2245), .A3(n2246), .A4(n2247), .ZN(n2242)
         );
  OR3_X1 U1933 ( .A1(n2083), .A2(n2248), .A3(n2249), .ZN(n2245) );
  OR4_X1 U1934 ( .A1(n2250), .A2(n2251), .A3(n17), .A4(n2252), .ZN(n2244) );
  OR2_X1 U1935 ( .A1(n2253), .A2(n2254), .ZN(n2252) );
  NOR4_X1 U1936 ( .A1(n2255), .A2(n2256), .A3(n2257), .A4(n2258), .ZN(n2241)
         );
  OR3_X1 U1937 ( .A1(n22), .A2(n20), .A3(n21), .ZN(n2256) );
  OR4_X1 U1938 ( .A1(n2259), .A2(n2260), .A3(n1354), .A4(n2261), .ZN(n2255) );
  INV_X1 U1939 ( .A(n2064), .ZN(n2239) );
  NAND2_X1 U1940 ( .A1(n16695), .A2(n17011), .ZN(n2064) );
  NAND3_X1 U1941 ( .A1(n2262), .A2(n2065), .A3(n2263), .ZN(n2238) );
  OAI221_X1 U1942 ( .B1(U189_Z_0), .B2(n2264), .C1(n16995), .C2(n1832), .A(
        n2265), .ZN(n2065) );
  NAND3_X1 U1943 ( .A1(U189_Z_0), .A2(n1832), .A3(n2131), .ZN(n2265) );
  NOR2_X1 U1944 ( .A1(n1680), .A2(n16993), .ZN(n2264) );
  INV_X1 U1945 ( .A(n1832), .ZN(n1680) );
  NAND4_X1 U1946 ( .A1(n2266), .A2(n2267), .A3(n2268), .A4(n2269), .ZN(n1832)
         );
  AOI222_X1 U1947 ( .A1(n16973), .A2(vis_msp_o[26]), .B1(n16972), .B2(n2271), 
        .C1(n16967), .C2(vis_psp_o[26]), .ZN(n2269) );
  AOI222_X1 U1949 ( .A1(n16982), .A2(vis_r14_o[28]), .B1(n16964), .B2(
        vis_r12_o[28]), .C1(n16985), .C2(vis_r11_o[28]), .ZN(n2268) );
  AOI222_X1 U1952 ( .A1(n16979), .A2(vis_r9_o[28]), .B1(n16961), .B2(
        vis_r10_o[28]), .C1(n16958), .C2(vis_r8_o[28]), .ZN(n2267) );
  AOI22_X1 U1954 ( .A1(n16976), .A2(n2279), .B1(n16954), .B2(n2280), .ZN(n2266) );
  AND3_X1 U1955 ( .A1(n2281), .A2(n2282), .A3(n2283), .ZN(n2236) );
  NAND4_X1 U1956 ( .A1(n2284), .A2(n2285), .A3(n2286), .A4(n2287), .ZN(n2098)
         );
  NOR4_X1 U1957 ( .A1(n2288), .A2(n2084), .A3(n2289), .A4(n2290), .ZN(n2287)
         );
  INV_X1 U1958 ( .A(n2291), .ZN(n2290) );
  AND3_X1 U1959 ( .A1(n16995), .A2(U180_Z_0), .A3(n1677), .ZN(n2084) );
  AND4_X1 U1960 ( .A1(n2292), .A2(n2293), .A3(n2294), .A4(n2295), .ZN(n1677)
         );
  AOI222_X1 U1961 ( .A1(n16973), .A2(vis_msp_o[28]), .B1(n16972), .B2(n2297), 
        .C1(n16967), .C2(vis_psp_o[28]), .ZN(n2295) );
  AOI222_X1 U1963 ( .A1(n16982), .A2(vis_r14_o[30]), .B1(n16965), .B2(
        vis_r12_o[30]), .C1(n16985), .C2(vis_r11_o[30]), .ZN(n2294) );
  AOI222_X1 U1966 ( .A1(n16979), .A2(vis_r9_o[30]), .B1(n16961), .B2(
        vis_r10_o[30]), .C1(n16958), .C2(vis_r8_o[30]), .ZN(n2293) );
  AOI22_X1 U1968 ( .A1(n16976), .A2(n874), .B1(n16954), .B2(n881), .ZN(n2292)
         );
  NAND3_X1 U1969 ( .A1(n2305), .A2(n2306), .A3(n2307), .ZN(n2288) );
  NOR3_X1 U1970 ( .A1(n2308), .A2(n2309), .A3(n2310), .ZN(n2286) );
  AOI221_X1 U1971 ( .B1(n2311), .B2(n2312), .C1(n2313), .C2(n2314), .A(n2315), 
        .ZN(n2096) );
  OAI221_X1 U1972 ( .B1(n2316), .B2(n2317), .C1(n2318), .C2(n2319), .A(n2320), 
        .ZN(n2315) );
  OAI33_X1 U1973 ( .A1(n2321), .A2(n2322), .A3(n2323), .B1(n2324), .B2(n2325), 
        .B3(n2326), .ZN(n2320) );
  NAND3_X1 U1974 ( .A1(n1781), .A2(n1789), .A3(n2327), .ZN(n2324) );
  OAI33_X1 U1975 ( .A1(n2328), .A2(n2329), .A3(n2330), .B1(n2331), .B2(n2332), 
        .B3(n2333), .ZN(n2327) );
  OR3_X1 U1976 ( .A1(n2334), .A2(n16788), .A3(n2336), .ZN(n2331) );
  OR3_X1 U1977 ( .A1(n2337), .A2(n2338), .A3(n2339), .ZN(n2328) );
  AOI21_X1 U1978 ( .B1(n2340), .B2(n2341), .A(n2342), .ZN(n2319) );
  NOR3_X1 U1979 ( .A1(n2343), .A2(n2344), .A3(n2345), .ZN(n2318) );
  NAND3_X1 U1980 ( .A1(n1779), .A2(n2346), .A3(n2347), .ZN(n2343) );
  OAI33_X1 U1981 ( .A1(n2348), .A2(n2349), .A3(n2350), .B1(n2351), .B2(n2352), 
        .B3(n2353), .ZN(n2347) );
  OR3_X1 U1982 ( .A1(n2354), .A2(n16789), .A3(n2355), .ZN(n2351) );
  OR3_X1 U1983 ( .A1(n2337), .A2(n2356), .A3(n2357), .ZN(n2348) );
  NOR4_X1 U1984 ( .A1(n2358), .A2(n2340), .A3(n2359), .A4(n2360), .ZN(n2317)
         );
  NOR4_X1 U1985 ( .A1(n2361), .A2(n2362), .A3(n2363), .A4(n2364), .ZN(n2316)
         );
  OAI22_X1 U1986 ( .A1(n2365), .A2(n2366), .B1(n2367), .B2(n2368), .ZN(n2362)
         );
  NOR2_X1 U1987 ( .A1(n2337), .A2(n2369), .ZN(n2367) );
  INV_X1 U1988 ( .A(n2370), .ZN(n2366) );
  INV_X1 U1989 ( .A(n2371), .ZN(n2365) );
  NAND4_X1 U1990 ( .A1(n2372), .A2(n2373), .A3(n2374), .A4(n2375), .ZN(n2361)
         );
  OAI21_X1 U1991 ( .B1(n2340), .B2(n2342), .A(n2376), .ZN(n2314) );
  INV_X1 U1992 ( .A(n2377), .ZN(n2342) );
  NAND4_X1 U1993 ( .A1(n2378), .A2(n2379), .A3(n2380), .A4(n2381), .ZN(n2312)
         );
  OAI33_X1 U1994 ( .A1(n2382), .A2(n2329), .A3(n2330), .B1(n2383), .B2(n2352), 
        .B3(n2353), .ZN(n2381) );
  OR3_X1 U1995 ( .A1(n2337), .A2(n2384), .A3(n2385), .ZN(n2383) );
  OR3_X1 U1996 ( .A1(n2386), .A2(n16789), .A3(n2387), .ZN(n2382) );
  AND2_X1 U1997 ( .A1(n1791), .A2(n1772), .ZN(n2380) );
  INV_X1 U1998 ( .A(n2388), .ZN(n2379) );
  OAI21_X1 U1999 ( .B1(n2389), .B2(n2390), .A(n2377), .ZN(n2311) );
  OAI22_X1 U2000 ( .A1(n5079), .A2(n17003), .B1(n2391), .B2(n17005), .ZN(
        U664_Z_0) );
  OAI22_X1 U2001 ( .A1(n5078), .A2(n16998), .B1(n2391), .B2(n17000), .ZN(
        U663_Z_0) );
  OAI22_X1 U2002 ( .A1(n5289), .A2(n17040), .B1(n2391), .B2(n17042), .ZN(
        U662_Z_0) );
  OAI22_X1 U2003 ( .A1(n5268), .A2(n17035), .B1(n2391), .B2(n17037), .ZN(
        U661_Z_0) );
  OAI22_X1 U2004 ( .A1(n5077), .A2(n17030), .B1(n2391), .B2(n17032), .ZN(
        U660_Z_0) );
  OAI22_X1 U2005 ( .A1(n5175), .A2(n17025), .B1(n2391), .B2(n17027), .ZN(
        U659_Z_0) );
  OAI22_X1 U2006 ( .A1(n5076), .A2(n17020), .B1(n2391), .B2(n17022), .ZN(
        U658_Z_0) );
  OAI22_X1 U2007 ( .A1(n5204), .A2(n17015), .B1(n2391), .B2(n17017), .ZN(
        U657_Z_0) );
  OAI22_X1 U2008 ( .A1(n5311), .A2(n17045), .B1(n2391), .B2(n17047), .ZN(
        U656_Z_0) );
  OAI22_X1 U2009 ( .A1(n5340), .A2(n17050), .B1(n2391), .B2(n17052), .ZN(
        U655_Z_0) );
  OAI22_X1 U2010 ( .A1(n5369), .A2(n17055), .B1(n2391), .B2(n17057), .ZN(
        U654_Z_0) );
  OAI22_X1 U2011 ( .A1(n5398), .A2(n17060), .B1(n2391), .B2(n17062), .ZN(
        U653_Z_0) );
  OAI22_X1 U2012 ( .A1(n5427), .A2(n17065), .B1(n2391), .B2(n17067), .ZN(
        U652_Z_0) );
  OAI22_X1 U2013 ( .A1(n5456), .A2(n17070), .B1(n2391), .B2(n17072), .ZN(
        U651_Z_0) );
  OAI22_X1 U2014 ( .A1(n5075), .A2(n17075), .B1(n2391), .B2(n17077), .ZN(
        U650_Z_0) );
  OAI22_X1 U2015 ( .A1(n5480), .A2(n17080), .B1(n2391), .B2(n17082), .ZN(
        U649_Z_0) );
  OAI211_X1 U2017 ( .C1(n2392), .C2(n2393), .A(n2394), .B(n2395), .ZN(n2233)
         );
  AOI222_X1 U2018 ( .A1(n2125), .A2(vis_apsr_o[1]), .B1(n17008), .B2(n1755), 
        .C1(n16693), .C2(n17009), .ZN(n2395) );
  AOI21_X1 U2020 ( .B1(n2396), .B2(n1870), .A(n2055), .ZN(n2394) );
  NOR2_X1 U2021 ( .A1(U158_Z_0), .A2(n16993), .ZN(n2396) );
  AOI22_X1 U2022 ( .A1(n1678), .A2(n16994), .B1(n1870), .B2(n2126), .ZN(n2393)
         );
  INV_X1 U2023 ( .A(n1870), .ZN(n1678) );
  NAND4_X1 U2024 ( .A1(n2397), .A2(n2398), .A3(n2399), .A4(n2400), .ZN(n1870)
         );
  AOI222_X1 U2025 ( .A1(n16974), .A2(vis_msp_o[27]), .B1(n16972), .B2(n2402), 
        .C1(n16967), .C2(vis_psp_o[27]), .ZN(n2400) );
  AOI222_X1 U2027 ( .A1(n16982), .A2(vis_r14_o[29]), .B1(n16965), .B2(
        vis_r12_o[29]), .C1(n16985), .C2(vis_r11_o[29]), .ZN(n2399) );
  AOI222_X1 U2030 ( .A1(n16979), .A2(vis_r9_o[29]), .B1(n16961), .B2(
        vis_r10_o[29]), .C1(n16958), .C2(vis_r8_o[29]), .ZN(n2398) );
  AOI22_X1 U2032 ( .A1(n16976), .A2(n881), .B1(n16954), .B2(n2279), .ZN(n2397)
         );
  INV_X1 U2035 ( .A(U158_Z_0), .ZN(n2392) );
  INV_X1 U2036 ( .A(n72), .ZN(n1754) );
  AOI221_X1 U2037 ( .B1(n2410), .B2(n2067), .C1(n2411), .C2(n2074), .A(n2412), 
        .ZN(n72) );
  INV_X1 U2038 ( .A(n2413), .ZN(n2412) );
  AOI221_X1 U2039 ( .B1(n2072), .B2(n2414), .C1(n2415), .C2(n2069), .A(n2076), 
        .ZN(n2413) );
  OAI22_X1 U2040 ( .A1(n5630), .A2(n17003), .B1(n2416), .B2(n17005), .ZN(
        U648_Z_0) );
  OAI22_X1 U2041 ( .A1(n5629), .A2(n16998), .B1(n2416), .B2(n17000), .ZN(
        U647_Z_0) );
  OAI22_X1 U2042 ( .A1(n5628), .A2(n17040), .B1(n2416), .B2(n17042), .ZN(
        U646_Z_0) );
  OAI22_X1 U2043 ( .A1(n5627), .A2(n17035), .B1(n2416), .B2(n17037), .ZN(
        U645_Z_0) );
  OAI22_X1 U2044 ( .A1(n5113), .A2(n17030), .B1(n2416), .B2(n17032), .ZN(
        U644_Z_0) );
  OAI22_X1 U2045 ( .A1(n5176), .A2(n17025), .B1(n2416), .B2(n17027), .ZN(
        U643_Z_0) );
  OAI22_X1 U2046 ( .A1(n5112), .A2(n17020), .B1(n2416), .B2(n17022), .ZN(
        U642_Z_0) );
  OAI22_X1 U2047 ( .A1(n5205), .A2(n17015), .B1(n2416), .B2(n17017), .ZN(
        U641_Z_0) );
  OAI22_X1 U2048 ( .A1(n5312), .A2(n17045), .B1(n2416), .B2(n17047), .ZN(
        U640_Z_0) );
  OAI22_X1 U2049 ( .A1(n5341), .A2(n17050), .B1(n2416), .B2(n17052), .ZN(
        U639_Z_0) );
  OAI22_X1 U2050 ( .A1(n5370), .A2(n17055), .B1(n2416), .B2(n17057), .ZN(
        U638_Z_0) );
  OAI22_X1 U2051 ( .A1(n5399), .A2(n17060), .B1(n2416), .B2(n17062), .ZN(
        U637_Z_0) );
  OAI22_X1 U2052 ( .A1(n5428), .A2(n17065), .B1(n2416), .B2(n17067), .ZN(
        U636_Z_0) );
  OAI22_X1 U2053 ( .A1(n5457), .A2(n17070), .B1(n2416), .B2(n17072), .ZN(
        U635_Z_0) );
  OAI22_X1 U2054 ( .A1(n5111), .A2(n17075), .B1(n2416), .B2(n17077), .ZN(
        U634_Z_0) );
  OAI22_X1 U2055 ( .A1(n5481), .A2(n17080), .B1(n2416), .B2(n17082), .ZN(
        U633_Z_0) );
  OAI221_X1 U2057 ( .B1(n2417), .B2(n2418), .C1(n2089), .C2(n2419), .A(n2420), 
        .ZN(n99) );
  AOI221_X1 U2058 ( .B1(n2074), .B2(n2421), .C1(n2422), .C2(n2069), .A(n2076), 
        .ZN(n2420) );
  OAI211_X1 U2059 ( .C1(n2423), .C2(n2424), .A(n2425), .B(n2426), .ZN(n2110)
         );
  AOI22_X1 U2060 ( .A1(n17008), .A2(n2427), .B1(n16698), .B2(n17010), .ZN(
        n2426) );
  NAND3_X1 U2061 ( .A1(n2127), .A2(n2423), .A3(n1644), .ZN(n2425) );
  AOI22_X1 U2062 ( .A1(n1681), .A2(n16994), .B1(n1644), .B2(n2126), .ZN(n2424)
         );
  INV_X1 U2063 ( .A(n1644), .ZN(n1681) );
  NAND4_X1 U2064 ( .A1(n2428), .A2(n2429), .A3(n2430), .A4(n2431), .ZN(n1644)
         );
  AOI222_X1 U2065 ( .A1(n16973), .A2(vis_msp_o[25]), .B1(n16972), .B2(n2433), 
        .C1(n16967), .C2(vis_psp_o[25]), .ZN(n2431) );
  AOI222_X1 U2067 ( .A1(n16982), .A2(vis_r14_o[27]), .B1(n16964), .B2(
        vis_r12_o[27]), .C1(n16985), .C2(vis_r11_o[27]), .ZN(n2430) );
  AOI222_X1 U2070 ( .A1(n16979), .A2(vis_r9_o[27]), .B1(n16961), .B2(
        vis_r10_o[27]), .C1(n16958), .C2(vis_r8_o[27]), .ZN(n2429) );
  AOI22_X1 U2072 ( .A1(n16976), .A2(n2280), .B1(n16954), .B2(n2441), .ZN(n2428) );
  INV_X1 U2074 ( .A(U175_Z_0), .ZN(n2423) );
  OAI22_X1 U2075 ( .A1(n4993), .A2(n17003), .B1(n2442), .B2(n17005), .ZN(
        U632_Z_0) );
  OAI22_X1 U2076 ( .A1(n4992), .A2(n16998), .B1(n2442), .B2(n17000), .ZN(
        U631_Z_0) );
  OAI22_X1 U2077 ( .A1(n5290), .A2(n17040), .B1(n2442), .B2(n17042), .ZN(
        U630_Z_0) );
  OAI22_X1 U2078 ( .A1(n5269), .A2(n17035), .B1(n2442), .B2(n17037), .ZN(
        U629_Z_0) );
  OAI22_X1 U2079 ( .A1(n4991), .A2(n17030), .B1(n2442), .B2(n17032), .ZN(
        U628_Z_0) );
  OAI22_X1 U2080 ( .A1(n5177), .A2(n17025), .B1(n2442), .B2(n17027), .ZN(
        U627_Z_0) );
  OAI22_X1 U2081 ( .A1(n4990), .A2(n17020), .B1(n2442), .B2(n17022), .ZN(
        U626_Z_0) );
  OAI22_X1 U2082 ( .A1(n5206), .A2(n17015), .B1(n2442), .B2(n17017), .ZN(
        U625_Z_0) );
  OAI22_X1 U2083 ( .A1(n5313), .A2(n17045), .B1(n2442), .B2(n17047), .ZN(
        U624_Z_0) );
  OAI22_X1 U2084 ( .A1(n5342), .A2(n17050), .B1(n2442), .B2(n17052), .ZN(
        U623_Z_0) );
  OAI22_X1 U2085 ( .A1(n5371), .A2(n17055), .B1(n2442), .B2(n17057), .ZN(
        U622_Z_0) );
  OAI22_X1 U2086 ( .A1(n5400), .A2(n17060), .B1(n2442), .B2(n17062), .ZN(
        U621_Z_0) );
  OAI22_X1 U2087 ( .A1(n5429), .A2(n17065), .B1(n2442), .B2(n17067), .ZN(
        U620_Z_0) );
  OAI22_X1 U2088 ( .A1(n5458), .A2(n17070), .B1(n2442), .B2(n17072), .ZN(
        U619_Z_0) );
  OAI22_X1 U2089 ( .A1(n4989), .A2(n17075), .B1(n2442), .B2(n17077), .ZN(
        U618_Z_0) );
  OAI22_X1 U2090 ( .A1(n5482), .A2(n17080), .B1(n2442), .B2(n17082), .ZN(
        U617_Z_0) );
  AOI221_X1 U2092 ( .B1(n17006), .B2(n2260), .C1(n16663), .C2(n17010), .A(
        n2055), .ZN(n2444) );
  OAI221_X1 U2093 ( .B1(n4952), .B2(n2445), .C1(n16995), .C2(n1645), .A(n2446), 
        .ZN(n2443) );
  NAND3_X1 U2094 ( .A1(n2131), .A2(n1645), .A3(n4952), .ZN(n2446) );
  NOR2_X1 U2095 ( .A1(n1682), .A2(n16993), .ZN(n2445) );
  INV_X1 U2096 ( .A(n1645), .ZN(n1682) );
  NAND4_X1 U2097 ( .A1(n2447), .A2(n2448), .A3(n2449), .A4(n2450), .ZN(n1645)
         );
  AOI222_X1 U2098 ( .A1(n16973), .A2(vis_msp_o[24]), .B1(n16972), .B2(n2452), 
        .C1(n16967), .C2(vis_psp_o[24]), .ZN(n2450) );
  AOI222_X1 U2100 ( .A1(n16982), .A2(vis_r14_o[26]), .B1(n16964), .B2(
        vis_r12_o[26]), .C1(n16985), .C2(vis_r11_o[26]), .ZN(n2449) );
  AOI222_X1 U2103 ( .A1(n16980), .A2(vis_r9_o[26]), .B1(n16961), .B2(
        vis_r10_o[26]), .C1(n16958), .C2(vis_r8_o[26]), .ZN(n2448) );
  AOI22_X1 U2105 ( .A1(n16976), .A2(n2441), .B1(n16954), .B2(n2460), .ZN(n2447) );
  INV_X1 U2108 ( .A(n2260), .ZN(n2463) );
  AOI221_X1 U2109 ( .B1(n2464), .B2(n2069), .C1(n2465), .C2(n2074), .A(n2466), 
        .ZN(n100) );
  INV_X1 U2110 ( .A(n2467), .ZN(n2466) );
  AOI221_X1 U2111 ( .B1(n2468), .B2(n2072), .C1(n2469), .C2(n2067), .A(n2076), 
        .ZN(n2467) );
  OAI22_X1 U2112 ( .A1(n5016), .A2(n17003), .B1(n2470), .B2(n17005), .ZN(
        U614_Z_0) );
  OAI22_X1 U2113 ( .A1(n5015), .A2(n16998), .B1(n2470), .B2(n17000), .ZN(
        U613_Z_0) );
  OAI22_X1 U2114 ( .A1(n5291), .A2(n17040), .B1(n2470), .B2(n17042), .ZN(
        U612_Z_0) );
  OAI22_X1 U2115 ( .A1(n5270), .A2(n17035), .B1(n2470), .B2(n17037), .ZN(
        U611_Z_0) );
  OAI22_X1 U2116 ( .A1(n5014), .A2(n17030), .B1(n2470), .B2(n17032), .ZN(
        U610_Z_0) );
  OAI22_X1 U2117 ( .A1(n5178), .A2(n17025), .B1(n2470), .B2(n17027), .ZN(
        U609_Z_0) );
  OAI22_X1 U2118 ( .A1(n5013), .A2(n17020), .B1(n2470), .B2(n17022), .ZN(
        U608_Z_0) );
  OAI22_X1 U2119 ( .A1(n5207), .A2(n17015), .B1(n2470), .B2(n17017), .ZN(
        U607_Z_0) );
  OAI22_X1 U2120 ( .A1(n5314), .A2(n17045), .B1(n2470), .B2(n17047), .ZN(
        U606_Z_0) );
  OAI22_X1 U2121 ( .A1(n5343), .A2(n17050), .B1(n2470), .B2(n17052), .ZN(
        U605_Z_0) );
  OAI22_X1 U2122 ( .A1(n5372), .A2(n17055), .B1(n2470), .B2(n17057), .ZN(
        U604_Z_0) );
  OAI22_X1 U2123 ( .A1(n5401), .A2(n17060), .B1(n2470), .B2(n17062), .ZN(
        U603_Z_0) );
  OAI22_X1 U2124 ( .A1(n5430), .A2(n17065), .B1(n2470), .B2(n17067), .ZN(
        U602_Z_0) );
  OAI22_X1 U2125 ( .A1(n5459), .A2(n17070), .B1(n2470), .B2(n17072), .ZN(
        U601_Z_0) );
  OAI22_X1 U2126 ( .A1(n5012), .A2(n17075), .B1(n2470), .B2(n17077), .ZN(
        U600_Z_0) );
  OAI22_X1 U2127 ( .A1(n5483), .A2(n17080), .B1(n2470), .B2(n17082), .ZN(
        U599_Z_0) );
  AOI221_X1 U2129 ( .B1(n16655), .B2(n17009), .C1(n17008), .C2(n2248), .A(n108), .ZN(n2471) );
  OAI221_X1 U2130 ( .B1(n2417), .B2(n2472), .C1(n2473), .C2(n2089), .A(n2474), 
        .ZN(n108) );
  AOI221_X1 U2131 ( .B1(n2074), .B2(n2003), .C1(n2005), .C2(n2069), .A(n2076), 
        .ZN(n2474) );
  NAND3_X1 U2132 ( .A1(n16995), .A2(n4951), .A3(n1683), .ZN(n2234) );
  INV_X1 U2133 ( .A(n1647), .ZN(n1683) );
  NAND2_X1 U2134 ( .A1(n2475), .A2(n1647), .ZN(n2291) );
  NAND4_X1 U2135 ( .A1(n2476), .A2(n2477), .A3(n2478), .A4(n2479), .ZN(n1647)
         );
  AOI222_X1 U2136 ( .A1(n16958), .A2(vis_r8_o[25]), .B1(n2481), .B2(n16954), 
        .C1(n16981), .C2(vis_r9_o[25]), .ZN(n2479) );
  AOI222_X1 U2138 ( .A1(n16985), .A2(vis_r11_o[25]), .B1(n16972), .B2(n2484), 
        .C1(n16984), .C2(vis_r14_o[25]), .ZN(n2478) );
  AOI222_X1 U2141 ( .A1(n16967), .A2(vis_psp_o[23]), .B1(n16961), .B2(
        vis_r10_o[25]), .C1(n16975), .C2(vis_msp_o[23]), .ZN(n2477) );
  AOI22_X1 U2143 ( .A1(n16966), .A2(vis_r12_o[25]), .B1(n16976), .B2(n2460), 
        .ZN(n2476) );
  OAI22_X1 U2145 ( .A1(n16992), .A2(n4951), .B1(n2131), .B2(n2490), .ZN(n2475)
         );
  INV_X1 U2146 ( .A(n2490), .ZN(n4951) );
  OAI22_X1 U2147 ( .A1(n2491), .A2(n2492), .B1(n2248), .B2(n2493), .ZN(n2490)
         );
  INV_X1 U2148 ( .A(n2248), .ZN(n2491) );
  OAI22_X1 U2149 ( .A1(n5647), .A2(n17002), .B1(n2494), .B2(n17005), .ZN(
        U598_Z_0) );
  OAI22_X1 U2150 ( .A1(n5646), .A2(n16997), .B1(n2494), .B2(n17000), .ZN(
        U597_Z_0) );
  OAI22_X1 U2151 ( .A1(n5645), .A2(n17039), .B1(n2494), .B2(n17042), .ZN(
        U596_Z_0) );
  OAI22_X1 U2152 ( .A1(n5644), .A2(n17034), .B1(n2494), .B2(n17037), .ZN(
        U595_Z_0) );
  OAI22_X1 U2153 ( .A1(n4972), .A2(n17029), .B1(n2494), .B2(n17032), .ZN(
        U594_Z_0) );
  OAI22_X1 U2154 ( .A1(n5179), .A2(n17024), .B1(n2494), .B2(n17027), .ZN(
        U593_Z_0) );
  OAI22_X1 U2155 ( .A1(n4980), .A2(n17019), .B1(n2494), .B2(n17022), .ZN(
        U592_Z_0) );
  OAI22_X1 U2156 ( .A1(n5208), .A2(n17014), .B1(n2494), .B2(n17017), .ZN(
        U591_Z_0) );
  OAI22_X1 U2157 ( .A1(n5315), .A2(n17044), .B1(n2494), .B2(n17047), .ZN(
        U590_Z_0) );
  OAI22_X1 U2158 ( .A1(n5344), .A2(n17049), .B1(n2494), .B2(n17052), .ZN(
        U589_Z_0) );
  OAI22_X1 U2159 ( .A1(n5373), .A2(n17054), .B1(n2494), .B2(n17057), .ZN(
        U588_Z_0) );
  OAI22_X1 U2160 ( .A1(n5402), .A2(n17059), .B1(n2494), .B2(n17062), .ZN(
        U587_Z_0) );
  OAI22_X1 U2161 ( .A1(n5431), .A2(n17064), .B1(n2494), .B2(n17067), .ZN(
        U586_Z_0) );
  OAI22_X1 U2162 ( .A1(n5460), .A2(n17069), .B1(n2494), .B2(n17072), .ZN(
        U585_Z_0) );
  OAI22_X1 U2163 ( .A1(n4982), .A2(n17074), .B1(n2494), .B2(n17077), .ZN(
        U584_Z_0) );
  OAI22_X1 U2164 ( .A1(n5484), .A2(n17079), .B1(n2494), .B2(n17082), .ZN(
        U583_Z_0) );
  AOI221_X1 U2166 ( .B1(n2495), .B2(n16701), .C1(n2496), .C2(n17007), .A(n2497), .ZN(n2109) );
  INV_X1 U2167 ( .A(n2498), .ZN(n2497) );
  AOI211_X1 U2168 ( .C1(n2499), .C2(U163_Z_0), .A(n2055), .B(n2500), .ZN(n2498) );
  NOR3_X1 U2169 ( .A1(n1684), .A2(U163_Z_0), .A3(n16992), .ZN(n2500) );
  OAI22_X1 U2170 ( .A1(n2131), .A2(n1684), .B1(n2501), .B2(n1648), .ZN(n2499)
         );
  INV_X1 U2171 ( .A(n1648), .ZN(n1684) );
  NAND4_X1 U2172 ( .A1(n2502), .A2(n2503), .A3(n2504), .A4(n2505), .ZN(n1648)
         );
  AOI222_X1 U2173 ( .A1(n16973), .A2(vis_msp_o[22]), .B1(n16972), .B2(n2507), 
        .C1(n16967), .C2(vis_psp_o[22]), .ZN(n2505) );
  AOI222_X1 U2175 ( .A1(n16983), .A2(vis_r14_o[24]), .B1(n16964), .B2(
        vis_r12_o[24]), .C1(n16986), .C2(vis_r11_o[24]), .ZN(n2504) );
  AOI222_X1 U2178 ( .A1(n16979), .A2(vis_r9_o[24]), .B1(n16961), .B2(
        vis_r10_o[24]), .C1(n16958), .C2(vis_r8_o[24]), .ZN(n2503) );
  AOI22_X1 U2180 ( .A1(n16977), .A2(n2481), .B1(n16954), .B2(n2515), .ZN(n2502) );
  INV_X1 U2182 ( .A(n1337), .ZN(n109) );
  OAI221_X1 U2183 ( .B1(n2516), .B2(n2089), .C1(n2517), .C2(n2091), .A(n2518), 
        .ZN(n1337) );
  AOI221_X1 U2184 ( .B1(n2074), .B2(n2019), .C1(n2023), .C2(n2067), .A(n2076), 
        .ZN(n2518) );
  INV_X1 U2185 ( .A(n2069), .ZN(n2091) );
  INV_X1 U2186 ( .A(n2072), .ZN(n2089) );
  OAI22_X1 U2187 ( .A1(n5045), .A2(n17002), .B1(n16791), .B2(n17005), .ZN(
        U582_Z_0) );
  OAI22_X1 U2188 ( .A1(n5044), .A2(n16997), .B1(n16791), .B2(n17000), .ZN(
        U581_Z_0) );
  OAI22_X1 U2189 ( .A1(n5292), .A2(n17039), .B1(n16791), .B2(n17042), .ZN(
        U580_Z_0) );
  OAI22_X1 U2190 ( .A1(n5271), .A2(n17034), .B1(n16791), .B2(n17037), .ZN(
        U579_Z_0) );
  OAI22_X1 U2191 ( .A1(n5043), .A2(n17029), .B1(n16791), .B2(n17032), .ZN(
        U578_Z_0) );
  OAI22_X1 U2192 ( .A1(n5180), .A2(n17024), .B1(n16791), .B2(n17027), .ZN(
        U577_Z_0) );
  OAI22_X1 U2193 ( .A1(n5042), .A2(n17019), .B1(n16791), .B2(n17022), .ZN(
        U576_Z_0) );
  OAI22_X1 U2194 ( .A1(n5209), .A2(n17014), .B1(n16791), .B2(n17017), .ZN(
        U575_Z_0) );
  OAI22_X1 U2195 ( .A1(n5316), .A2(n17044), .B1(n16791), .B2(n17047), .ZN(
        U574_Z_0) );
  OAI22_X1 U2196 ( .A1(n5345), .A2(n17049), .B1(n16791), .B2(n17052), .ZN(
        U573_Z_0) );
  OAI22_X1 U2197 ( .A1(n5374), .A2(n17054), .B1(n16791), .B2(n17057), .ZN(
        U572_Z_0) );
  OAI22_X1 U2198 ( .A1(n5403), .A2(n17059), .B1(n16791), .B2(n17062), .ZN(
        U571_Z_0) );
  OAI22_X1 U2199 ( .A1(n5432), .A2(n17064), .B1(n16791), .B2(n17067), .ZN(
        U570_Z_0) );
  OAI22_X1 U2200 ( .A1(n5461), .A2(n17069), .B1(n16791), .B2(n17072), .ZN(
        U569_Z_0) );
  OAI22_X1 U2201 ( .A1(n5041), .A2(n17074), .B1(n16791), .B2(n17077), .ZN(
        U568_Z_0) );
  OAI22_X1 U2202 ( .A1(n5485), .A2(n17079), .B1(n16791), .B2(n17082), .ZN(
        U567_Z_0) );
  OR3_X1 U2204 ( .A1(n2522), .A2(n2523), .A3(n2524), .ZN(n2521) );
  NOR3_X1 U2205 ( .A1(n2161), .A2(n2501), .A3(n2525), .ZN(n2524) );
  INV_X1 U2206 ( .A(n2235), .ZN(n2523) );
  OAI221_X1 U2207 ( .B1(n2126), .B2(n2525), .C1(n5817), .C2(n2127), .A(n2161), 
        .ZN(n2235) );
  NAND4_X1 U2208 ( .A1(n2526), .A2(n2527), .A3(n2528), .A4(n2529), .ZN(n2161)
         );
  AOI222_X1 U2209 ( .A1(n16973), .A2(vis_msp_o[4]), .B1(n16972), .B2(n2531), 
        .C1(n16967), .C2(vis_psp_o[4]), .ZN(n2529) );
  AOI222_X1 U2210 ( .A1(n16982), .A2(vis_r14_o[6]), .B1(n16964), .B2(
        vis_r12_o[6]), .C1(n16985), .C2(vis_r11_o[6]), .ZN(n2528) );
  AOI222_X1 U2211 ( .A1(n16979), .A2(vis_r9_o[6]), .B1(n16961), .B2(
        vis_r10_o[6]), .C1(n16958), .C2(vis_r8_o[6]), .ZN(n2527) );
  AOI22_X1 U2212 ( .A1(n16977), .A2(n1152), .B1(n16954), .B2(n2539), .ZN(n2526) );
  INV_X1 U2213 ( .A(n5817), .ZN(n2525) );
  XOR2_X1 U2214 ( .A(n16990), .B(n2540), .Z(n5817) );
  AOI221_X1 U2215 ( .B1(n2541), .B2(n16671), .C1(n16988), .C2(n2250), .A(n2542), .ZN(n2540) );
  OAI22_X1 U2216 ( .A1(n5244), .A2(n2543), .B1(n5257), .B2(n2201), .ZN(n2542)
         );
  INV_X1 U2217 ( .A(n2200), .ZN(n2541) );
  AOI21_X1 U2218 ( .B1(n2124), .B2(n16782), .A(n2544), .ZN(n2522) );
  INV_X1 U2220 ( .A(n148), .ZN(n2520) );
  AOI221_X1 U2221 ( .B1(n2004), .B2(n2545), .C1(n2008), .C2(n2546), .A(n2547), 
        .ZN(n148) );
  INV_X1 U2222 ( .A(n2548), .ZN(n2547) );
  AOI221_X1 U2223 ( .B1(n2093), .B2(n2002), .C1(n2094), .C2(n2011), .A(n2012), 
        .ZN(n2548) );
  OAI22_X1 U2224 ( .A1(n5095), .A2(n17002), .B1(n2549), .B2(n17005), .ZN(
        U566_Z_0) );
  OAI22_X1 U2225 ( .A1(n5094), .A2(n16997), .B1(n2549), .B2(n17000), .ZN(
        U565_Z_0) );
  OAI22_X1 U2226 ( .A1(n5293), .A2(n17039), .B1(n2549), .B2(n17042), .ZN(
        U564_Z_0) );
  OAI22_X1 U2227 ( .A1(n5272), .A2(n17034), .B1(n2549), .B2(n17037), .ZN(
        U563_Z_0) );
  OAI22_X1 U2228 ( .A1(n5093), .A2(n17029), .B1(n2549), .B2(n17032), .ZN(
        U562_Z_0) );
  OAI22_X1 U2229 ( .A1(n5181), .A2(n17024), .B1(n2549), .B2(n17027), .ZN(
        U561_Z_0) );
  OAI22_X1 U2230 ( .A1(n5092), .A2(n17019), .B1(n2549), .B2(n17022), .ZN(
        U560_Z_0) );
  OAI22_X1 U2231 ( .A1(n5210), .A2(n17014), .B1(n2549), .B2(n17017), .ZN(
        U559_Z_0) );
  OAI22_X1 U2232 ( .A1(n5317), .A2(n17044), .B1(n2549), .B2(n17047), .ZN(
        U558_Z_0) );
  OAI22_X1 U2233 ( .A1(n5346), .A2(n17049), .B1(n2549), .B2(n17052), .ZN(
        U557_Z_0) );
  OAI22_X1 U2234 ( .A1(n5375), .A2(n17054), .B1(n2549), .B2(n17057), .ZN(
        U556_Z_0) );
  OAI22_X1 U2235 ( .A1(n5404), .A2(n17059), .B1(n2549), .B2(n17062), .ZN(
        U555_Z_0) );
  OAI22_X1 U2236 ( .A1(n5433), .A2(n17064), .B1(n2549), .B2(n17067), .ZN(
        U554_Z_0) );
  OAI22_X1 U2237 ( .A1(n5462), .A2(n17069), .B1(n2549), .B2(n17072), .ZN(
        U553_Z_0) );
  OAI22_X1 U2238 ( .A1(n5091), .A2(n17074), .B1(n2549), .B2(n17077), .ZN(
        U552_Z_0) );
  OAI22_X1 U2239 ( .A1(n5486), .A2(n17079), .B1(n2549), .B2(n17082), .ZN(
        U551_Z_0) );
  OAI221_X1 U2241 ( .B1(n2550), .B2(n5802), .C1(n16995), .C2(n1634), .A(n2551), 
        .ZN(n2281) );
  NAND3_X1 U2242 ( .A1(n2131), .A2(n1634), .A3(n5802), .ZN(n2551) );
  XOR2_X1 U2243 ( .A(n2552), .B(n16991), .Z(n5802) );
  OAI221_X1 U2244 ( .B1(n5256), .B2(n2201), .C1(n5100), .C2(n2554), .A(n2555), 
        .ZN(n2552) );
  AOI22_X1 U2245 ( .A1(n16988), .A2(n2556), .B1(n2198), .B2(n781), .ZN(n2555)
         );
  NOR2_X1 U2246 ( .A1(n1673), .A2(n16993), .ZN(n2550) );
  INV_X1 U2247 ( .A(n1634), .ZN(n1673) );
  NAND4_X1 U2248 ( .A1(n2557), .A2(n2558), .A3(n2559), .A4(n2560), .ZN(n1634)
         );
  AOI222_X1 U2249 ( .A1(n16973), .A2(vis_msp_o[3]), .B1(n16971), .B2(n2562), 
        .C1(n16967), .C2(vis_psp_o[3]), .ZN(n2560) );
  AOI222_X1 U2250 ( .A1(n16982), .A2(vis_r14_o[5]), .B1(n16964), .B2(
        vis_r12_o[5]), .C1(n16986), .C2(vis_r11_o[5]), .ZN(n2559) );
  AOI222_X1 U2251 ( .A1(n16979), .A2(vis_r9_o[5]), .B1(n16962), .B2(
        vis_r10_o[5]), .C1(n16958), .C2(vis_r8_o[5]), .ZN(n2558) );
  AOI22_X1 U2252 ( .A1(n16977), .A2(n2539), .B1(n16954), .B2(n2570), .ZN(n2557) );
  NAND2_X1 U2253 ( .A1(n16731), .A2(n17011), .ZN(n2263) );
  AOI221_X1 U2254 ( .B1(vis_ipsr_o[5]), .B2(n2227), .C1(n2556), .C2(n17007), 
        .A(n2055), .ZN(n2107) );
  AOI221_X1 U2255 ( .B1(n2410), .B2(n2011), .C1(n2415), .C2(n2004), .A(n2571), 
        .ZN(n152) );
  INV_X1 U2256 ( .A(n2572), .ZN(n2571) );
  AOI221_X1 U2257 ( .B1(n2008), .B2(n2414), .C1(n2411), .C2(n2002), .A(n2012), 
        .ZN(n2572) );
  OAI22_X1 U2258 ( .A1(n5125), .A2(n17002), .B1(n2573), .B2(n17005), .ZN(
        U550_Z_0) );
  OAI22_X1 U2259 ( .A1(n5124), .A2(n16997), .B1(n2573), .B2(n17000), .ZN(
        U549_Z_0) );
  OAI22_X1 U2260 ( .A1(n5294), .A2(n17039), .B1(n2573), .B2(n17042), .ZN(
        U548_Z_0) );
  OAI22_X1 U2261 ( .A1(n5273), .A2(n17034), .B1(n2573), .B2(n17037), .ZN(
        U547_Z_0) );
  OAI22_X1 U2262 ( .A1(n5123), .A2(n17029), .B1(n2573), .B2(n17032), .ZN(
        U546_Z_0) );
  OAI22_X1 U2263 ( .A1(n5182), .A2(n17024), .B1(n2573), .B2(n17027), .ZN(
        U545_Z_0) );
  OAI22_X1 U2264 ( .A1(n5122), .A2(n17019), .B1(n2573), .B2(n17022), .ZN(
        U544_Z_0) );
  OAI22_X1 U2265 ( .A1(n5211), .A2(n17014), .B1(n2573), .B2(n17017), .ZN(
        U543_Z_0) );
  OAI22_X1 U2266 ( .A1(n5318), .A2(n17044), .B1(n2573), .B2(n17047), .ZN(
        U542_Z_0) );
  OAI22_X1 U2267 ( .A1(n5347), .A2(n17049), .B1(n2573), .B2(n17052), .ZN(
        U541_Z_0) );
  OAI22_X1 U2268 ( .A1(n5376), .A2(n17054), .B1(n2573), .B2(n17057), .ZN(
        U540_Z_0) );
  OAI22_X1 U2269 ( .A1(n5405), .A2(n17059), .B1(n2573), .B2(n17062), .ZN(
        U539_Z_0) );
  OAI22_X1 U2270 ( .A1(n5434), .A2(n17064), .B1(n2573), .B2(n17067), .ZN(
        U538_Z_0) );
  OAI22_X1 U2271 ( .A1(n5463), .A2(n17069), .B1(n2573), .B2(n17072), .ZN(
        U537_Z_0) );
  OAI22_X1 U2272 ( .A1(n5121), .A2(n17074), .B1(n2573), .B2(n17077), .ZN(
        U536_Z_0) );
  OAI22_X1 U2273 ( .A1(n5487), .A2(n17079), .B1(n2573), .B2(n17082), .ZN(
        U535_Z_0) );
  OAI221_X1 U2275 ( .B1(n2574), .B2(n5801), .C1(n16995), .C2(n1636), .A(n2575), 
        .ZN(n2283) );
  NAND3_X1 U2276 ( .A1(n2131), .A2(n1636), .A3(n5801), .ZN(n2575) );
  XOR2_X1 U2277 ( .A(n16990), .B(n2576), .Z(n5801) );
  AOI221_X1 U2278 ( .B1(n16656), .B2(n2577), .C1(n16988), .C2(n2578), .A(n2579), .ZN(n2576) );
  OAI22_X1 U2279 ( .A1(n16794), .A2(n2543), .B1(n16810), .B2(n2201), .ZN(n2579) );
  NOR2_X1 U2280 ( .A1(n1674), .A2(n16993), .ZN(n2574) );
  INV_X1 U2281 ( .A(n1636), .ZN(n1674) );
  NAND4_X1 U2282 ( .A1(n2580), .A2(n2581), .A3(n2582), .A4(n2583), .ZN(n1636)
         );
  AOI222_X1 U2283 ( .A1(n16973), .A2(vis_msp_o[2]), .B1(n16971), .B2(n2585), 
        .C1(n16967), .C2(vis_psp_o[2]), .ZN(n2583) );
  AOI222_X1 U2284 ( .A1(n16982), .A2(vis_r14_o[4]), .B1(n16965), .B2(
        vis_r12_o[4]), .C1(n16986), .C2(vis_r11_o[4]), .ZN(n2582) );
  AOI222_X1 U2285 ( .A1(n16979), .A2(vis_r9_o[4]), .B1(n16962), .B2(
        vis_r10_o[4]), .C1(n16959), .C2(vis_r8_o[4]), .ZN(n2581) );
  AOI22_X1 U2286 ( .A1(n16977), .A2(n2570), .B1(n16954), .B2(n2593), .ZN(n2580) );
  NAND2_X1 U2287 ( .A1(n16730), .A2(n17011), .ZN(n2262) );
  AOI221_X1 U2288 ( .B1(vis_ipsr_o[4]), .B2(n2227), .C1(n2578), .C2(n17007), 
        .A(n2055), .ZN(n2112) );
  AOI221_X1 U2289 ( .B1(n2066), .B2(n2011), .C1(n2068), .C2(n2004), .A(n2594), 
        .ZN(n160) );
  INV_X1 U2290 ( .A(n2595), .ZN(n2594) );
  AOI221_X1 U2291 ( .B1(n2008), .B2(n2073), .C1(n2002), .C2(n2075), .A(n2012), 
        .ZN(n2595) );
  INV_X1 U2292 ( .A(n2596), .ZN(n2073) );
  OAI22_X1 U2293 ( .A1(n5032), .A2(n17002), .B1(n2597), .B2(n17005), .ZN(
        U534_Z_0) );
  OAI22_X1 U2294 ( .A1(n5031), .A2(n16997), .B1(n2597), .B2(n17000), .ZN(
        U533_Z_0) );
  OAI22_X1 U2295 ( .A1(n5295), .A2(n17039), .B1(n2597), .B2(n17042), .ZN(
        U532_Z_0) );
  OAI22_X1 U2296 ( .A1(n5274), .A2(n17034), .B1(n2597), .B2(n17037), .ZN(
        U531_Z_0) );
  OAI22_X1 U2297 ( .A1(n5030), .A2(n17029), .B1(n2597), .B2(n17032), .ZN(
        U530_Z_0) );
  OAI22_X1 U2298 ( .A1(n5183), .A2(n17024), .B1(n2597), .B2(n17027), .ZN(
        U529_Z_0) );
  OAI22_X1 U2299 ( .A1(n5029), .A2(n17019), .B1(n2597), .B2(n17022), .ZN(
        U528_Z_0) );
  OAI22_X1 U2300 ( .A1(n5212), .A2(n17014), .B1(n2597), .B2(n17017), .ZN(
        U527_Z_0) );
  OAI22_X1 U2301 ( .A1(n5319), .A2(n17044), .B1(n2597), .B2(n17047), .ZN(
        U526_Z_0) );
  OAI22_X1 U2302 ( .A1(n5348), .A2(n17049), .B1(n2597), .B2(n17052), .ZN(
        U525_Z_0) );
  OAI22_X1 U2303 ( .A1(n5377), .A2(n17054), .B1(n2597), .B2(n17057), .ZN(
        U524_Z_0) );
  OAI22_X1 U2304 ( .A1(n5406), .A2(n17059), .B1(n2597), .B2(n17062), .ZN(
        U523_Z_0) );
  OAI22_X1 U2305 ( .A1(n5435), .A2(n17064), .B1(n2597), .B2(n17067), .ZN(
        U522_Z_0) );
  OAI22_X1 U2306 ( .A1(n5464), .A2(n17069), .B1(n2597), .B2(n17072), .ZN(
        U521_Z_0) );
  OAI22_X1 U2307 ( .A1(n5028), .A2(n17074), .B1(n2597), .B2(n17077), .ZN(
        U520_Z_0) );
  OAI22_X1 U2308 ( .A1(n5488), .A2(n17079), .B1(n2597), .B2(n17082), .ZN(
        U519_Z_0) );
  AOI222_X1 U2310 ( .A1(n17006), .A2(n2257), .B1(n16682), .B2(n17010), .C1(
        n2032), .C2(n2055), .ZN(n2598) );
  INV_X1 U2311 ( .A(n2599), .ZN(n2032) );
  INV_X1 U2312 ( .A(n2600), .ZN(n2111) );
  OAI221_X1 U2313 ( .B1(n2601), .B2(n2602), .C1(n170), .C2(n2164), .A(n2603), 
        .ZN(n2600) );
  NAND3_X1 U2314 ( .A1(n2604), .A2(n2127), .A3(n2602), .ZN(n2603) );
  INV_X1 U2315 ( .A(n2227), .ZN(n2164) );
  INV_X1 U2316 ( .A(add_2082_B_4_), .ZN(n2602) );
  XOR2_X1 U2317 ( .A(n2605), .B(n16991), .Z(add_2082_B_4_) );
  OAI221_X1 U2318 ( .B1(n5100), .B2(n2201), .C1(n5027), .C2(n2554), .A(n2606), 
        .ZN(n2605) );
  AOI22_X1 U2319 ( .A1(n16989), .A2(n2257), .B1(n2198), .B2(n454), .ZN(n2606)
         );
  AOI22_X1 U2320 ( .A1(n1638), .A2(n16994), .B1(n2604), .B2(n2126), .ZN(n2601)
         );
  INV_X1 U2321 ( .A(n2604), .ZN(n1638) );
  NAND4_X1 U2322 ( .A1(n2607), .A2(n2608), .A3(n2609), .A4(n2610), .ZN(n2604)
         );
  AOI222_X1 U2323 ( .A1(n16973), .A2(vis_msp_o[1]), .B1(n16971), .B2(n2612), 
        .C1(n16968), .C2(vis_psp_o[1]), .ZN(n2610) );
  AOI222_X1 U2324 ( .A1(n16982), .A2(vis_r14_o[3]), .B1(n16965), .B2(
        vis_r12_o[3]), .C1(n16986), .C2(vis_r11_o[3]), .ZN(n2609) );
  AOI222_X1 U2325 ( .A1(n16979), .A2(vis_r9_o[3]), .B1(n16962), .B2(
        vis_r10_o[3]), .C1(n16959), .C2(vis_r8_o[3]), .ZN(n2608) );
  AOI22_X1 U2326 ( .A1(n16977), .A2(n2593), .B1(n16955), .B2(n2620), .ZN(n2607) );
  AOI221_X1 U2327 ( .B1(n2421), .B2(n2002), .C1(n2422), .C2(n2004), .A(n2621), 
        .ZN(n166) );
  INV_X1 U2328 ( .A(n2622), .ZN(n2621) );
  AOI221_X1 U2329 ( .B1(n2623), .B2(n2008), .C1(n2624), .C2(n2011), .A(n2012), 
        .ZN(n2622) );
  OAI22_X1 U2330 ( .A1(n5102), .A2(n980), .B1(n683), .B2(n1811), .ZN(U518_Z_0)
         );
  OAI222_X1 U2334 ( .A1(n16957), .A2(n2628), .B1(n16837), .B2(n1027), .C1(
        n16856), .C2(n782), .ZN(n2627) );
  OAI221_X1 U2335 ( .B1(n2629), .B2(n16829), .C1(n16826), .C2(n1857), .A(n2630), .ZN(n2626) );
  NAND3_X1 U2336 ( .A1(n16806), .A2(n16851), .A3(n2631), .ZN(n2630) );
  AOI21_X1 U2337 ( .B1(n1564), .B2(n565), .A(n1606), .ZN(n2629) );
  NAND3_X1 U2338 ( .A1(n2632), .A2(n2633), .A3(n2634), .ZN(n2232) );
  AOI221_X1 U2339 ( .B1(n16976), .B2(n2635), .C1(n16956), .C2(n2188), .A(n2636), .ZN(n2634) );
  OAI22_X1 U2340 ( .A1(n5366), .A2(n2637), .B1(n5395), .B2(n2190), .ZN(n2636)
         );
  AOI222_X1 U2342 ( .A1(n16985), .A2(vis_r11_o[1]), .B1(n16971), .B2(n2639), 
        .C1(n16964), .C2(vis_r12_o[1]), .ZN(n2633) );
  AOI22_X1 U2343 ( .A1(n16984), .A2(vis_r14_o[1]), .B1(n16963), .B2(
        vis_r10_o[1]), .ZN(n2632) );
  AOI222_X1 U2348 ( .A1(n1806), .A2(n16836), .B1(n2628), .B2(n16954), .C1(
        n2646), .C2(n16828), .ZN(n2645) );
  INV_X1 U2349 ( .A(n919), .ZN(n1806) );
  NAND4_X1 U2350 ( .A1(n1103), .A2(n16867), .A3(n673), .A4(n2647), .ZN(n2643)
         );
  AOI21_X1 U2351 ( .B1(n1561), .B2(n502), .A(n611), .ZN(n2647) );
  INV_X1 U2352 ( .A(n1218), .ZN(n502) );
  XOR2_X1 U2353 ( .A(n4973), .B(n1106), .Z(n2625) );
  OAI21_X1 U2354 ( .B1(n1007), .B2(n187), .A(n1008), .ZN(n1106) );
  AOI21_X1 U2356 ( .B1(n16845), .B2(n1563), .A(n943), .ZN(n187) );
  INV_X1 U2357 ( .A(n1217), .ZN(n943) );
  NAND2_X1 U2358 ( .A1(n483), .A2(n16728), .ZN(n1217) );
  INV_X1 U2359 ( .A(n846), .ZN(n1563) );
  NAND2_X1 U2360 ( .A1(n16869), .A2(n16839), .ZN(n846) );
  AND3_X1 U2361 ( .A1(n2648), .A2(n2649), .A3(n2650), .ZN(n1007) );
  NOR4_X1 U2362 ( .A1(n2651), .A2(n2652), .A3(n2653), .A4(n2654), .ZN(n2650)
         );
  NOR4_X1 U2363 ( .A1(n16836), .A2(n16819), .A3(n1519), .A4(n604), .ZN(n2654)
         );
  NOR4_X1 U2364 ( .A1(n1086), .A2(n16858), .A3(n1104), .A4(n498), .ZN(n2653)
         );
  NAND2_X1 U2365 ( .A1(n16834), .A2(n16821), .ZN(n498) );
  INV_X1 U2366 ( .A(n2655), .ZN(n2652) );
  OAI211_X1 U2367 ( .C1(n998), .C2(n542), .A(n566), .B(n715), .ZN(n2655) );
  OAI33_X1 U2368 ( .A1(n532), .A2(n1218), .A3(n917), .B1(n648), .B2(n16833), 
        .B3(n16805), .ZN(n2651) );
  AOI22_X1 U2369 ( .A1(n2656), .A2(n596), .B1(n757), .B2(n2657), .ZN(n2649) );
  NAND4_X1 U2370 ( .A1(n16866), .A2(n918), .A3(n1856), .A4(n1579), .ZN(n2657)
         );
  NAND2_X1 U2371 ( .A1(n2658), .A2(n2659), .ZN(n2656) );
  NAND3_X1 U2372 ( .A1(n991), .A2(n1574), .A3(n1095), .ZN(n2659) );
  AOI22_X1 U2373 ( .A1(n2660), .A2(n16826), .B1(n2661), .B2(n2662), .ZN(n2648)
         );
  NAND4_X1 U2374 ( .A1(n1857), .A2(n694), .A3(n2663), .A4(n2664), .ZN(n2660)
         );
  AOI221_X1 U2375 ( .B1(n897), .B2(n16728), .C1(n527), .C2(n16808), .A(n2665), 
        .ZN(n2664) );
  OAI22_X1 U2376 ( .A1(n605), .A2(n745), .B1(n556), .B2(n616), .ZN(n2665) );
  AOI21_X1 U2377 ( .B1(n2666), .B2(n596), .A(n2667), .ZN(n2663) );
  NOR3_X1 U2378 ( .A1(n16808), .A2(n16845), .A3(n585), .ZN(n2667) );
  OAI21_X1 U2380 ( .B1(n2668), .B2(n16830), .A(n2669), .ZN(n2666) );
  NAND3_X1 U2381 ( .A1(n592), .A2(n1574), .A3(n16804), .ZN(n2669) );
  AOI222_X1 U2382 ( .A1(n592), .A2(n2670), .B1(n2671), .B2(n466), .C1(n2672), 
        .C2(n1468), .ZN(n2668) );
  NOR2_X1 U2383 ( .A1(n16851), .A2(n1469), .ZN(n2671) );
  INV_X1 U2384 ( .A(n2673), .ZN(n2670) );
  NOR4_X1 U2387 ( .A1(n2678), .A2(n2679), .A3(n2680), .A4(n2681), .ZN(n2677)
         );
  NOR4_X1 U2388 ( .A1(n16694), .A2(n1086), .A3(n917), .A4(n762), .ZN(n2681) );
  INV_X1 U2389 ( .A(n1177), .ZN(n2680) );
  AND3_X1 U2390 ( .A1(n1561), .A2(n1094), .A3(n809), .ZN(n2679) );
  NOR2_X1 U2391 ( .A1(n16826), .A2(n16851), .ZN(n1561) );
  OAI33_X1 U2392 ( .A1(n713), .A2(n16836), .A3(n616), .B1(n524), .B2(n16858), 
        .B3(n16808), .ZN(n2678) );
  AOI21_X1 U2393 ( .B1(n2682), .B2(n16864), .A(n2683), .ZN(n2676) );
  OAI33_X1 U2394 ( .A1(n696), .A2(n16821), .A3(n715), .B1(n945), .B2(n16845), 
        .B3(n16828), .ZN(n2683) );
  OAI211_X1 U2395 ( .C1(n16824), .C2(n1857), .A(n2684), .B(n1279), .ZN(n2682)
         );
  NAND3_X1 U2396 ( .A1(n809), .A2(n16824), .A3(n5165), .ZN(n1279) );
  INV_X1 U2397 ( .A(n609), .ZN(n2684) );
  NAND2_X1 U2398 ( .A1(n563), .A2(n1574), .ZN(n1857) );
  NAND2_X1 U2399 ( .A1(n660), .A2(n1034), .ZN(n2675) );
  INV_X1 U2400 ( .A(n1811), .ZN(n980) );
  NAND2_X1 U2401 ( .A1(n17124), .A2(hprot_o[0]), .ZN(n1811) );
  NOR4_X1 U2403 ( .A1(n2687), .A2(n1272), .A3(n615), .A4(n2688), .ZN(n2686) );
  INV_X1 U2404 ( .A(n1025), .ZN(n2688) );
  NAND3_X1 U2405 ( .A1(n827), .A2(n16824), .A3(n660), .ZN(n1025) );
  NOR2_X1 U2406 ( .A1(n558), .A2(n16871), .ZN(n660) );
  INV_X1 U2407 ( .A(n646), .ZN(n615) );
  NAND2_X1 U2408 ( .A1(n798), .A2(n590), .ZN(n646) );
  NOR3_X1 U2409 ( .A1(n641), .A2(n745), .A3(n808), .ZN(n1272) );
  OAI33_X1 U2410 ( .A1(n650), .A2(n16833), .A3(n16826), .B1(n2689), .B2(n16858), .B3(n640), .ZN(n2687) );
  AOI222_X1 U2411 ( .A1(n1037), .A2(n16856), .B1(n2690), .B2(n506), .C1(n609), 
        .C2(n991), .ZN(n2685) );
  NOR2_X1 U2412 ( .A1(n1307), .A2(n558), .ZN(n609) );
  NOR2_X1 U2413 ( .A1(n16848), .A2(n808), .ZN(n2690) );
  NOR3_X1 U2415 ( .A1(n16821), .A2(n1467), .A3(n699), .ZN(n1037) );
  INV_X1 U2416 ( .A(n2691), .ZN(n2674) );
  OAI211_X1 U2417 ( .C1(n16833), .C2(n499), .A(n1024), .B(n1476), .ZN(n2691)
         );
  AND2_X1 U2418 ( .A1(n2692), .A2(n1957), .ZN(n1476) );
  OAI21_X1 U2419 ( .B1(n506), .B2(n1306), .A(n526), .ZN(n2692) );
  NOR2_X1 U2420 ( .A1(n610), .A2(n696), .ZN(n1306) );
  NAND2_X1 U2421 ( .A1(n695), .A2(n590), .ZN(n1024) );
  INV_X1 U2422 ( .A(n650), .ZN(n590) );
  NOR2_X1 U2423 ( .A1(n16859), .A2(n16856), .ZN(n695) );
  INV_X1 U2424 ( .A(n2693), .ZN(n1876) );
  OAI33_X1 U2425 ( .A1(n1517), .A2(n16826), .A3(n1882), .B1(n558), .B2(n16833), 
        .B3(n715), .ZN(n2693) );
  NAND2_X1 U2426 ( .A1(n16680), .A2(n592), .ZN(n558) );
  OAI22_X1 U2427 ( .A1(n5052), .A2(n17002), .B1(n2694), .B2(n17005), .ZN(
        U517_Z_0) );
  OAI22_X1 U2428 ( .A1(n5051), .A2(n16997), .B1(n2694), .B2(n17000), .ZN(
        U516_Z_0) );
  OAI22_X1 U2429 ( .A1(n5296), .A2(n17039), .B1(n2694), .B2(n17042), .ZN(
        U515_Z_0) );
  OAI22_X1 U2430 ( .A1(n5275), .A2(n17034), .B1(n2694), .B2(n17037), .ZN(
        U514_Z_0) );
  OAI22_X1 U2431 ( .A1(n5050), .A2(n17029), .B1(n2694), .B2(n17032), .ZN(
        U513_Z_0) );
  OAI22_X1 U2432 ( .A1(n5184), .A2(n17024), .B1(n2694), .B2(n17027), .ZN(
        U512_Z_0) );
  OAI22_X1 U2433 ( .A1(n5049), .A2(n17019), .B1(n2694), .B2(n17022), .ZN(
        U511_Z_0) );
  OAI22_X1 U2434 ( .A1(n5213), .A2(n17014), .B1(n2694), .B2(n17017), .ZN(
        U510_Z_0) );
  OAI22_X1 U2435 ( .A1(n5320), .A2(n17044), .B1(n2694), .B2(n17047), .ZN(
        U509_Z_0) );
  OAI22_X1 U2436 ( .A1(n5349), .A2(n17049), .B1(n2694), .B2(n17052), .ZN(
        U508_Z_0) );
  OAI22_X1 U2437 ( .A1(n5378), .A2(n17054), .B1(n2694), .B2(n17057), .ZN(
        U507_Z_0) );
  OAI22_X1 U2438 ( .A1(n5407), .A2(n17059), .B1(n2694), .B2(n17062), .ZN(
        U506_Z_0) );
  OAI22_X1 U2439 ( .A1(n5436), .A2(n17064), .B1(n2694), .B2(n17067), .ZN(
        U505_Z_0) );
  OAI22_X1 U2440 ( .A1(n5465), .A2(n17069), .B1(n2694), .B2(n17072), .ZN(
        U504_Z_0) );
  OAI22_X1 U2441 ( .A1(n5048), .A2(n17074), .B1(n2694), .B2(n17077), .ZN(
        U503_Z_0) );
  OAI22_X1 U2442 ( .A1(n5489), .A2(n17079), .B1(n2694), .B2(n17082), .ZN(
        U502_Z_0) );
  AOI221_X1 U2444 ( .B1(n17006), .B2(n2251), .C1(n16702), .C2(n17010), .A(
        n2698), .ZN(n2697) );
  INV_X1 U2445 ( .A(n2282), .ZN(n2698) );
  OAI221_X1 U2446 ( .B1(n2126), .B2(n2699), .C1(n5816), .C2(n2127), .A(n1650), 
        .ZN(n2282) );
  INV_X1 U2447 ( .A(n5816), .ZN(n2699) );
  NAND3_X1 U2448 ( .A1(n5816), .A2(n16994), .A3(n1686), .ZN(n2695) );
  INV_X1 U2449 ( .A(n1650), .ZN(n1686) );
  NAND4_X1 U2450 ( .A1(n2700), .A2(n2701), .A3(n2702), .A4(n2703), .ZN(n1650)
         );
  AOI222_X1 U2451 ( .A1(n16973), .A2(vis_msp_o[20]), .B1(n16971), .B2(n2705), 
        .C1(n16968), .C2(vis_psp_o[20]), .ZN(n2703) );
  AOI222_X1 U2453 ( .A1(n16982), .A2(vis_r14_o[22]), .B1(n16965), .B2(
        vis_r12_o[22]), .C1(n16986), .C2(vis_r11_o[22]), .ZN(n2702) );
  AOI222_X1 U2456 ( .A1(n16980), .A2(vis_r9_o[22]), .B1(n16962), .B2(
        vis_r10_o[22]), .C1(n16959), .C2(vis_r8_o[22]), .ZN(n2701) );
  AOI22_X1 U2458 ( .A1(n16977), .A2(n2713), .B1(n16955), .B2(n2714), .ZN(n2700) );
  XOR2_X1 U2459 ( .A(n16990), .B(n2715), .Z(n5816) );
  AOI221_X1 U2460 ( .B1(n2716), .B2(n16813), .C1(n16988), .C2(n2251), .A(n2717), .ZN(n2715) );
  NAND2_X1 U2461 ( .A1(n2718), .A2(n2719), .ZN(n2717) );
  NAND3_X1 U2462 ( .A1(n5254), .A2(n2198), .A3(n16812), .ZN(n2718) );
  AOI221_X1 U2463 ( .B1(n2720), .B2(n2094), .C1(n2721), .C2(n2093), .A(n2722), 
        .ZN(n61) );
  OAI22_X1 U2464 ( .A1(n2723), .A2(n2090), .B1(n2088), .B2(n2724), .ZN(n2722)
         );
  OAI22_X1 U2465 ( .A1(n5624), .A2(n17002), .B1(n2725), .B2(n17005), .ZN(
        U501_Z_0) );
  OAI22_X1 U2466 ( .A1(n5623), .A2(n16997), .B1(n2725), .B2(n17000), .ZN(
        U500_Z_0) );
  OAI22_X1 U2467 ( .A1(n5622), .A2(n17039), .B1(n2725), .B2(n17042), .ZN(
        U499_Z_0) );
  OAI22_X1 U2468 ( .A1(n5621), .A2(n17034), .B1(n2725), .B2(n17037), .ZN(
        U498_Z_0) );
  OAI22_X1 U2469 ( .A1(n5117), .A2(n17029), .B1(n2725), .B2(n17032), .ZN(
        U497_Z_0) );
  OAI22_X1 U2470 ( .A1(n5185), .A2(n17024), .B1(n2725), .B2(n17027), .ZN(
        U496_Z_0) );
  OAI22_X1 U2471 ( .A1(n5116), .A2(n17019), .B1(n2725), .B2(n17022), .ZN(
        U495_Z_0) );
  OAI22_X1 U2472 ( .A1(n5214), .A2(n17014), .B1(n2725), .B2(n17017), .ZN(
        U494_Z_0) );
  OAI22_X1 U2473 ( .A1(n5321), .A2(n17044), .B1(n2725), .B2(n17047), .ZN(
        U493_Z_0) );
  OAI22_X1 U2474 ( .A1(n5350), .A2(n17049), .B1(n2725), .B2(n17052), .ZN(
        U492_Z_0) );
  OAI22_X1 U2475 ( .A1(n5379), .A2(n17054), .B1(n2725), .B2(n17057), .ZN(
        U491_Z_0) );
  OAI22_X1 U2476 ( .A1(n5408), .A2(n17059), .B1(n2725), .B2(n17062), .ZN(
        U490_Z_0) );
  OAI22_X1 U2477 ( .A1(n5437), .A2(n17064), .B1(n2725), .B2(n17067), .ZN(
        U489_Z_0) );
  OAI22_X1 U2478 ( .A1(n5466), .A2(n17069), .B1(n2725), .B2(n17072), .ZN(
        U488_Z_0) );
  OAI22_X1 U2479 ( .A1(n5115), .A2(n17074), .B1(n2725), .B2(n17077), .ZN(
        U487_Z_0) );
  OAI22_X1 U2480 ( .A1(n5490), .A2(n17079), .B1(n2725), .B2(n17082), .ZN(
        U486_Z_0) );
  AOI222_X1 U2482 ( .A1(n17007), .A2(n21), .B1(n2727), .B2(n2728), .C1(n16668), 
        .C2(n17009), .ZN(n2726) );
  NAND3_X1 U2483 ( .A1(n2131), .A2(n1651), .A3(n5815), .ZN(n2728) );
  OAI21_X1 U2484 ( .B1(n16993), .B2(n1687), .A(n2729), .ZN(n2727) );
  OAI21_X1 U2485 ( .B1(n16994), .B2(n1651), .A(n5815), .ZN(n2729) );
  AOI221_X1 U2487 ( .B1(n16989), .B2(n21), .C1(n2198), .C2(n2731), .A(n2732), 
        .ZN(n2730) );
  INV_X1 U2488 ( .A(n1651), .ZN(n1687) );
  NAND4_X1 U2489 ( .A1(n2733), .A2(n2734), .A3(n2735), .A4(n2736), .ZN(n1651)
         );
  AOI222_X1 U2490 ( .A1(n16974), .A2(vis_msp_o[19]), .B1(n16971), .B2(n2738), 
        .C1(n16968), .C2(vis_psp_o[19]), .ZN(n2736) );
  AOI222_X1 U2492 ( .A1(n16983), .A2(vis_r14_o[21]), .B1(n16965), .B2(
        vis_r12_o[21]), .C1(n16986), .C2(vis_r11_o[21]), .ZN(n2735) );
  AOI222_X1 U2495 ( .A1(n16980), .A2(vis_r9_o[21]), .B1(n16962), .B2(
        vis_r10_o[21]), .C1(n16959), .C2(vis_r8_o[21]), .ZN(n2734) );
  AOI22_X1 U2497 ( .A1(n16977), .A2(n2714), .B1(n16955), .B2(n2746), .ZN(n2733) );
  AOI221_X1 U2499 ( .B1(n2720), .B2(n2410), .C1(n2721), .C2(n2411), .A(n2747), 
        .ZN(n58) );
  INV_X1 U2500 ( .A(n2748), .ZN(n2747) );
  AOI22_X1 U2501 ( .A1(n2074), .A2(n2415), .B1(n2414), .B2(n2749), .ZN(n2748)
         );
  OAI22_X1 U2502 ( .A1(n5617), .A2(n17002), .B1(n2750), .B2(n17005), .ZN(
        U483_Z_0) );
  OAI22_X1 U2503 ( .A1(n5616), .A2(n16997), .B1(n2750), .B2(n17000), .ZN(
        U482_Z_0) );
  OAI22_X1 U2504 ( .A1(n5615), .A2(n17039), .B1(n2750), .B2(n17042), .ZN(
        U481_Z_0) );
  OAI22_X1 U2505 ( .A1(n5614), .A2(n17034), .B1(n2750), .B2(n17037), .ZN(
        U480_Z_0) );
  OAI22_X1 U2506 ( .A1(n5613), .A2(n17029), .B1(n2750), .B2(n17032), .ZN(
        U479_Z_0) );
  OAI22_X1 U2507 ( .A1(n5612), .A2(n17024), .B1(n2750), .B2(n17027), .ZN(
        U478_Z_0) );
  OAI22_X1 U2508 ( .A1(n5611), .A2(n17019), .B1(n2750), .B2(n17022), .ZN(
        U477_Z_0) );
  OAI22_X1 U2509 ( .A1(n5610), .A2(n17014), .B1(n2750), .B2(n17017), .ZN(
        U476_Z_0) );
  OAI22_X1 U2510 ( .A1(n5609), .A2(n17044), .B1(n2750), .B2(n17047), .ZN(
        U475_Z_0) );
  OAI22_X1 U2511 ( .A1(n5608), .A2(n17049), .B1(n2750), .B2(n17052), .ZN(
        U474_Z_0) );
  OAI22_X1 U2512 ( .A1(n5607), .A2(n17054), .B1(n2750), .B2(n17057), .ZN(
        U473_Z_0) );
  OAI22_X1 U2513 ( .A1(n5606), .A2(n17059), .B1(n2750), .B2(n17062), .ZN(
        U472_Z_0) );
  OAI22_X1 U2514 ( .A1(n5605), .A2(n17064), .B1(n2750), .B2(n17067), .ZN(
        U471_Z_0) );
  OAI22_X1 U2515 ( .A1(n5604), .A2(n17069), .B1(n2750), .B2(n17072), .ZN(
        U470_Z_0) );
  OAI22_X1 U2516 ( .A1(n5603), .A2(n17074), .B1(n2750), .B2(n17077), .ZN(
        U469_Z_0) );
  OAI22_X1 U2517 ( .A1(n5602), .A2(n17079), .B1(n2750), .B2(n17082), .ZN(
        U468_Z_0) );
  AOI221_X1 U2519 ( .B1(n17006), .B2(n20), .C1(n16706), .C2(n17010), .A(n2754), 
        .ZN(n2753) );
  INV_X1 U2520 ( .A(n2284), .ZN(n2754) );
  OAI221_X1 U2521 ( .B1(n2126), .B2(n2755), .C1(n5814), .C2(n2127), .A(n1653), 
        .ZN(n2284) );
  INV_X1 U2522 ( .A(n5814), .ZN(n2755) );
  INV_X1 U2523 ( .A(n55), .ZN(n2752) );
  OAI221_X1 U2524 ( .B1(n2756), .B2(n2757), .C1(n2724), .C2(n2596), .A(n2758), 
        .ZN(n55) );
  AOI22_X1 U2525 ( .A1(n2074), .A2(n2068), .B1(n2075), .B2(n2721), .ZN(n2758)
         );
  NAND3_X1 U2526 ( .A1(n5814), .A2(n16994), .A3(n1688), .ZN(n2751) );
  INV_X1 U2527 ( .A(n1653), .ZN(n1688) );
  NAND4_X1 U2528 ( .A1(n2759), .A2(n2760), .A3(n2761), .A4(n2762), .ZN(n1653)
         );
  AOI222_X1 U2529 ( .A1(n16974), .A2(vis_msp_o[18]), .B1(n16971), .B2(n2764), 
        .C1(n16968), .C2(vis_psp_o[18]), .ZN(n2762) );
  AOI222_X1 U2531 ( .A1(n16983), .A2(vis_r14_o[20]), .B1(n16965), .B2(
        vis_r12_o[20]), .C1(n16986), .C2(vis_r11_o[20]), .ZN(n2761) );
  AOI222_X1 U2534 ( .A1(n16980), .A2(vis_r9_o[20]), .B1(n16962), .B2(
        vis_r10_o[20]), .C1(n16959), .C2(vis_r8_o[20]), .ZN(n2760) );
  AOI22_X1 U2536 ( .A1(n16977), .A2(n2746), .B1(n16955), .B2(n2772), .ZN(n2759) );
  XOR2_X1 U2538 ( .A(n16990), .B(n2773), .Z(n5814) );
  AOI221_X1 U2539 ( .B1(n16989), .B2(n20), .C1(n2198), .C2(n2774), .A(n2732), 
        .ZN(n2773) );
  OAI22_X1 U2540 ( .A1(n5638), .A2(n17002), .B1(n2775), .B2(n17005), .ZN(
        U467_Z_0) );
  OAI22_X1 U2541 ( .A1(n5637), .A2(n16997), .B1(n2775), .B2(n17000), .ZN(
        U466_Z_0) );
  OAI22_X1 U2542 ( .A1(n5636), .A2(n17039), .B1(n2775), .B2(n17042), .ZN(
        U465_Z_0) );
  OAI22_X1 U2543 ( .A1(n5635), .A2(n17034), .B1(n2775), .B2(n17037), .ZN(
        U464_Z_0) );
  OAI22_X1 U2544 ( .A1(n5090), .A2(n17029), .B1(n2775), .B2(n17032), .ZN(
        U463_Z_0) );
  OAI22_X1 U2545 ( .A1(n5186), .A2(n17024), .B1(n2775), .B2(n17027), .ZN(
        U462_Z_0) );
  OAI22_X1 U2546 ( .A1(n5089), .A2(n17019), .B1(n2775), .B2(n17022), .ZN(
        U461_Z_0) );
  OAI22_X1 U2547 ( .A1(n5215), .A2(n17014), .B1(n2775), .B2(n17017), .ZN(
        U460_Z_0) );
  OAI22_X1 U2548 ( .A1(n5322), .A2(n17044), .B1(n2775), .B2(n17047), .ZN(
        U459_Z_0) );
  OAI22_X1 U2549 ( .A1(n5351), .A2(n17049), .B1(n2775), .B2(n17052), .ZN(
        U458_Z_0) );
  OAI22_X1 U2550 ( .A1(n5380), .A2(n17054), .B1(n2775), .B2(n17057), .ZN(
        U457_Z_0) );
  OAI22_X1 U2551 ( .A1(n5409), .A2(n17059), .B1(n2775), .B2(n17062), .ZN(
        U456_Z_0) );
  OAI22_X1 U2552 ( .A1(n5438), .A2(n17064), .B1(n2775), .B2(n17067), .ZN(
        U455_Z_0) );
  OAI22_X1 U2553 ( .A1(n5467), .A2(n17069), .B1(n2775), .B2(n17072), .ZN(
        U454_Z_0) );
  OAI22_X1 U2554 ( .A1(n5088), .A2(n17074), .B1(n2775), .B2(n17077), .ZN(
        U453_Z_0) );
  OAI22_X1 U2555 ( .A1(n5491), .A2(n17079), .B1(n2775), .B2(n17082), .ZN(
        U452_Z_0) );
  AOI222_X1 U2557 ( .A1(n17007), .A2(n22), .B1(n2778), .B2(n2779), .C1(n16709), 
        .C2(n17009), .ZN(n2777) );
  NAND3_X1 U2558 ( .A1(n2131), .A2(n2156), .A3(n5813), .ZN(n2779) );
  OAI21_X1 U2559 ( .B1(n16993), .B2(n1654), .A(n2780), .ZN(n2778) );
  OAI21_X1 U2560 ( .B1(n16994), .B2(n2156), .A(n5813), .ZN(n2780) );
  XOR2_X1 U2561 ( .A(n16990), .B(n2781), .Z(n5813) );
  AOI221_X1 U2562 ( .B1(n16989), .B2(n22), .C1(n2198), .C2(n486), .A(n2732), 
        .ZN(n2781) );
  INV_X1 U2563 ( .A(n2156), .ZN(n1654) );
  NAND4_X1 U2564 ( .A1(n2782), .A2(n2783), .A3(n2784), .A4(n2785), .ZN(n2156)
         );
  AOI222_X1 U2565 ( .A1(n16974), .A2(vis_msp_o[17]), .B1(n16971), .B2(n2787), 
        .C1(n16968), .C2(vis_psp_o[17]), .ZN(n2785) );
  AOI222_X1 U2567 ( .A1(n16983), .A2(vis_r14_o[19]), .B1(n16965), .B2(
        vis_r12_o[19]), .C1(n16986), .C2(vis_r11_o[19]), .ZN(n2784) );
  AOI222_X1 U2570 ( .A1(n16980), .A2(vis_r9_o[19]), .B1(n16962), .B2(
        vis_r10_o[19]), .C1(n16959), .C2(vis_r8_o[19]), .ZN(n2783) );
  AOI22_X1 U2572 ( .A1(n16977), .A2(n2772), .B1(n16955), .B2(n2795), .ZN(n2782) );
  INV_X1 U2574 ( .A(n70), .ZN(n2776) );
  OAI221_X1 U2575 ( .B1(n2756), .B2(n2418), .C1(n2724), .C2(n2419), .A(n2796), 
        .ZN(n70) );
  AOI22_X1 U2576 ( .A1(n2074), .A2(n2422), .B1(n2421), .B2(n2721), .ZN(n2796)
         );
  OAI22_X1 U2577 ( .A1(n5066), .A2(n17002), .B1(n2797), .B2(n17005), .ZN(
        U449_Z_0) );
  OAI22_X1 U2578 ( .A1(n5065), .A2(n16997), .B1(n2797), .B2(n17000), .ZN(
        U448_Z_0) );
  OAI22_X1 U2579 ( .A1(n5297), .A2(n17039), .B1(n2797), .B2(n17042), .ZN(
        U447_Z_0) );
  OAI22_X1 U2580 ( .A1(n5276), .A2(n17034), .B1(n2797), .B2(n17037), .ZN(
        U446_Z_0) );
  OAI22_X1 U2581 ( .A1(n5064), .A2(n17029), .B1(n2797), .B2(n17032), .ZN(
        U445_Z_0) );
  OAI22_X1 U2582 ( .A1(n5187), .A2(n17024), .B1(n2797), .B2(n17027), .ZN(
        U444_Z_0) );
  OAI22_X1 U2583 ( .A1(n5063), .A2(n17019), .B1(n2797), .B2(n17022), .ZN(
        U443_Z_0) );
  OAI22_X1 U2584 ( .A1(n5216), .A2(n17014), .B1(n2797), .B2(n17017), .ZN(
        U442_Z_0) );
  OAI22_X1 U2585 ( .A1(n5323), .A2(n17044), .B1(n2797), .B2(n17047), .ZN(
        U441_Z_0) );
  OAI22_X1 U2586 ( .A1(n5352), .A2(n17049), .B1(n2797), .B2(n17052), .ZN(
        U440_Z_0) );
  OAI22_X1 U2587 ( .A1(n5381), .A2(n17054), .B1(n2797), .B2(n17057), .ZN(
        U439_Z_0) );
  OAI22_X1 U2588 ( .A1(n5410), .A2(n17059), .B1(n2797), .B2(n17062), .ZN(
        U438_Z_0) );
  OAI22_X1 U2589 ( .A1(n5439), .A2(n17064), .B1(n2797), .B2(n17067), .ZN(
        U437_Z_0) );
  OAI22_X1 U2590 ( .A1(n5468), .A2(n17069), .B1(n2797), .B2(n17072), .ZN(
        U436_Z_0) );
  OAI22_X1 U2591 ( .A1(n5062), .A2(n17074), .B1(n2797), .B2(n17077), .ZN(
        U435_Z_0) );
  OAI22_X1 U2592 ( .A1(n5492), .A2(n17079), .B1(n2797), .B2(n17082), .ZN(
        U434_Z_0) );
  AOI221_X1 U2594 ( .B1(n17006), .B2(n2249), .C1(n16672), .C2(n17010), .A(
        n2289), .ZN(n2799) );
  AND2_X1 U2595 ( .A1(n2800), .A2(n1657), .ZN(n2289) );
  OAI22_X1 U2596 ( .A1(n16993), .A2(n5812), .B1(n2131), .B2(n2801), .ZN(n2800)
         );
  INV_X1 U2597 ( .A(n5812), .ZN(n2801) );
  AOI221_X1 U2598 ( .B1(n2464), .B2(n2074), .C1(n2720), .C2(n2469), .A(n2802), 
        .ZN(n64) );
  INV_X1 U2599 ( .A(n2803), .ZN(n2802) );
  AOI22_X1 U2600 ( .A1(n2468), .A2(n2749), .B1(n2465), .B2(n2721), .ZN(n2803)
         );
  NAND3_X1 U2601 ( .A1(n5812), .A2(n16994), .A3(n1690), .ZN(n2798) );
  INV_X1 U2602 ( .A(n1657), .ZN(n1690) );
  NAND4_X1 U2603 ( .A1(n2804), .A2(n2805), .A3(n2806), .A4(n2807), .ZN(n1657)
         );
  AOI222_X1 U2604 ( .A1(n16974), .A2(vis_msp_o[16]), .B1(n16971), .B2(n2809), 
        .C1(n16968), .C2(vis_psp_o[16]), .ZN(n2807) );
  AOI222_X1 U2606 ( .A1(n16983), .A2(vis_r14_o[18]), .B1(n16965), .B2(
        vis_r12_o[18]), .C1(n16986), .C2(vis_r11_o[18]), .ZN(n2806) );
  AOI222_X1 U2609 ( .A1(n16980), .A2(vis_r9_o[18]), .B1(n16962), .B2(
        vis_r10_o[18]), .C1(n16959), .C2(vis_r8_o[18]), .ZN(n2805) );
  AOI22_X1 U2611 ( .A1(n16977), .A2(n2795), .B1(n16955), .B2(n2817), .ZN(n2804) );
  XOR2_X1 U2613 ( .A(n16990), .B(n2818), .Z(n5812) );
  AOI221_X1 U2614 ( .B1(n16989), .B2(n2249), .C1(n2198), .C2(n2819), .A(n2732), 
        .ZN(n2818) );
  OAI22_X1 U2615 ( .A1(n5087), .A2(n17002), .B1(n2820), .B2(n17005), .ZN(
        U433_Z_0) );
  OAI22_X1 U2616 ( .A1(n5086), .A2(n16997), .B1(n2820), .B2(n17000), .ZN(
        U432_Z_0) );
  OAI22_X1 U2617 ( .A1(n5298), .A2(n17039), .B1(n2820), .B2(n17042), .ZN(
        U431_Z_0) );
  OAI22_X1 U2618 ( .A1(n5277), .A2(n17034), .B1(n2820), .B2(n17037), .ZN(
        U430_Z_0) );
  OAI22_X1 U2619 ( .A1(n5085), .A2(n17029), .B1(n2820), .B2(n17032), .ZN(
        U429_Z_0) );
  OAI22_X1 U2620 ( .A1(n5188), .A2(n17024), .B1(n2820), .B2(n17027), .ZN(
        U428_Z_0) );
  OAI22_X1 U2621 ( .A1(n5084), .A2(n17019), .B1(n2820), .B2(n17022), .ZN(
        U427_Z_0) );
  OAI22_X1 U2622 ( .A1(n5217), .A2(n17014), .B1(n2820), .B2(n17017), .ZN(
        U426_Z_0) );
  OAI22_X1 U2623 ( .A1(n5324), .A2(n17044), .B1(n2820), .B2(n17047), .ZN(
        U425_Z_0) );
  OAI22_X1 U2624 ( .A1(n5353), .A2(n17049), .B1(n2820), .B2(n17052), .ZN(
        U424_Z_0) );
  OAI22_X1 U2625 ( .A1(n5382), .A2(n17054), .B1(n2820), .B2(n17057), .ZN(
        U423_Z_0) );
  OAI22_X1 U2626 ( .A1(n5411), .A2(n17059), .B1(n2820), .B2(n17062), .ZN(
        U422_Z_0) );
  OAI22_X1 U2627 ( .A1(n5440), .A2(n17064), .B1(n2820), .B2(n17067), .ZN(
        U421_Z_0) );
  OAI22_X1 U2628 ( .A1(n5469), .A2(n17069), .B1(n2820), .B2(n17072), .ZN(
        U420_Z_0) );
  OAI22_X1 U2629 ( .A1(n5083), .A2(n17074), .B1(n2820), .B2(n17077), .ZN(
        U419_Z_0) );
  OAI22_X1 U2630 ( .A1(n5493), .A2(n17079), .B1(n2820), .B2(n17082), .ZN(
        U418_Z_0) );
  AOI222_X1 U2632 ( .A1(n17007), .A2(n2258), .B1(n2823), .B2(n2824), .C1(
        n16710), .C2(n17009), .ZN(n2822) );
  NAND3_X1 U2633 ( .A1(n2131), .A2(n1658), .A3(n5811), .ZN(n2824) );
  OAI21_X1 U2634 ( .B1(n16993), .B2(n1691), .A(n2825), .ZN(n2823) );
  OAI21_X1 U2635 ( .B1(n16994), .B2(n1658), .A(n5811), .ZN(n2825) );
  XOR2_X1 U2636 ( .A(n16990), .B(n2826), .Z(n5811) );
  AOI221_X1 U2637 ( .B1(n16989), .B2(n2258), .C1(n2198), .C2(n2827), .A(n2732), 
        .ZN(n2826) );
  INV_X1 U2638 ( .A(n1658), .ZN(n1691) );
  NAND4_X1 U2639 ( .A1(n2828), .A2(n2829), .A3(n2830), .A4(n2831), .ZN(n1658)
         );
  AOI222_X1 U2640 ( .A1(n16974), .A2(vis_msp_o[15]), .B1(n16971), .B2(n2833), 
        .C1(n16968), .C2(vis_psp_o[15]), .ZN(n2831) );
  AOI222_X1 U2642 ( .A1(n16983), .A2(vis_r14_o[17]), .B1(n16965), .B2(
        vis_r12_o[17]), .C1(n16986), .C2(vis_r11_o[17]), .ZN(n2830) );
  AOI222_X1 U2645 ( .A1(n16980), .A2(vis_r9_o[17]), .B1(n16962), .B2(
        vis_r10_o[17]), .C1(n16959), .C2(vis_r8_o[17]), .ZN(n2829) );
  AOI22_X1 U2647 ( .A1(n16977), .A2(n2817), .B1(n16955), .B2(n2841), .ZN(n2828) );
  INV_X1 U2649 ( .A(n66), .ZN(n2821) );
  OAI221_X1 U2650 ( .B1(n2756), .B2(n2472), .C1(n2724), .C2(n2473), .A(n2842), 
        .ZN(n66) );
  AOI22_X1 U2651 ( .A1(n2074), .A2(n2005), .B1(n2003), .B2(n2721), .ZN(n2842)
         );
  OAI22_X1 U2652 ( .A1(n5073), .A2(n17001), .B1(n2843), .B2(n17005), .ZN(
        U415_Z_0) );
  OAI22_X1 U2653 ( .A1(n5072), .A2(n16996), .B1(n2843), .B2(n17000), .ZN(
        U414_Z_0) );
  OAI22_X1 U2654 ( .A1(n5299), .A2(n17038), .B1(n2843), .B2(n17042), .ZN(
        U413_Z_0) );
  OAI22_X1 U2655 ( .A1(n5278), .A2(n17033), .B1(n2843), .B2(n17037), .ZN(
        U412_Z_0) );
  OAI22_X1 U2656 ( .A1(n5071), .A2(n17028), .B1(n2843), .B2(n17032), .ZN(
        U411_Z_0) );
  OAI22_X1 U2657 ( .A1(n5189), .A2(n17023), .B1(n2843), .B2(n17027), .ZN(
        U410_Z_0) );
  OAI22_X1 U2658 ( .A1(n5070), .A2(n17018), .B1(n2843), .B2(n17022), .ZN(
        U409_Z_0) );
  OAI22_X1 U2659 ( .A1(n5218), .A2(n17013), .B1(n2843), .B2(n17017), .ZN(
        U408_Z_0) );
  OAI22_X1 U2660 ( .A1(n5325), .A2(n17043), .B1(n2843), .B2(n17047), .ZN(
        U407_Z_0) );
  OAI22_X1 U2661 ( .A1(n5354), .A2(n17048), .B1(n2843), .B2(n17052), .ZN(
        U406_Z_0) );
  OAI22_X1 U2662 ( .A1(n5383), .A2(n17053), .B1(n2843), .B2(n17057), .ZN(
        U405_Z_0) );
  OAI22_X1 U2663 ( .A1(n5412), .A2(n17058), .B1(n2843), .B2(n17062), .ZN(
        U404_Z_0) );
  OAI22_X1 U2664 ( .A1(n5441), .A2(n17063), .B1(n2843), .B2(n17067), .ZN(
        U403_Z_0) );
  OAI22_X1 U2665 ( .A1(n5470), .A2(n17068), .B1(n2843), .B2(n17072), .ZN(
        U402_Z_0) );
  OAI22_X1 U2666 ( .A1(n5069), .A2(n17073), .B1(n2843), .B2(n17077), .ZN(
        U401_Z_0) );
  OAI22_X1 U2667 ( .A1(n5494), .A2(n17078), .B1(n2843), .B2(n17082), .ZN(
        U400_Z_0) );
  AOI221_X1 U2669 ( .B1(n17006), .B2(n17), .C1(n16711), .C2(n17010), .A(n2847), 
        .ZN(n2846) );
  INV_X1 U2670 ( .A(n2307), .ZN(n2847) );
  NAND2_X1 U2671 ( .A1(n2848), .A2(n1660), .ZN(n2307) );
  OAI22_X1 U2672 ( .A1(n16992), .A2(n5810), .B1(n2131), .B2(n2849), .ZN(n2848)
         );
  INV_X1 U2673 ( .A(n5810), .ZN(n2849) );
  INV_X1 U2674 ( .A(n68), .ZN(n2845) );
  OAI221_X1 U2675 ( .B1(n2517), .B2(n2723), .C1(n2724), .C2(n2516), .A(n2850), 
        .ZN(n68) );
  AOI22_X1 U2676 ( .A1(n2023), .A2(n2720), .B1(n2019), .B2(n2721), .ZN(n2850)
         );
  INV_X1 U2677 ( .A(n2749), .ZN(n2724) );
  NAND3_X1 U2678 ( .A1(n5810), .A2(n16994), .A3(n1692), .ZN(n2844) );
  INV_X1 U2679 ( .A(n1660), .ZN(n1692) );
  NAND4_X1 U2680 ( .A1(n2851), .A2(n2852), .A3(n2853), .A4(n2854), .ZN(n1660)
         );
  AOI222_X1 U2681 ( .A1(n16974), .A2(vis_msp_o[14]), .B1(n16971), .B2(n2856), 
        .C1(n16968), .C2(vis_psp_o[14]), .ZN(n2854) );
  AOI222_X1 U2683 ( .A1(n16983), .A2(vis_r14_o[16]), .B1(n16965), .B2(
        vis_r12_o[16]), .C1(n16986), .C2(vis_r11_o[16]), .ZN(n2853) );
  AOI222_X1 U2686 ( .A1(n16980), .A2(vis_r9_o[16]), .B1(n16963), .B2(
        vis_r10_o[16]), .C1(n16959), .C2(vis_r8_o[16]), .ZN(n2852) );
  AOI22_X1 U2688 ( .A1(n16977), .A2(n2841), .B1(n16955), .B2(n1163), .ZN(n2851) );
  XOR2_X1 U2690 ( .A(n16990), .B(n2864), .Z(n5810) );
  AOI221_X1 U2691 ( .B1(n16989), .B2(n17), .C1(n2198), .C2(n2865), .A(n2732), 
        .ZN(n2864) );
  NOR2_X1 U2692 ( .A1(n2055), .A2(n71), .ZN(n2696) );
  OAI22_X1 U2693 ( .A1(n5107), .A2(n17001), .B1(n2866), .B2(n17005), .ZN(
        U399_Z_0) );
  OAI22_X1 U2694 ( .A1(n5106), .A2(n16996), .B1(n2866), .B2(n17000), .ZN(
        U398_Z_0) );
  OAI22_X1 U2695 ( .A1(n5300), .A2(n17038), .B1(n2866), .B2(n17042), .ZN(
        U397_Z_0) );
  OAI22_X1 U2696 ( .A1(n5279), .A2(n17033), .B1(n2866), .B2(n17037), .ZN(
        U396_Z_0) );
  OAI22_X1 U2697 ( .A1(n5105), .A2(n17028), .B1(n2866), .B2(n17032), .ZN(
        U395_Z_0) );
  OAI22_X1 U2698 ( .A1(n5190), .A2(n17023), .B1(n2866), .B2(n17027), .ZN(
        U394_Z_0) );
  OAI22_X1 U2699 ( .A1(n5104), .A2(n17018), .B1(n2866), .B2(n17022), .ZN(
        U393_Z_0) );
  OAI22_X1 U2700 ( .A1(n5219), .A2(n17013), .B1(n2866), .B2(n17017), .ZN(
        U392_Z_0) );
  OAI22_X1 U2701 ( .A1(n5326), .A2(n17043), .B1(n2866), .B2(n17047), .ZN(
        U391_Z_0) );
  OAI22_X1 U2702 ( .A1(n5355), .A2(n17048), .B1(n2866), .B2(n17052), .ZN(
        U390_Z_0) );
  OAI22_X1 U2703 ( .A1(n5384), .A2(n17053), .B1(n2866), .B2(n17057), .ZN(
        U389_Z_0) );
  OAI22_X1 U2704 ( .A1(n5413), .A2(n17058), .B1(n2866), .B2(n17062), .ZN(
        U388_Z_0) );
  OAI22_X1 U2705 ( .A1(n5442), .A2(n17063), .B1(n2866), .B2(n17067), .ZN(
        U387_Z_0) );
  OAI22_X1 U2706 ( .A1(n5471), .A2(n17068), .B1(n2866), .B2(n17072), .ZN(
        U386_Z_0) );
  OAI22_X1 U2707 ( .A1(n5103), .A2(n17073), .B1(n2866), .B2(n17077), .ZN(
        U385_Z_0) );
  OAI22_X1 U2708 ( .A1(n5495), .A2(n17078), .B1(n2866), .B2(n17082), .ZN(
        U384_Z_0) );
  AOI221_X1 U2710 ( .B1(n16658), .B2(n17009), .C1(n17008), .C2(n2253), .A(n135), .ZN(n2867) );
  OAI221_X1 U2711 ( .B1(n2868), .B2(n2090), .C1(n2869), .C2(n2088), .A(n2870), 
        .ZN(n135) );
  AOI221_X1 U2712 ( .B1(n2093), .B2(n2871), .C1(n2094), .C2(n2872), .A(n2873), 
        .ZN(n2870) );
  OAI211_X1 U2713 ( .C1(n2874), .C2(n2875), .A(n2876), .B(n2877), .ZN(n2094)
         );
  AOI222_X1 U2714 ( .A1(sub_2068_A_22_), .A2(n2878), .B1(hrdata_i[22]), .B2(
        n2879), .C1(n16787), .C2(n2881), .ZN(n2877) );
  AOI22_X1 U2716 ( .A1(n2882), .A2(n2883), .B1(n16645), .B2(n2344), .ZN(n2876)
         );
  OAI221_X1 U2717 ( .B1(n1896), .B2(n2885), .C1(n5053), .C2(n2886), .A(n2887), 
        .ZN(n2883) );
  AOI222_X1 U2718 ( .A1(n1890), .A2(n2888), .B1(n1191), .B2(n2889), .C1(n1887), 
        .C2(n2890), .ZN(n2887) );
  NAND4_X1 U2720 ( .A1(n2891), .A2(n2892), .A3(n2893), .A4(n2894), .ZN(n2093)
         );
  AOI221_X1 U2721 ( .B1(n407), .B2(n2895), .C1(n2882), .C2(n2896), .A(n2897), 
        .ZN(n2894) );
  OAI221_X1 U2722 ( .B1(n5151), .B2(n2898), .C1(n5157), .C2(n2899), .A(n2900), 
        .ZN(n2896) );
  AOI22_X1 U2723 ( .A1(n1897), .A2(n2901), .B1(n1893), .B2(n2902), .ZN(n2900)
         );
  INV_X1 U2724 ( .A(n426), .ZN(n407) );
  OAI211_X1 U2725 ( .C1(n2903), .C2(n1372), .A(n2904), .B(n2905), .ZN(n426) );
  NAND3_X1 U2726 ( .A1(n2906), .A2(n1372), .A3(n2907), .ZN(n2904) );
  OAI22_X1 U2727 ( .A1(n2908), .A2(n2909), .B1(n2910), .B2(n2911), .ZN(n2906)
         );
  AOI22_X1 U2728 ( .A1(n2912), .A2(n2352), .B1(n16645), .B2(n2388), .ZN(n2893)
         );
  AOI222_X1 U2729 ( .A1(hrdata_i[14]), .A2(n2879), .B1(n2913), .B2(n2914), 
        .C1(n2915), .C2(n2916), .ZN(n2892) );
  AOI22_X1 U2730 ( .A1(n16787), .A2(n2917), .B1(sub_2068_A_14_), .B2(n2878), 
        .ZN(n2891) );
  INV_X1 U2732 ( .A(n2546), .ZN(n2088) );
  OAI211_X1 U2733 ( .C1(n2918), .C2(n1145), .A(n2919), .B(n2920), .ZN(n2546)
         );
  AOI211_X1 U2734 ( .C1(n2921), .C2(n2922), .A(n2923), .B(n2897), .ZN(n2920)
         );
  AOI21_X1 U2735 ( .B1(n2924), .B2(n2925), .A(n2926), .ZN(n2923) );
  AOI222_X1 U2736 ( .A1(n1887), .A2(n2927), .B1(n2928), .B2(n1189), .C1(n1191), 
        .C2(n2929), .ZN(n2925) );
  NOR2_X1 U2737 ( .A1(n5503), .A2(n2930), .ZN(n2928) );
  AOI222_X1 U2738 ( .A1(n1893), .A2(n2931), .B1(n1890), .B2(n2932), .C1(n1897), 
        .C2(n2933), .ZN(n2924) );
  INV_X1 U2739 ( .A(n2373), .ZN(n2921) );
  OAI22_X1 U2740 ( .A1(n2313), .A2(n2934), .B1(n2935), .B2(n2936), .ZN(n2373)
         );
  INV_X1 U2741 ( .A(n2934), .ZN(n2936) );
  AOI22_X1 U2742 ( .A1(n2937), .A2(n2337), .B1(n2938), .B2(n16789), .ZN(n2935)
         );
  INV_X1 U2743 ( .A(n2332), .ZN(n2938) );
  AOI22_X1 U2744 ( .A1(n2939), .A2(n2940), .B1(n2941), .B2(n2942), .ZN(n2934)
         );
  INV_X1 U2745 ( .A(hrdata_i[30]), .ZN(n1145) );
  INV_X1 U2746 ( .A(n2545), .ZN(n2090) );
  NAND3_X1 U2747 ( .A1(n2943), .A2(n2944), .A3(n2945), .ZN(n2545) );
  AOI221_X1 U2748 ( .B1(n16787), .B2(n2946), .C1(sub_2068_A_6_), .C2(n2878), 
        .A(n2947), .ZN(n2945) );
  OAI22_X1 U2749 ( .A1(n2918), .A2(n397), .B1(n4798), .B2(n2948), .ZN(n2947)
         );
  INV_X1 U2750 ( .A(hrdata_i[6]), .ZN(n397) );
  AOI22_X1 U2752 ( .A1(n2882), .A2(n2949), .B1(n16645), .B2(n2325), .ZN(n2944)
         );
  OAI221_X1 U2753 ( .B1(n1885), .B2(n2898), .C1(n5518), .C2(n2899), .A(n2950), 
        .ZN(n2949) );
  AOI22_X1 U2754 ( .A1(n1897), .A2(n2951), .B1(n1893), .B2(n2952), .ZN(n2950)
         );
  AOI22_X1 U2756 ( .A1(n2912), .A2(n2329), .B1(n2913), .B2(n2953), .ZN(n2943)
         );
  INV_X1 U2757 ( .A(n2954), .ZN(n2868) );
  NAND3_X1 U2758 ( .A1(n5809), .A2(n16994), .A3(n1693), .ZN(n2285) );
  INV_X1 U2759 ( .A(n1663), .ZN(n1693) );
  NAND2_X1 U2760 ( .A1(n2955), .A2(n1663), .ZN(n2305) );
  NAND4_X1 U2761 ( .A1(n2956), .A2(n2957), .A3(n2958), .A4(n2959), .ZN(n1663)
         );
  AOI222_X1 U2762 ( .A1(n16958), .A2(vis_r8_o[14]), .B1(n16976), .B2(n2961), 
        .C1(n16981), .C2(vis_r9_o[14]), .ZN(n2959) );
  AOI222_X1 U2764 ( .A1(n16985), .A2(vis_r11_o[14]), .B1(n16970), .B2(n2964), 
        .C1(n16984), .C2(vis_r14_o[14]), .ZN(n2958) );
  AOI222_X1 U2767 ( .A1(n16967), .A2(vis_psp_o[12]), .B1(n16963), .B2(
        vis_r10_o[14]), .C1(n16975), .C2(vis_msp_o[12]), .ZN(n2957) );
  AOI22_X1 U2769 ( .A1(n16966), .A2(vis_r12_o[14]), .B1(n2970), .B2(n16956), 
        .ZN(n2956) );
  OAI22_X1 U2770 ( .A1(n16993), .A2(n5809), .B1(n2131), .B2(n2971), .ZN(n2955)
         );
  INV_X1 U2771 ( .A(n5809), .ZN(n2971) );
  XOR2_X1 U2772 ( .A(n2169), .B(n2972), .Z(n5809) );
  AOI221_X1 U2773 ( .B1(n16989), .B2(n2253), .C1(n2198), .C2(n795), .A(n2732), 
        .ZN(n2972) );
  OAI22_X1 U2774 ( .A1(n5599), .A2(n17001), .B1(n2973), .B2(n17005), .ZN(
        U383_Z_0) );
  OAI22_X1 U2775 ( .A1(n5598), .A2(n16996), .B1(n2973), .B2(n17000), .ZN(
        U382_Z_0) );
  OAI22_X1 U2776 ( .A1(n5597), .A2(n17038), .B1(n2973), .B2(n17042), .ZN(
        U381_Z_0) );
  OAI22_X1 U2777 ( .A1(n5596), .A2(n17033), .B1(n2973), .B2(n17037), .ZN(
        U380_Z_0) );
  OAI22_X1 U2778 ( .A1(n5134), .A2(n17028), .B1(n2973), .B2(n17032), .ZN(
        U379_Z_0) );
  OAI22_X1 U2779 ( .A1(n5191), .A2(n17023), .B1(n2973), .B2(n17027), .ZN(
        U378_Z_0) );
  OAI22_X1 U2780 ( .A1(n5133), .A2(n17018), .B1(n2973), .B2(n17022), .ZN(
        U377_Z_0) );
  OAI22_X1 U2781 ( .A1(n5220), .A2(n17013), .B1(n2973), .B2(n17017), .ZN(
        U376_Z_0) );
  OAI22_X1 U2782 ( .A1(n5327), .A2(n17043), .B1(n2973), .B2(n17047), .ZN(
        U375_Z_0) );
  OAI22_X1 U2783 ( .A1(n5356), .A2(n17048), .B1(n2973), .B2(n17052), .ZN(
        U374_Z_0) );
  OAI22_X1 U2784 ( .A1(n5385), .A2(n17053), .B1(n2973), .B2(n17057), .ZN(
        U373_Z_0) );
  OAI22_X1 U2785 ( .A1(n5414), .A2(n17058), .B1(n2973), .B2(n17062), .ZN(
        U372_Z_0) );
  OAI22_X1 U2786 ( .A1(n5443), .A2(n17063), .B1(n2973), .B2(n17067), .ZN(
        U371_Z_0) );
  OAI22_X1 U2787 ( .A1(n5472), .A2(n17068), .B1(n2973), .B2(n17072), .ZN(
        U370_Z_0) );
  OAI22_X1 U2788 ( .A1(n5132), .A2(n17073), .B1(n2973), .B2(n17077), .ZN(
        U369_Z_0) );
  OAI22_X1 U2789 ( .A1(n5496), .A2(n17078), .B1(n2973), .B2(n17082), .ZN(
        U368_Z_0) );
  AOI221_X1 U2791 ( .B1(n16679), .B2(n17009), .C1(n17008), .C2(n2259), .A(
        n2976), .ZN(n2975) );
  INV_X1 U2792 ( .A(n118), .ZN(n2976) );
  AOI221_X1 U2793 ( .B1(n2954), .B2(n2415), .C1(n2414), .C2(n2977), .A(n2978), 
        .ZN(n118) );
  INV_X1 U2794 ( .A(n2979), .ZN(n2978) );
  AOI221_X1 U2795 ( .B1(n2411), .B2(n2871), .C1(n2410), .C2(n2872), .A(n2873), 
        .ZN(n2979) );
  OAI221_X1 U2796 ( .B1(n5625), .B2(n16685), .C1(n2981), .C2(n270), .A(n2982), 
        .ZN(n2410) );
  AOI222_X1 U2797 ( .A1(hrdata_i[21]), .A2(n2879), .B1(n16645), .B2(n2345), 
        .C1(n2912), .C2(n2357), .ZN(n2982) );
  NAND3_X1 U2799 ( .A1(n2983), .A2(n2984), .A3(n2985), .ZN(n2411) );
  AOI221_X1 U2800 ( .B1(n16787), .B2(n2986), .C1(sub_2068_A_13_), .C2(n2878), 
        .A(n2987), .ZN(n2985) );
  OAI22_X1 U2801 ( .A1(n2918), .A2(n382), .B1(n244), .B2(n2948), .ZN(n2987) );
  INV_X1 U2802 ( .A(hrdata_i[13]), .ZN(n382) );
  AOI22_X1 U2804 ( .A1(n2895), .A2(n410), .B1(n16645), .B2(n2988), .ZN(n2984)
         );
  OAI211_X1 U2805 ( .C1(n1067), .C2(n2989), .A(n5229), .B(n4965), .ZN(n410) );
  AOI211_X1 U2806 ( .C1(n2908), .C2(n2990), .A(n2991), .B(n1370), .ZN(n2989)
         );
  OAI21_X1 U2807 ( .B1(n2908), .B2(n2992), .A(n2907), .ZN(n2991) );
  AOI22_X1 U2808 ( .A1(n2993), .A2(n2994), .B1(n2909), .B2(n2995), .ZN(n2992)
         );
  OAI21_X1 U2809 ( .B1(n2996), .B2(n2910), .A(n2997), .ZN(n2990) );
  AOI22_X1 U2810 ( .A1(n2912), .A2(n2353), .B1(n2913), .B2(n4751), .ZN(n2983)
         );
  OAI221_X1 U2811 ( .B1(n2998), .B2(n2374), .C1(n2918), .C2(n1144), .A(n2999), 
        .ZN(n2414) );
  INV_X1 U2812 ( .A(n3000), .ZN(n2999) );
  OAI21_X1 U2813 ( .B1(n3001), .B2(n3002), .A(n3003), .ZN(n3000) );
  INV_X1 U2814 ( .A(hrdata_i[29]), .ZN(n1144) );
  OAI221_X1 U2815 ( .B1(n2337), .B2(n2336), .C1(n16788), .C2(n3004), .A(n3002), 
        .ZN(n2374) );
  AOI22_X1 U2816 ( .A1(n3005), .A2(n2940), .B1(n2941), .B2(n3006), .ZN(n3002)
         );
  NAND2_X1 U2817 ( .A1(n3007), .A2(n3008), .ZN(n2415) );
  AOI221_X1 U2818 ( .B1(n16645), .B2(n2326), .C1(n2912), .C2(n2330), .A(n3009), 
        .ZN(n3008) );
  OAI22_X1 U2819 ( .A1(n3010), .A2(n2948), .B1(n5533), .B2(n3011), .ZN(n3009)
         );
  AOI222_X1 U2820 ( .A1(sub_2068_A_5_), .A2(n2878), .B1(hrdata_i[5]), .B2(
        n2879), .C1(n16787), .C2(n3012), .ZN(n3007) );
  INV_X1 U2822 ( .A(n2308), .ZN(n2974) );
  NOR3_X1 U2823 ( .A1(n3013), .A2(n2501), .A3(n1664), .ZN(n2308) );
  NAND2_X1 U2824 ( .A1(n3014), .A2(n1664), .ZN(n2306) );
  NAND4_X1 U2825 ( .A1(n3015), .A2(n3016), .A3(n3017), .A4(n3018), .ZN(n1664)
         );
  AOI222_X1 U2826 ( .A1(n16958), .A2(vis_r8_o[13]), .B1(n16976), .B2(n2970), 
        .C1(n16981), .C2(vis_r9_o[13]), .ZN(n3018) );
  AOI222_X1 U2829 ( .A1(n16961), .A2(vis_r10_o[13]), .B1(n16970), .B2(n3022), 
        .C1(n16987), .C2(vis_r11_o[13]), .ZN(n3017) );
  AOI222_X1 U2831 ( .A1(n16974), .A2(vis_msp_o[11]), .B1(n16984), .B2(
        vis_r14_o[13]), .C1(n16964), .C2(vis_r12_o[13]), .ZN(n3016) );
  AOI22_X1 U2834 ( .A1(n16969), .A2(vis_psp_o[11]), .B1(n3028), .B2(n16956), 
        .ZN(n3015) );
  OAI22_X1 U2835 ( .A1(n16992), .A2(n5808), .B1(n2131), .B2(n3013), .ZN(n3014)
         );
  INV_X1 U2836 ( .A(n5808), .ZN(n3013) );
  XOR2_X1 U2837 ( .A(n2169), .B(n3029), .Z(n5808) );
  AOI221_X1 U2838 ( .B1(n16989), .B2(n2259), .C1(n2198), .C2(n16656), .A(n2732), .ZN(n3029) );
  OAI22_X1 U2839 ( .A1(n5131), .A2(n17001), .B1(n3030), .B2(n17005), .ZN(
        U367_Z_0) );
  OAI22_X1 U2840 ( .A1(n5130), .A2(n16996), .B1(n3030), .B2(n17000), .ZN(
        U366_Z_0) );
  OAI22_X1 U2841 ( .A1(n5301), .A2(n17038), .B1(n3030), .B2(n17042), .ZN(
        U365_Z_0) );
  OAI22_X1 U2842 ( .A1(n5280), .A2(n17033), .B1(n3030), .B2(n17037), .ZN(
        U364_Z_0) );
  OAI22_X1 U2843 ( .A1(n5129), .A2(n17028), .B1(n3030), .B2(n17032), .ZN(
        U363_Z_0) );
  OAI22_X1 U2844 ( .A1(n5192), .A2(n17023), .B1(n3030), .B2(n17027), .ZN(
        U362_Z_0) );
  OAI22_X1 U2845 ( .A1(n5128), .A2(n17018), .B1(n3030), .B2(n17022), .ZN(
        U361_Z_0) );
  OAI22_X1 U2846 ( .A1(n5221), .A2(n17013), .B1(n3030), .B2(n17017), .ZN(
        U360_Z_0) );
  OAI22_X1 U2847 ( .A1(n5328), .A2(n17043), .B1(n3030), .B2(n17047), .ZN(
        U359_Z_0) );
  OAI22_X1 U2848 ( .A1(n5357), .A2(n17048), .B1(n3030), .B2(n17052), .ZN(
        U358_Z_0) );
  OAI22_X1 U2849 ( .A1(n5386), .A2(n17053), .B1(n3030), .B2(n17057), .ZN(
        U357_Z_0) );
  OAI22_X1 U2850 ( .A1(n5415), .A2(n17058), .B1(n3030), .B2(n17062), .ZN(
        U356_Z_0) );
  OAI22_X1 U2851 ( .A1(n5444), .A2(n17063), .B1(n3030), .B2(n17067), .ZN(
        U355_Z_0) );
  OAI22_X1 U2852 ( .A1(n5473), .A2(n17068), .B1(n3030), .B2(n17072), .ZN(
        U354_Z_0) );
  OAI22_X1 U2853 ( .A1(n5127), .A2(n17073), .B1(n3030), .B2(n17077), .ZN(
        U353_Z_0) );
  OAI22_X1 U2854 ( .A1(n5497), .A2(n17078), .B1(n3030), .B2(n17082), .ZN(
        U352_Z_0) );
  AOI221_X1 U2856 ( .B1(n17006), .B2(n2247), .C1(n16653), .C2(n17010), .A(
        n2055), .ZN(n3032) );
  OAI221_X1 U2857 ( .B1(n3033), .B2(n5807), .C1(n16995), .C2(n1665), .A(n3034), 
        .ZN(n3031) );
  NAND3_X1 U2858 ( .A1(n2131), .A2(n1665), .A3(n5807), .ZN(n3034) );
  AOI221_X1 U2860 ( .B1(n16989), .B2(n2247), .C1(n2198), .C2(n2231), .A(n2732), 
        .ZN(n3035) );
  NOR2_X1 U2861 ( .A1(n1694), .A2(n16993), .ZN(n3033) );
  INV_X1 U2862 ( .A(n1665), .ZN(n1694) );
  NAND4_X1 U2863 ( .A1(n3036), .A2(n3037), .A3(n3038), .A4(n3039), .ZN(n1665)
         );
  AOI222_X1 U2864 ( .A1(n16974), .A2(vis_msp_o[10]), .B1(n16970), .B2(n3041), 
        .C1(n16968), .C2(vis_psp_o[10]), .ZN(n3039) );
  AOI222_X1 U2866 ( .A1(n16983), .A2(vis_r14_o[12]), .B1(n16966), .B2(
        vis_r12_o[12]), .C1(n16987), .C2(vis_r11_o[12]), .ZN(n3038) );
  AOI222_X1 U2869 ( .A1(n16980), .A2(vis_r9_o[12]), .B1(n16962), .B2(
        vis_r10_o[12]), .C1(n16959), .C2(vis_r8_o[12]), .ZN(n3037) );
  AOI22_X1 U2871 ( .A1(n16978), .A2(n3028), .B1(n16955), .B2(n3049), .ZN(n3036) );
  INV_X1 U2873 ( .A(n3050), .ZN(n136) );
  OAI221_X1 U2874 ( .B1(n2757), .B2(n3051), .C1(n2596), .C2(n2869), .A(n3052), 
        .ZN(n3050) );
  AOI221_X1 U2875 ( .B1(n2871), .B2(n2075), .C1(n2068), .C2(n2954), .A(n2873), 
        .ZN(n3052) );
  NAND3_X1 U2876 ( .A1(n3053), .A2(n3054), .A3(n3055), .ZN(n2068) );
  AOI221_X1 U2877 ( .B1(n16787), .B2(n3056), .C1(sub_2068_A_4_), .C2(n2878), 
        .A(n3057), .ZN(n3055) );
  OAI22_X1 U2878 ( .A1(n2918), .A2(n420), .B1(n4800), .B2(n2948), .ZN(n3057)
         );
  INV_X1 U2879 ( .A(hrdata_i[4]), .ZN(n420) );
  AOI22_X1 U2881 ( .A1(n3058), .A2(n3059), .B1(n16645), .B2(n2333), .ZN(n3054)
         );
  AOI22_X1 U2883 ( .A1(n2912), .A2(n2339), .B1(n2913), .B2(n3060), .ZN(n3053)
         );
  NAND3_X1 U2884 ( .A1(n3061), .A2(n3062), .A3(n3063), .ZN(n2075) );
  AOI221_X1 U2885 ( .B1(hrdata_i[12]), .B2(n2879), .C1(sub_2068_A_12_), .C2(
        n2878), .A(n3064), .ZN(n3063) );
  OAI22_X1 U2886 ( .A1(n5507), .A2(n16685), .B1(n4795), .B2(n2948), .ZN(n3064)
         );
  AOI22_X1 U2887 ( .A1(n417), .A2(n2895), .B1(n16645), .B2(n2387), .ZN(n3062)
         );
  INV_X1 U2888 ( .A(n412), .ZN(n417) );
  OAI21_X1 U2889 ( .B1(n3065), .B2(n3066), .A(n4965), .ZN(n412) );
  AOI211_X1 U2890 ( .C1(n1370), .C2(n2903), .A(n1067), .B(n3067), .ZN(n3065)
         );
  AOI211_X1 U2891 ( .C1(n3068), .C2(n2911), .A(n3069), .B(n1370), .ZN(n3067)
         );
  OAI21_X1 U2892 ( .B1(n3070), .B2(n2911), .A(n2907), .ZN(n3069) );
  AOI221_X1 U2893 ( .B1(n3071), .B2(n3072), .C1(n3073), .C2(n3074), .A(n3075), 
        .ZN(n3070) );
  NOR3_X1 U2894 ( .A1(n3076), .A2(n3073), .A3(n3077), .ZN(n3075) );
  OAI21_X1 U2895 ( .B1(n3078), .B2(n3079), .A(n3080), .ZN(n3074) );
  INV_X1 U2896 ( .A(n2997), .ZN(n3071) );
  OAI22_X1 U2897 ( .A1(n2993), .A2(n3081), .B1(n3082), .B2(n2909), .ZN(n3068)
         );
  INV_X1 U2898 ( .A(n3083), .ZN(n3082) );
  OAI21_X1 U2899 ( .B1(n2994), .B2(n3084), .A(n3085), .ZN(n3083) );
  AOI22_X1 U2900 ( .A1(n3086), .A2(n3087), .B1(n2995), .B2(n3088), .ZN(n3081)
         );
  AOI22_X1 U2901 ( .A1(n2912), .A2(n2385), .B1(n2913), .B2(n3089), .ZN(n3061)
         );
  AOI221_X1 U2902 ( .B1(n209), .B2(n2895), .C1(n2364), .C2(n2922), .A(n3090), 
        .ZN(n2596) );
  OAI21_X1 U2903 ( .B1(n1143), .B2(n2918), .A(n3003), .ZN(n3090) );
  INV_X1 U2904 ( .A(hrdata_i[28]), .ZN(n1143) );
  OAI22_X1 U2905 ( .A1(n3091), .A2(n3092), .B1(n2940), .B2(n3093), .ZN(n2364)
         );
  AOI22_X1 U2906 ( .A1(n16788), .A2(n3094), .B1(n2337), .B2(n3095), .ZN(n3093)
         );
  INV_X1 U2907 ( .A(n2066), .ZN(n2757) );
  OAI221_X1 U2908 ( .B1(n5618), .B2(n16685), .C1(n2981), .C2(n272), .A(n3096), 
        .ZN(n2066) );
  AOI222_X1 U2909 ( .A1(hrdata_i[20]), .A2(n2879), .B1(n16645), .B2(n2355), 
        .C1(n2912), .C2(n2350), .ZN(n3096) );
  OAI22_X1 U2911 ( .A1(n5569), .A2(n17001), .B1(n3097), .B2(n17005), .ZN(
        U349_Z_0) );
  OAI22_X1 U2912 ( .A1(n5568), .A2(n16996), .B1(n3097), .B2(n17000), .ZN(
        U348_Z_0) );
  OAI22_X1 U2913 ( .A1(n5567), .A2(n17038), .B1(n3097), .B2(n17042), .ZN(
        U347_Z_0) );
  OAI22_X1 U2914 ( .A1(n5566), .A2(n17033), .B1(n3097), .B2(n17037), .ZN(
        U346_Z_0) );
  OAI22_X1 U2915 ( .A1(n5565), .A2(n17028), .B1(n3097), .B2(n17032), .ZN(
        U345_Z_0) );
  OAI22_X1 U2916 ( .A1(n5564), .A2(n17023), .B1(n3097), .B2(n17027), .ZN(
        U344_Z_0) );
  OAI22_X1 U2917 ( .A1(n5563), .A2(n17018), .B1(n3097), .B2(n17022), .ZN(
        U343_Z_0) );
  OAI22_X1 U2918 ( .A1(n5562), .A2(n17013), .B1(n3097), .B2(n17017), .ZN(
        U342_Z_0) );
  OAI22_X1 U2919 ( .A1(n5561), .A2(n17043), .B1(n3097), .B2(n17047), .ZN(
        U341_Z_0) );
  OAI22_X1 U2920 ( .A1(n5560), .A2(n17048), .B1(n3097), .B2(n17052), .ZN(
        U340_Z_0) );
  OAI22_X1 U2921 ( .A1(n5559), .A2(n17053), .B1(n3097), .B2(n17057), .ZN(
        U339_Z_0) );
  OAI22_X1 U2922 ( .A1(n5558), .A2(n17058), .B1(n3097), .B2(n17062), .ZN(
        U338_Z_0) );
  OAI22_X1 U2923 ( .A1(n5557), .A2(n17063), .B1(n3097), .B2(n17067), .ZN(
        U337_Z_0) );
  OAI22_X1 U2924 ( .A1(n5556), .A2(n17068), .B1(n3097), .B2(n17072), .ZN(
        U336_Z_0) );
  OAI22_X1 U2925 ( .A1(n5555), .A2(n17073), .B1(n3097), .B2(n17077), .ZN(
        U335_Z_0) );
  OAI22_X1 U2926 ( .A1(n5554), .A2(n17078), .B1(n3097), .B2(n17082), .ZN(
        U334_Z_0) );
  INV_X1 U2928 ( .A(n3099), .ZN(n3098) );
  AOI221_X1 U2929 ( .B1(n16719), .B2(n17009), .C1(n17008), .C2(n2246), .A(n126), .ZN(n3099) );
  OAI221_X1 U2930 ( .B1(n3051), .B2(n2418), .C1(n2869), .C2(n2419), .A(n3100), 
        .ZN(n126) );
  AOI221_X1 U2931 ( .B1(n2421), .B2(n2871), .C1(n2422), .C2(n2954), .A(n2873), 
        .ZN(n3100) );
  NAND3_X1 U2932 ( .A1(n3101), .A2(n3102), .A3(n3103), .ZN(n2422) );
  AOI221_X1 U2933 ( .B1(n16787), .B2(n3104), .C1(sub_2068_A_3_), .C2(n2878), 
        .A(n3105), .ZN(n3103) );
  OAI22_X1 U2934 ( .A1(n2918), .A2(n423), .B1(n5536), .B2(n2948), .ZN(n3105)
         );
  INV_X1 U2935 ( .A(hrdata_i[3]), .ZN(n423) );
  AOI21_X1 U2937 ( .B1(n16645), .B2(n2334), .A(n3106), .ZN(n3102) );
  AOI22_X1 U2938 ( .A1(n2912), .A2(n2338), .B1(n2913), .B2(n3107), .ZN(n3101)
         );
  NAND3_X1 U2939 ( .A1(n3108), .A2(n3109), .A3(n3110), .ZN(n2421) );
  AOI222_X1 U2940 ( .A1(sub_2068_A_11_), .A2(n2878), .B1(hrdata_i[11]), .B2(
        n2879), .C1(n16787), .C2(n3111), .ZN(n3110) );
  AOI22_X1 U2942 ( .A1(n16645), .A2(n2386), .B1(n2912), .B2(n2384), .ZN(n3109)
         );
  INV_X1 U2943 ( .A(n3112), .ZN(n3108) );
  OAI22_X1 U2944 ( .A1(n3011), .A2(n5572), .B1(n2948), .B2(n5570), .ZN(n3112)
         );
  INV_X1 U2945 ( .A(n2623), .ZN(n2419) );
  OAI211_X1 U2946 ( .C1(n3113), .C2(n2368), .A(n3003), .B(n3114), .ZN(n2623)
         );
  INV_X1 U2947 ( .A(n3115), .ZN(n3114) );
  OAI22_X1 U2948 ( .A1(n3116), .A2(n3001), .B1(n1142), .B2(n2918), .ZN(n3115)
         );
  INV_X1 U2949 ( .A(hrdata_i[27]), .ZN(n1142) );
  OAI21_X1 U2950 ( .B1(n16788), .B2(n3117), .A(n3116), .ZN(n2368) );
  OAI221_X1 U2951 ( .B1(n3118), .B2(n3119), .C1(n3120), .C2(n16952), .A(n3122), 
        .ZN(n3116) );
  AOI21_X1 U2952 ( .B1(n2922), .B2(n2369), .A(n16645), .ZN(n3113) );
  INV_X1 U2953 ( .A(n2624), .ZN(n2418) );
  OAI211_X1 U2954 ( .C1(n3123), .C2(n2875), .A(n3124), .B(n3125), .ZN(n2624)
         );
  AOI222_X1 U2955 ( .A1(sub_2068_A_19_), .A2(n2878), .B1(hrdata_i[19]), .B2(
        n2879), .C1(n16787), .C2(n3126), .ZN(n3125) );
  AOI21_X1 U2957 ( .B1(n16645), .B2(n2354), .A(n2897), .ZN(n3124) );
  INV_X1 U2958 ( .A(n2356), .ZN(n3123) );
  AOI221_X1 U2959 ( .B1(n5820), .B2(n2131), .C1(n3127), .C2(n16992), .A(n1695), 
        .ZN(n2310) );
  INV_X1 U2960 ( .A(n3128), .ZN(n1695) );
  NOR3_X1 U2961 ( .A1(n3127), .A2(n2501), .A3(n3128), .ZN(n2309) );
  NAND4_X1 U2962 ( .A1(n3129), .A2(n3130), .A3(n3131), .A4(n3132), .ZN(n3128)
         );
  AOI222_X1 U2963 ( .A1(n16974), .A2(vis_msp_o[9]), .B1(n16970), .B2(n3134), 
        .C1(n16968), .C2(vis_psp_o[9]), .ZN(n3132) );
  AOI222_X1 U2965 ( .A1(n16983), .A2(vis_r14_o[11]), .B1(n16966), .B2(
        vis_r12_o[11]), .C1(n16987), .C2(vis_r11_o[11]), .ZN(n3131) );
  AOI222_X1 U2968 ( .A1(n16980), .A2(vis_r9_o[11]), .B1(n16963), .B2(
        vis_r10_o[11]), .C1(n16960), .C2(vis_r8_o[11]), .ZN(n3130) );
  AOI22_X1 U2970 ( .A1(n16978), .A2(n3049), .B1(n16956), .B2(n3142), .ZN(n3129) );
  INV_X1 U2972 ( .A(n5820), .ZN(n3127) );
  XOR2_X1 U2973 ( .A(n2169), .B(n3143), .Z(n5820) );
  AOI221_X1 U2974 ( .B1(n16989), .B2(n2246), .C1(n2198), .C2(n16817), .A(n2732), .ZN(n3143) );
  OAI22_X1 U2975 ( .A1(n5148), .A2(n17001), .B1(n3144), .B2(n17005), .ZN(
        U333_Z_0) );
  OAI22_X1 U2976 ( .A1(n5147), .A2(n16996), .B1(n3144), .B2(n17000), .ZN(
        U332_Z_0) );
  OAI22_X1 U2977 ( .A1(n5302), .A2(n17038), .B1(n3144), .B2(n17042), .ZN(
        U331_Z_0) );
  OAI22_X1 U2978 ( .A1(n5281), .A2(n17033), .B1(n3144), .B2(n17037), .ZN(
        U330_Z_0) );
  OAI22_X1 U2979 ( .A1(n5146), .A2(n17028), .B1(n3144), .B2(n17032), .ZN(
        U329_Z_0) );
  OAI22_X1 U2980 ( .A1(n5193), .A2(n17023), .B1(n3144), .B2(n17027), .ZN(
        U328_Z_0) );
  OAI22_X1 U2981 ( .A1(n5145), .A2(n17018), .B1(n3144), .B2(n17022), .ZN(
        U327_Z_0) );
  OAI22_X1 U2982 ( .A1(n5222), .A2(n17013), .B1(n3144), .B2(n17017), .ZN(
        U326_Z_0) );
  OAI22_X1 U2983 ( .A1(n5329), .A2(n17043), .B1(n3144), .B2(n17047), .ZN(
        U325_Z_0) );
  OAI22_X1 U2984 ( .A1(n5358), .A2(n17048), .B1(n3144), .B2(n17052), .ZN(
        U324_Z_0) );
  OAI22_X1 U2985 ( .A1(n5387), .A2(n17053), .B1(n3144), .B2(n17057), .ZN(
        U323_Z_0) );
  OAI22_X1 U2986 ( .A1(n5416), .A2(n17058), .B1(n3144), .B2(n17062), .ZN(
        U322_Z_0) );
  OAI22_X1 U2987 ( .A1(n5445), .A2(n17063), .B1(n3144), .B2(n17067), .ZN(
        U321_Z_0) );
  OAI22_X1 U2988 ( .A1(n5474), .A2(n17068), .B1(n3144), .B2(n17072), .ZN(
        U320_Z_0) );
  OAI22_X1 U2989 ( .A1(n5144), .A2(n17073), .B1(n3144), .B2(n17077), .ZN(
        U319_Z_0) );
  OAI22_X1 U2990 ( .A1(n5498), .A2(n17078), .B1(n3144), .B2(n17082), .ZN(
        U318_Z_0) );
  AOI221_X1 U2992 ( .B1(n2495), .B2(n16723), .C1(n3145), .C2(n17007), .A(n3146), .ZN(n2114) );
  INV_X1 U2993 ( .A(n3147), .ZN(n3146) );
  AOI211_X1 U2994 ( .C1(n5804), .C2(n3148), .A(n2055), .B(n3149), .ZN(n3147)
         );
  NOR3_X1 U2995 ( .A1(n5804), .A2(n16992), .A3(n1696), .ZN(n3149) );
  OAI22_X1 U2996 ( .A1(n2131), .A2(n1696), .B1(n2501), .B2(n1667), .ZN(n3148)
         );
  INV_X1 U2997 ( .A(n1667), .ZN(n1696) );
  NAND4_X1 U2998 ( .A1(n3150), .A2(n3151), .A3(n3152), .A4(n3153), .ZN(n1667)
         );
  AOI222_X1 U2999 ( .A1(n16974), .A2(vis_msp_o[8]), .B1(n16970), .B2(n3155), 
        .C1(n16969), .C2(vis_psp_o[8]), .ZN(n3153) );
  AOI222_X1 U3001 ( .A1(n16983), .A2(vis_r14_o[10]), .B1(n16966), .B2(
        vis_r12_o[10]), .C1(n16987), .C2(vis_r11_o[10]), .ZN(n3152) );
  AOI222_X1 U3004 ( .A1(n16980), .A2(vis_r9_o[10]), .B1(n16963), .B2(
        vis_r10_o[10]), .C1(n16960), .C2(vis_r8_o[10]), .ZN(n3151) );
  AOI22_X1 U3006 ( .A1(n16978), .A2(n3142), .B1(n16956), .B2(n869), .ZN(n3150)
         );
  XOR2_X1 U3008 ( .A(n2169), .B(n3163), .Z(n5804) );
  AOI222_X1 U3009 ( .A1(n16988), .A2(n3145), .B1(n2198), .B2(n16657), .C1(
        n3164), .C2(n2731), .ZN(n3163) );
  AOI221_X1 U3010 ( .B1(n2464), .B2(n2954), .C1(n2465), .C2(n2871), .A(n3165), 
        .ZN(n140) );
  INV_X1 U3011 ( .A(n3166), .ZN(n3165) );
  AOI221_X1 U3012 ( .B1(n2468), .B2(n2977), .C1(n2469), .C2(n2872), .A(n2873), 
        .ZN(n3166) );
  OAI22_X1 U3013 ( .A1(n5546), .A2(n3167), .B1(n3168), .B2(n3169), .ZN(
        U317_Z_0) );
  AOI22_X1 U3014 ( .A1(n1040), .A2(n1640), .B1(n3170), .B2(n1058), .ZN(n3168)
         );
  INV_X1 U3015 ( .A(n3169), .ZN(n3167) );
  OAI211_X1 U3016 ( .C1(n1173), .C2(n1880), .A(n17123), .B(n195), .ZN(n3169)
         );
  INV_X1 U3017 ( .A(n890), .ZN(n1880) );
  OAI22_X1 U3018 ( .A1(n5060), .A2(n17001), .B1(n3171), .B2(n17005), .ZN(
        U315_Z_0) );
  OAI22_X1 U3019 ( .A1(n5059), .A2(n16996), .B1(n3171), .B2(n17000), .ZN(
        U314_Z_0) );
  OAI22_X1 U3020 ( .A1(n5303), .A2(n17038), .B1(n3171), .B2(n17042), .ZN(
        U313_Z_0) );
  OAI22_X1 U3021 ( .A1(n5282), .A2(n17033), .B1(n3171), .B2(n17037), .ZN(
        U312_Z_0) );
  OAI22_X1 U3022 ( .A1(n5058), .A2(n17028), .B1(n3171), .B2(n17032), .ZN(
        U311_Z_0) );
  OAI22_X1 U3023 ( .A1(n5194), .A2(n17023), .B1(n3171), .B2(n17027), .ZN(
        U310_Z_0) );
  OAI22_X1 U3024 ( .A1(n5057), .A2(n17018), .B1(n3171), .B2(n17022), .ZN(
        U309_Z_0) );
  OAI22_X1 U3025 ( .A1(n5223), .A2(n17013), .B1(n3171), .B2(n17017), .ZN(
        U308_Z_0) );
  OAI22_X1 U3026 ( .A1(n5330), .A2(n17043), .B1(n3171), .B2(n17047), .ZN(
        U307_Z_0) );
  OAI22_X1 U3027 ( .A1(n5359), .A2(n17048), .B1(n3171), .B2(n17052), .ZN(
        U306_Z_0) );
  OAI22_X1 U3028 ( .A1(n5388), .A2(n17053), .B1(n3171), .B2(n17057), .ZN(
        U305_Z_0) );
  OAI22_X1 U3029 ( .A1(n5417), .A2(n17058), .B1(n3171), .B2(n17062), .ZN(
        U304_Z_0) );
  OAI22_X1 U3030 ( .A1(n5446), .A2(n17063), .B1(n3171), .B2(n17067), .ZN(
        U303_Z_0) );
  OAI22_X1 U3031 ( .A1(n5475), .A2(n17068), .B1(n3171), .B2(n17072), .ZN(
        U302_Z_0) );
  OAI22_X1 U3032 ( .A1(n5056), .A2(n17073), .B1(n3171), .B2(n17077), .ZN(
        U301_Z_0) );
  OAI22_X1 U3033 ( .A1(n5499), .A2(n17078), .B1(n3171), .B2(n17082), .ZN(
        U300_Z_0) );
  AND4_X1 U3035 ( .A1(n3172), .A2(n3173), .A3(n3174), .A4(n3175), .ZN(n2115)
         );
  AOI222_X1 U3036 ( .A1(n16729), .A2(n17009), .B1(n2055), .B2(vis_control_o), 
        .C1(n17007), .C2(n3177), .ZN(n3175) );
  AOI22_X1 U3038 ( .A1(n5806), .A2(n3178), .B1(n2227), .B2(vis_ipsr_o[2]), 
        .ZN(n3174) );
  NOR3_X1 U3039 ( .A1(n16671), .A2(n5120), .A3(n2168), .ZN(n2227) );
  OAI22_X1 U3040 ( .A1(n2131), .A2(n1676), .B1(n2501), .B2(n1640), .ZN(n3178)
         );
  OR4_X1 U3041 ( .A1(n1308), .A2(n5546), .A3(n16853), .A4(n4950), .ZN(n3173)
         );
  NAND2_X1 U3042 ( .A1(n17096), .A2(n16728), .ZN(n1308) );
  OR3_X1 U3043 ( .A1(n1676), .A2(n16992), .A3(n5806), .ZN(n3172) );
  XNOR2_X1 U3044 ( .A(n16990), .B(n3179), .ZN(n5806) );
  OAI221_X1 U3045 ( .B1(n5120), .B2(n2554), .C1(n3180), .C2(n3181), .A(n3182), 
        .ZN(n3179) );
  AOI22_X1 U3046 ( .A1(n461), .A2(n2198), .B1(n16656), .B2(n2173), .ZN(n3182)
         );
  NAND2_X1 U3047 ( .A1(n2201), .A2(n3183), .ZN(n2173) );
  NAND4_X1 U3048 ( .A1(n1097), .A2(n2661), .A3(n16841), .A4(n1697), .ZN(n3183)
         );
  INV_X1 U3049 ( .A(n3184), .ZN(n2201) );
  OAI21_X1 U3050 ( .B1(n4950), .B2(n3185), .A(n3186), .ZN(n3184) );
  AOI221_X1 U3051 ( .B1(n16862), .B2(n3187), .C1(n3188), .C2(n16871), .A(n3189), .ZN(n3185) );
  OAI22_X1 U3052 ( .A1(n1104), .A2(n1517), .B1(n919), .B2(n655), .ZN(n3189) );
  NAND2_X1 U3053 ( .A1(n17097), .A2(n16838), .ZN(n655) );
  OAI21_X1 U3054 ( .B1(n16837), .B2(n1211), .A(n919), .ZN(n3188) );
  NAND2_X1 U3055 ( .A1(n16830), .A2(n16856), .ZN(n919) );
  OAI22_X1 U3056 ( .A1(n16851), .A2(n1104), .B1(n16805), .B2(n648), .ZN(n3187)
         );
  INV_X1 U3057 ( .A(n3177), .ZN(n3181) );
  INV_X1 U3058 ( .A(n2577), .ZN(n2554) );
  OAI21_X1 U3059 ( .B1(n4950), .B2(n3190), .A(n2200), .ZN(n2577) );
  AOI221_X1 U3060 ( .B1(n3191), .B2(n16868), .C1(n507), .C2(n16839), .A(n3192), 
        .ZN(n3190) );
  OAI22_X1 U3061 ( .A1(n16806), .A2(n673), .B1(n585), .B2(n1211), .ZN(n3192)
         );
  NAND2_X1 U3062 ( .A1(n499), .A2(n994), .ZN(n507) );
  AOI21_X1 U3063 ( .B1(n1603), .B2(n3193), .A(n16866), .ZN(n3191) );
  NAND2_X1 U3064 ( .A1(n1564), .A2(n16858), .ZN(n3193) );
  INV_X1 U3065 ( .A(n1640), .ZN(n1676) );
  NAND4_X1 U3066 ( .A1(n3194), .A2(n3195), .A3(n3196), .A4(n3197), .ZN(n1640)
         );
  AOI222_X1 U3067 ( .A1(n16975), .A2(vis_msp_o[0]), .B1(n16970), .B2(n3199), 
        .C1(n16969), .C2(vis_psp_o[0]), .ZN(n3197) );
  AOI222_X1 U3068 ( .A1(n16984), .A2(vis_r14_o[2]), .B1(n16966), .B2(
        vis_r12_o[2]), .C1(n16987), .C2(vis_r11_o[2]), .ZN(n3196) );
  AOI222_X1 U3069 ( .A1(n16981), .A2(vis_r9_o[2]), .B1(n16963), .B2(
        vis_r10_o[2]), .C1(n16960), .C2(vis_r8_o[2]), .ZN(n3195) );
  AOI22_X1 U3070 ( .A1(n16978), .A2(n2620), .B1(n16955), .B2(n2635), .ZN(n3194) );
  AOI221_X1 U3072 ( .B1(n2008), .B2(n2468), .C1(n2002), .C2(n2465), .A(n3207), 
        .ZN(n171) );
  INV_X1 U3073 ( .A(n3208), .ZN(n3207) );
  AOI221_X1 U3074 ( .B1(n2469), .B2(n2011), .C1(n2464), .C2(n2004), .A(n2012), 
        .ZN(n3208) );
  AND4_X1 U3075 ( .A1(n3209), .A2(n3210), .A3(n3211), .A4(n3212), .ZN(n2012)
         );
  AOI222_X1 U3076 ( .A1(n2360), .A2(n3213), .B1(n3214), .B2(n2341), .C1(n3215), 
        .C2(n3216), .ZN(n3212) );
  INV_X1 U3077 ( .A(n3217), .ZN(n2360) );
  AOI211_X1 U3079 ( .C1(n3219), .C2(n606), .A(n1712), .B(n3220), .ZN(n3218) );
  AOI211_X1 U3080 ( .C1(n16841), .C2(n3221), .A(n3222), .B(n3223), .ZN(n3220)
         );
  NAND2_X1 U3081 ( .A1(n16838), .A2(n16856), .ZN(n3219) );
  NAND3_X1 U3082 ( .A1(n3224), .A2(n3225), .A3(n3226), .ZN(n2464) );
  AOI221_X1 U3083 ( .B1(n16787), .B2(n3227), .C1(sub_2068_A_2_), .C2(n2878), 
        .A(n3228), .ZN(n3226) );
  OAI22_X1 U3084 ( .A1(n2918), .A2(n425), .B1(n4801), .B2(n2948), .ZN(n3228)
         );
  INV_X1 U3085 ( .A(hrdata_i[2]), .ZN(n425) );
  AOI221_X1 U3087 ( .B1(n2912), .B2(n2325), .C1(n3058), .C2(n3229), .A(n3230), 
        .ZN(n3225) );
  OAI221_X1 U3089 ( .B1(n3231), .B2(n16949), .C1(n3233), .C2(n16951), .A(n3234), .ZN(n2325) );
  AOI22_X1 U3090 ( .A1(n16946), .A2(n2209), .B1(n16944), .B2(n3237), .ZN(n3234) );
  AOI22_X1 U3091 ( .A1(n16645), .A2(n2332), .B1(n2913), .B2(n3238), .ZN(n3224)
         );
  OAI221_X1 U3092 ( .B1(n3239), .B2(n16948), .C1(n3240), .C2(n16951), .A(n3241), .ZN(n2332) );
  AOI22_X1 U3093 ( .A1(n16945), .A2(n2612), .B1(n16944), .B2(n2562), .ZN(n3241) );
  NAND3_X1 U3095 ( .A1(n5227), .A2(n3223), .A3(n3246), .ZN(n3244) );
  NAND4_X1 U3096 ( .A1(n3247), .A2(n3003), .A3(n3248), .A4(n3249), .ZN(n2469)
         );
  AOI222_X1 U3097 ( .A1(sub_2068_A_18_), .A2(n2878), .B1(hrdata_i[18]), .B2(
        n2879), .C1(n16787), .C2(n3250), .ZN(n3249) );
  AOI22_X1 U3099 ( .A1(n16645), .A2(n2352), .B1(n2912), .B2(n2344), .ZN(n3248)
         );
  OAI221_X1 U3100 ( .B1(n3251), .B2(n16948), .C1(n3252), .C2(n16951), .A(n3253), .ZN(n2344) );
  AOI22_X1 U3101 ( .A1(n16945), .A2(n3254), .B1(n16944), .B2(n2484), .ZN(n3253) );
  OAI221_X1 U3102 ( .B1(n3255), .B2(n16948), .C1(n3256), .C2(n16951), .A(n3257), .ZN(n2352) );
  AOI22_X1 U3103 ( .A1(n16945), .A2(n2787), .B1(n16944), .B2(n2738), .ZN(n3257) );
  NAND2_X1 U3104 ( .A1(n3258), .A2(n3259), .ZN(n2465) );
  AOI221_X1 U3105 ( .B1(n2912), .B2(n2388), .C1(n16645), .C2(n2329), .A(n3260), 
        .ZN(n3259) );
  OAI22_X1 U3106 ( .A1(n5537), .A2(n2948), .B1(n4748), .B2(n3011), .ZN(n3260)
         );
  OAI221_X1 U3107 ( .B1(n3261), .B2(n16948), .C1(n3262), .C2(n16951), .A(n3263), .ZN(n2329) );
  AOI22_X1 U3108 ( .A1(n16945), .A2(n3134), .B1(n16944), .B2(n3022), .ZN(n3263) );
  OAI221_X1 U3109 ( .B1(n3264), .B2(n16948), .C1(n3265), .C2(n16951), .A(n3266), .ZN(n2388) );
  AOI22_X1 U3110 ( .A1(n16945), .A2(n3267), .B1(n16944), .B2(n2833), .ZN(n3266) );
  AOI222_X1 U3111 ( .A1(sub_2068_A_10_), .A2(n2878), .B1(hrdata_i[10]), .B2(
        n2879), .C1(n16787), .C2(n3268), .ZN(n3258) );
  NAND3_X1 U3113 ( .A1(n3269), .A2(n3210), .A3(n3270), .ZN(n2002) );
  AOI22_X1 U3114 ( .A1(n3271), .A2(n3246), .B1(n1207), .B2(n3215), .ZN(n3270)
         );
  NOR2_X1 U3115 ( .A1(n5227), .A2(n3223), .ZN(n3271) );
  OAI211_X1 U3116 ( .C1(n3001), .C2(n2371), .A(n3272), .B(n3273), .ZN(n2468)
         );
  AOI22_X1 U3117 ( .A1(n2895), .A2(n203), .B1(hrdata_i[26]), .B2(n2879), .ZN(
        n3273) );
  NAND3_X1 U3118 ( .A1(n2370), .A2(n2371), .A3(n2922), .ZN(n3272) );
  OAI22_X1 U3119 ( .A1(n2874), .A2(n16789), .B1(n2937), .B2(n2337), .ZN(n2370)
         );
  AOI221_X1 U3120 ( .B1(n3274), .B2(n3275), .C1(n2297), .C2(n3118), .A(n3276), 
        .ZN(n2937) );
  OAI22_X1 U3121 ( .A1(n3277), .A2(n3278), .B1(n3279), .B2(n3280), .ZN(n3276)
         );
  INV_X1 U3122 ( .A(n2349), .ZN(n2874) );
  OAI221_X1 U3123 ( .B1(n3281), .B2(n16948), .C1(n3282), .C2(n16951), .A(n3283), .ZN(n2349) );
  AOI22_X1 U3124 ( .A1(n16945), .A2(n2433), .B1(n16944), .B2(n2402), .ZN(n3283) );
  OAI221_X1 U3125 ( .B1(n2939), .B2(n3119), .C1(n3120), .C2(n2942), .A(n3122), 
        .ZN(n2371) );
  INV_X1 U3126 ( .A(n2942), .ZN(n2939) );
  NAND3_X1 U3128 ( .A1(n3222), .A2(n3223), .A3(n3246), .ZN(n3284) );
  NOR3_X1 U3129 ( .A1(n17096), .A2(n16841), .A3(n3213), .ZN(n3246) );
  OAI22_X1 U3131 ( .A1(n5577), .A2(n17001), .B1(n3286), .B2(n17005), .ZN(
        U299_Z_0) );
  OAI22_X1 U3132 ( .A1(n5576), .A2(n16996), .B1(n3286), .B2(n17000), .ZN(
        U298_Z_0) );
  OAI22_X1 U3133 ( .A1(n5575), .A2(n17038), .B1(n3286), .B2(n17042), .ZN(
        U297_Z_0) );
  OAI22_X1 U3134 ( .A1(n5574), .A2(n17033), .B1(n3286), .B2(n17037), .ZN(
        U296_Z_0) );
  OAI22_X1 U3135 ( .A1(n5143), .A2(n17028), .B1(n3286), .B2(n17032), .ZN(
        U295_Z_0) );
  OAI22_X1 U3136 ( .A1(n5195), .A2(n17023), .B1(n3286), .B2(n17027), .ZN(
        U294_Z_0) );
  OAI22_X1 U3137 ( .A1(n5142), .A2(n17018), .B1(n3286), .B2(n17022), .ZN(
        U293_Z_0) );
  OAI22_X1 U3138 ( .A1(n5224), .A2(n17013), .B1(n3286), .B2(n17017), .ZN(
        U292_Z_0) );
  OAI22_X1 U3139 ( .A1(n5331), .A2(n17043), .B1(n3286), .B2(n17047), .ZN(
        U291_Z_0) );
  OAI22_X1 U3140 ( .A1(n5360), .A2(n17048), .B1(n3286), .B2(n17052), .ZN(
        U290_Z_0) );
  OAI22_X1 U3142 ( .A1(n5389), .A2(n17053), .B1(n3286), .B2(n17057), .ZN(
        U289_Z_0) );
  OAI22_X1 U3143 ( .A1(n5418), .A2(n17058), .B1(n3286), .B2(n17062), .ZN(
        U288_Z_0) );
  OAI22_X1 U3144 ( .A1(n5447), .A2(n17063), .B1(n3286), .B2(n17067), .ZN(
        U287_Z_0) );
  OAI22_X1 U3145 ( .A1(n5476), .A2(n17068), .B1(n3286), .B2(n17072), .ZN(
        U286_Z_0) );
  OAI22_X1 U3146 ( .A1(n5141), .A2(n17073), .B1(n3286), .B2(n17077), .ZN(
        U285_Z_0) );
  OAI22_X1 U3147 ( .A1(n5541), .A2(n17078), .B1(n3286), .B2(n17082), .ZN(
        U284_Z_0) );
  AOI221_X1 U3149 ( .B1(n2495), .B2(n16727), .C1(n3287), .C2(n17007), .A(n3288), .ZN(n2113) );
  INV_X1 U3150 ( .A(n3289), .ZN(n3288) );
  AOI211_X1 U3151 ( .C1(n5805), .C2(n3290), .A(n2055), .B(n3291), .ZN(n3289)
         );
  NOR3_X1 U3152 ( .A1(n5805), .A2(n16992), .A3(n1621), .ZN(n3291) );
  OAI22_X1 U3153 ( .A1(n2131), .A2(n1621), .B1(n2501), .B2(n3292), .ZN(n3290)
         );
  INV_X1 U3154 ( .A(n3292), .ZN(n1621) );
  NAND4_X1 U3155 ( .A1(n3293), .A2(n3294), .A3(n3295), .A4(n3296), .ZN(n3292)
         );
  AOI222_X1 U3156 ( .A1(n16975), .A2(vis_msp_o[7]), .B1(n16970), .B2(n3237), 
        .C1(n16969), .C2(vis_psp_o[7]), .ZN(n3296) );
  AOI222_X1 U3158 ( .A1(n16984), .A2(vis_r14_o[9]), .B1(n16966), .B2(
        vis_r12_o[9]), .C1(n16987), .C2(vis_r11_o[9]), .ZN(n3295) );
  AOI222_X1 U3161 ( .A1(n16981), .A2(vis_r9_o[9]), .B1(n16963), .B2(
        vis_r10_o[9]), .C1(n16960), .C2(vis_r8_o[9]), .ZN(n3294) );
  AOI22_X1 U3163 ( .A1(n16978), .A2(n869), .B1(n16956), .B2(n1161), .ZN(n3293)
         );
  XOR2_X1 U3165 ( .A(n2169), .B(n3305), .Z(n5805) );
  AOI221_X1 U3166 ( .B1(n2198), .B2(n17098), .C1(n16988), .C2(n3287), .A(n3306), .ZN(n3305) );
  OAI22_X1 U3167 ( .A1(n5003), .A2(n3186), .B1(n5258), .B2(n2200), .ZN(n3306)
         );
  INV_X1 U3168 ( .A(n3170), .ZN(n127) );
  OAI221_X1 U3169 ( .B1(n3051), .B2(n2472), .C1(n2473), .C2(n2869), .A(n3307), 
        .ZN(n3170) );
  AOI221_X1 U3170 ( .B1(n2003), .B2(n2871), .C1(n2005), .C2(n2954), .A(n2873), 
        .ZN(n3307) );
  NAND3_X1 U3171 ( .A1(n3308), .A2(n3309), .A3(n3310), .ZN(n2005) );
  AOI221_X1 U3172 ( .B1(n16787), .B2(n3311), .C1(sub_2068_A_1_), .C2(n2878), 
        .A(n3312), .ZN(n3310) );
  OAI22_X1 U3173 ( .A1(n2918), .A2(n427), .B1(n5535), .B2(n2948), .ZN(n3312)
         );
  INV_X1 U3174 ( .A(hrdata_i[1]), .ZN(n427) );
  AOI222_X1 U3176 ( .A1(n16645), .A2(n2336), .B1(n3058), .B2(n3313), .C1(n2912), .C2(n2326), .ZN(n3309) );
  OAI221_X1 U3177 ( .B1(n3314), .B2(n16948), .C1(n3315), .C2(n16951), .A(n3316), .ZN(n2326) );
  AOI22_X1 U3178 ( .A1(n16945), .A2(n2531), .B1(n16943), .B2(n3317), .ZN(n3316) );
  AND2_X1 U3179 ( .A1(n3318), .A2(n1111), .ZN(n3058) );
  OAI221_X1 U3180 ( .B1(n3319), .B2(n16948), .C1(n3280), .C2(n16951), .A(n3320), .ZN(n2336) );
  AOI22_X1 U3181 ( .A1(n16945), .A2(n3199), .B1(n16943), .B2(n2585), .ZN(n3320) );
  INV_X1 U3182 ( .A(n3321), .ZN(n3308) );
  OAI22_X1 U3183 ( .A1(n3322), .A2(n4833), .B1(n3011), .B2(n5534), .ZN(n3321)
         );
  NAND3_X1 U3184 ( .A1(n3323), .A2(n3324), .A3(n3325), .ZN(n2003) );
  AOI221_X1 U3185 ( .B1(n16787), .B2(n3326), .C1(sub_2068_A_9_), .C2(n2878), 
        .A(n3327), .ZN(n3325) );
  OAI22_X1 U3186 ( .A1(n2918), .A2(n391), .B1(n5578), .B2(n2948), .ZN(n3327)
         );
  INV_X1 U3187 ( .A(hrdata_i[9]), .ZN(n391) );
  AOI211_X1 U3189 ( .C1(n16645), .C2(n2330), .A(n3106), .B(n2897), .ZN(n3324)
         );
  AND4_X1 U3190 ( .A1(n3318), .A2(n1189), .A3(n5096), .A4(n251), .ZN(n3106) );
  OAI221_X1 U3191 ( .B1(n3328), .B2(n16948), .C1(n3329), .C2(n16952), .A(n3330), .ZN(n2330) );
  AOI22_X1 U3192 ( .A1(n16945), .A2(n3155), .B1(n16943), .B2(n3041), .ZN(n3330) );
  INV_X1 U3193 ( .A(n3331), .ZN(n3323) );
  OAI22_X1 U3194 ( .A1(n2875), .A2(n2378), .B1(n3011), .B2(n5011), .ZN(n3331)
         );
  INV_X1 U3195 ( .A(n2988), .ZN(n2378) );
  OAI221_X1 U3196 ( .B1(n3332), .B2(n16948), .C1(n3333), .C2(n16952), .A(n3334), .ZN(n2988) );
  AOI22_X1 U3197 ( .A1(n16945), .A2(n2964), .B1(n16943), .B2(n2856), .ZN(n3334) );
  INV_X1 U3198 ( .A(n2977), .ZN(n2869) );
  INV_X1 U3199 ( .A(n2009), .ZN(n2473) );
  OAI211_X1 U3200 ( .C1(n3001), .C2(n3335), .A(n3003), .B(n3336), .ZN(n2009)
         );
  INV_X1 U3201 ( .A(n3337), .ZN(n3336) );
  OAI22_X1 U3202 ( .A1(n2372), .A2(n2998), .B1(n1140), .B2(n2918), .ZN(n3337)
         );
  INV_X1 U3203 ( .A(hrdata_i[25]), .ZN(n1140) );
  OAI221_X1 U3204 ( .B1(n2337), .B2(n3004), .C1(n16789), .C2(n2357), .A(n3335), 
        .ZN(n2372) );
  OAI221_X1 U3205 ( .B1(n3338), .B2(n16949), .C1(n3339), .C2(n16952), .A(n3340), .ZN(n2357) );
  AOI22_X1 U3206 ( .A1(n16946), .A2(n2452), .B1(n16943), .B2(n2271), .ZN(n3340) );
  OAI221_X1 U3207 ( .B1(n3278), .B2(n16949), .C1(n3341), .C2(n16952), .A(n3342), .ZN(n3004) );
  AOI22_X1 U3208 ( .A1(n16946), .A2(n2297), .B1(n16943), .B2(n3274), .ZN(n3342) );
  OAI221_X1 U3209 ( .B1(n3005), .B2(n3119), .C1(n3120), .C2(n3006), .A(n3122), 
        .ZN(n3335) );
  AOI21_X1 U3210 ( .B1(n3343), .B2(n2337), .A(n16851), .ZN(n3122) );
  INV_X1 U3211 ( .A(n3005), .ZN(n3006) );
  NAND2_X1 U3212 ( .A1(n2942), .A2(n16950), .ZN(n3005) );
  NOR2_X1 U3213 ( .A1(n3118), .A2(n16947), .ZN(n2942) );
  NAND2_X1 U3214 ( .A1(n2313), .A2(n2922), .ZN(n3001) );
  INV_X1 U3215 ( .A(n2010), .ZN(n2472) );
  OAI221_X1 U3216 ( .B1(n5639), .B2(n16685), .C1(n2981), .C2(n278), .A(n3344), 
        .ZN(n2010) );
  AOI222_X1 U3217 ( .A1(hrdata_i[17]), .A2(n2879), .B1(n16645), .B2(n2353), 
        .C1(n2912), .C2(n2345), .ZN(n3344) );
  OAI221_X1 U3218 ( .B1(n3345), .B2(n16949), .C1(n3346), .C2(n16952), .A(n3347), .ZN(n2345) );
  AOI22_X1 U3219 ( .A1(n16946), .A2(n2705), .B1(n16943), .B2(n2507), .ZN(n3347) );
  NAND2_X1 U3221 ( .A1(n2922), .A2(n16788), .ZN(n2875) );
  OAI221_X1 U3222 ( .B1(n3348), .B2(n16949), .C1(n3349), .C2(n16952), .A(n3350), .ZN(n2353) );
  AOI22_X1 U3223 ( .A1(n16946), .A2(n2809), .B1(n16943), .B2(n2764), .ZN(n3350) );
  INV_X1 U3226 ( .A(n2872), .ZN(n3051) );
  OAI22_X1 U3227 ( .A1(n5139), .A2(n17001), .B1(n3351), .B2(n17005), .ZN(
        U283_Z_0) );
  OAI22_X1 U3228 ( .A1(n5138), .A2(n16996), .B1(n3351), .B2(n17000), .ZN(
        U282_Z_0) );
  OAI22_X1 U3229 ( .A1(n5304), .A2(n17038), .B1(n3351), .B2(n17042), .ZN(
        U281_Z_0) );
  OAI22_X1 U3230 ( .A1(n5283), .A2(n17033), .B1(n3351), .B2(n17037), .ZN(
        U280_Z_0) );
  OAI22_X1 U3231 ( .A1(n5137), .A2(n17028), .B1(n3351), .B2(n17032), .ZN(
        U279_Z_0) );
  OAI22_X1 U3232 ( .A1(n5196), .A2(n17023), .B1(n3351), .B2(n17027), .ZN(
        U278_Z_0) );
  OAI22_X1 U3233 ( .A1(n5136), .A2(n17018), .B1(n3351), .B2(n17022), .ZN(
        U277_Z_0) );
  OAI22_X1 U3234 ( .A1(n5225), .A2(n17013), .B1(n3351), .B2(n17017), .ZN(
        U276_Z_0) );
  OAI22_X1 U3235 ( .A1(n5332), .A2(n17043), .B1(n3351), .B2(n17047), .ZN(
        U275_Z_0) );
  OAI22_X1 U3236 ( .A1(n5361), .A2(n17048), .B1(n3351), .B2(n17052), .ZN(
        U274_Z_0) );
  OAI22_X1 U3237 ( .A1(n5390), .A2(n17053), .B1(n3351), .B2(n17057), .ZN(
        U273_Z_0) );
  OAI22_X1 U3238 ( .A1(n5419), .A2(n17058), .B1(n3351), .B2(n17062), .ZN(
        U272_Z_0) );
  OAI22_X1 U3239 ( .A1(n5448), .A2(n17063), .B1(n3351), .B2(n17067), .ZN(
        U271_Z_0) );
  OAI22_X1 U3240 ( .A1(n5477), .A2(n17068), .B1(n3351), .B2(n17072), .ZN(
        U270_Z_0) );
  OAI22_X1 U3242 ( .A1(n5135), .A2(n17073), .B1(n3351), .B2(n17077), .ZN(
        U269_Z_0) );
  OAI22_X1 U3243 ( .A1(n5542), .A2(n17078), .B1(n3351), .B2(n17082), .ZN(
        U268_Z_0) );
  AOI221_X1 U3245 ( .B1(n17006), .B2(n2261), .C1(n16722), .C2(n17010), .A(
        n2055), .ZN(n3353) );
  OAI221_X1 U3246 ( .B1(n3354), .B2(n5819), .C1(n16995), .C2(n2148), .A(n3355), 
        .ZN(n3352) );
  NAND3_X1 U3247 ( .A1(n2131), .A2(n2148), .A3(n5819), .ZN(n3355) );
  AOI221_X1 U3249 ( .B1(n2198), .B2(n16798), .C1(n16988), .C2(n2261), .A(n3357), .ZN(n3356) );
  OAI22_X1 U3250 ( .A1(n5162), .A2(n3186), .B1(n5257), .B2(n2200), .ZN(n3357)
         );
  OAI21_X1 U3251 ( .B1(n3358), .B2(n3359), .A(n1697), .ZN(n2200) );
  OAI22_X1 U3252 ( .A1(n3360), .A2(n745), .B1(n758), .B2(n3361), .ZN(n3359) );
  NAND2_X1 U3253 ( .A1(n16851), .A2(n991), .ZN(n3361) );
  NOR3_X1 U3254 ( .A1(n16847), .A2(n760), .A3(n798), .ZN(n3360) );
  INV_X1 U3255 ( .A(n3362), .ZN(n798) );
  OAI33_X1 U3256 ( .A1(n3363), .A2(n1086), .A3(n653), .B1(n863), .B2(n16851), 
        .B3(n3362), .ZN(n3358) );
  NAND2_X1 U3257 ( .A1(n991), .A2(n16860), .ZN(n863) );
  NOR2_X1 U3258 ( .A1(n1625), .A2(n16993), .ZN(n3354) );
  INV_X1 U3259 ( .A(n2148), .ZN(n1625) );
  NAND4_X1 U3260 ( .A1(n3364), .A2(n3365), .A3(n3366), .A4(n3367), .ZN(n2148)
         );
  AOI222_X1 U3261 ( .A1(n16975), .A2(vis_msp_o[6]), .B1(n16970), .B2(n3317), 
        .C1(n16969), .C2(vis_psp_o[6]), .ZN(n3367) );
  AOI222_X1 U3263 ( .A1(n16983), .A2(vis_r14_o[8]), .B1(n16966), .B2(
        vis_r12_o[8]), .C1(n16987), .C2(vis_r11_o[8]), .ZN(n3366) );
  AOI222_X1 U3266 ( .A1(n16981), .A2(vis_r9_o[8]), .B1(n16963), .B2(
        vis_r10_o[8]), .C1(n16960), .C2(vis_r8_o[8]), .ZN(n3365) );
  AOI22_X1 U3268 ( .A1(n16978), .A2(n1161), .B1(n16956), .B2(n2221), .ZN(n3364) );
  AOI221_X1 U3270 ( .B1(n2022), .B2(n2977), .C1(n2018), .C2(n2954), .A(n3376), 
        .ZN(n144) );
  INV_X1 U3271 ( .A(n3377), .ZN(n3376) );
  AOI221_X1 U3272 ( .B1(n2871), .B2(n2019), .C1(n2023), .C2(n2872), .A(n2873), 
        .ZN(n3377) );
  NAND4_X1 U3273 ( .A1(n3378), .A2(n3003), .A3(n3379), .A4(n3380), .ZN(n2023)
         );
  AOI222_X1 U3274 ( .A1(sub_2068_A_16_), .A2(n2878), .B1(hrdata_i[16]), .B2(
        n2879), .C1(n16787), .C2(n3381), .ZN(n3380) );
  INV_X1 U3276 ( .A(n3382), .ZN(n3379) );
  OAI22_X1 U3277 ( .A1(n1779), .A2(n2998), .B1(n3322), .B2(n5068), .ZN(n3382)
         );
  OAI22_X1 U3278 ( .A1(n2337), .A2(n2355), .B1(n16789), .B2(n2385), .ZN(n1779)
         );
  OAI221_X1 U3279 ( .B1(n3256), .B2(n16949), .C1(n3264), .C2(n16952), .A(n3383), .ZN(n2385) );
  AOI22_X1 U3280 ( .A1(n16946), .A2(n2833), .B1(n16943), .B2(n2787), .ZN(n3383) );
  OAI221_X1 U3281 ( .B1(n3252), .B2(n16949), .C1(n3255), .C2(n16952), .A(n3384), .ZN(n2355) );
  AOI22_X1 U3282 ( .A1(n16946), .A2(n2738), .B1(n16943), .B2(n3254), .ZN(n3384) );
  NAND2_X1 U3283 ( .A1(n405), .A2(n2895), .ZN(n3378) );
  INV_X1 U3284 ( .A(n421), .ZN(n405) );
  NAND3_X1 U3285 ( .A1(n2907), .A2(n1372), .A3(n2905), .ZN(n421) );
  INV_X1 U3286 ( .A(n3385), .ZN(n2019) );
  AOI211_X1 U3287 ( .C1(n2878), .C2(sub_2068_A_8_), .A(n3386), .B(n3387), .ZN(
        n3385) );
  OAI222_X1 U3288 ( .A1(n3011), .A2(n4747), .B1(n2948), .B2(n4796), .C1(n393), 
        .C2(n2918), .ZN(n3387) );
  INV_X1 U3289 ( .A(hrdata_i[8]), .ZN(n393) );
  OAI22_X1 U3290 ( .A1(n1772), .A2(n2998), .B1(n16685), .B2(n5581), .ZN(n3386)
         );
  OAI22_X1 U3291 ( .A1(n2337), .A2(n2387), .B1(n16789), .B2(n2339), .ZN(n1772)
         );
  OAI221_X1 U3292 ( .B1(n3262), .B2(n16949), .C1(n3231), .C2(n16952), .A(n3388), .ZN(n2339) );
  AOI22_X1 U3293 ( .A1(n16946), .A2(n3237), .B1(n16943), .B2(n3134), .ZN(n3388) );
  OAI221_X1 U3294 ( .B1(n3265), .B2(n16949), .C1(n3261), .C2(n16952), .A(n3389), .ZN(n2387) );
  AOI22_X1 U3295 ( .A1(n16946), .A2(n3022), .B1(n16942), .B2(n3267), .ZN(n3389) );
  INV_X1 U3297 ( .A(n2517), .ZN(n2018) );
  NOR2_X1 U3298 ( .A1(n3390), .A2(n3391), .ZN(n2517) );
  OAI221_X1 U3299 ( .B1(n3322), .B2(n5516), .C1(n1781), .C2(n2998), .A(n3392), 
        .ZN(n3391) );
  INV_X1 U3300 ( .A(n3393), .ZN(n3392) );
  OAI22_X1 U3301 ( .A1(n5540), .A2(n2948), .B1(n5005), .B2(n3011), .ZN(n3393)
         );
  OAI22_X1 U3302 ( .A1(n2337), .A2(n2333), .B1(n16789), .B2(n3094), .ZN(n1781)
         );
  OAI221_X1 U3303 ( .B1(n3240), .B2(n16949), .C1(n2183), .C2(n16953), .A(n3394), .ZN(n3094) );
  AOI22_X1 U3304 ( .A1(n16946), .A2(n2639), .B1(n16942), .B2(n2612), .ZN(n3394) );
  OAI221_X1 U3305 ( .B1(n3314), .B2(n3279), .C1(n3239), .C2(n16953), .A(n3395), 
        .ZN(n2333) );
  AOI22_X1 U3306 ( .A1(n16946), .A2(n2562), .B1(n3275), .B2(n2531), .ZN(n3395)
         );
  INV_X1 U3307 ( .A(n3230), .ZN(n3322) );
  NOR3_X1 U3308 ( .A1(n251), .A2(n2926), .A3(n261), .ZN(n3230) );
  OAI222_X1 U3309 ( .A1(n260), .A2(n2981), .B1(n429), .B2(n2918), .C1(n16685), 
        .C2(n5510), .ZN(n3390) );
  INV_X1 U3310 ( .A(hrdata_i[0]), .ZN(n429) );
  INV_X1 U3311 ( .A(n2516), .ZN(n2022) );
  AOI221_X1 U3312 ( .B1(n2879), .B2(hrdata_i[24]), .C1(n2363), .C2(n2922), .A(
        n2897), .ZN(n2516) );
  OAI22_X1 U3313 ( .A1(n1782), .A2(n3396), .B1(n3092), .B2(n3397), .ZN(n2363)
         );
  INV_X1 U3314 ( .A(n3397), .ZN(n3396) );
  NAND2_X1 U3315 ( .A1(n3120), .A2(n16849), .ZN(n3397) );
  AOI22_X1 U3316 ( .A1(n2350), .A2(n2337), .B1(n3095), .B2(n16788), .ZN(n1782)
         );
  OAI221_X1 U3317 ( .B1(n3398), .B2(n16949), .C1(n3281), .C2(n16953), .A(n3399), .ZN(n3095) );
  AOI22_X1 U3318 ( .A1(n16947), .A2(n2402), .B1(n16942), .B2(n3400), .ZN(n3399) );
  OAI221_X1 U3319 ( .B1(n3282), .B2(n16950), .C1(n3251), .C2(n16953), .A(n3401), .ZN(n2350) );
  AOI22_X1 U3320 ( .A1(n16947), .A2(n2484), .B1(n16942), .B2(n2433), .ZN(n3401) );
  OAI22_X1 U3321 ( .A1(n5634), .A2(n17001), .B1(n3402), .B2(n17005), .ZN(
        U265_Z_0) );
  OAI22_X1 U3322 ( .A1(n5633), .A2(n16996), .B1(n3402), .B2(n17000), .ZN(
        U264_Z_0) );
  OAI22_X1 U3323 ( .A1(n5632), .A2(n17038), .B1(n3402), .B2(n17042), .ZN(
        U263_Z_0) );
  OAI22_X1 U3324 ( .A1(n5631), .A2(n17033), .B1(n3402), .B2(n17037), .ZN(
        U262_Z_0) );
  OAI22_X1 U3325 ( .A1(n5110), .A2(n17028), .B1(n3402), .B2(n17032), .ZN(
        U261_Z_0) );
  OAI22_X1 U3326 ( .A1(n5197), .A2(n17023), .B1(n3402), .B2(n17027), .ZN(
        U260_Z_0) );
  OAI22_X1 U3328 ( .A1(n5109), .A2(n17018), .B1(n3402), .B2(n17022), .ZN(
        U259_Z_0) );
  OAI22_X1 U3329 ( .A1(n5226), .A2(n17013), .B1(n3402), .B2(n17017), .ZN(
        U258_Z_0) );
  OAI22_X1 U3330 ( .A1(n5333), .A2(n17043), .B1(n3402), .B2(n17047), .ZN(
        U257_Z_0) );
  OAI22_X1 U3331 ( .A1(n5362), .A2(n17048), .B1(n3402), .B2(n17052), .ZN(
        U256_Z_0) );
  OAI22_X1 U3332 ( .A1(n5391), .A2(n17053), .B1(n3402), .B2(n17057), .ZN(
        U255_Z_0) );
  OAI22_X1 U3333 ( .A1(n5420), .A2(n17058), .B1(n3402), .B2(n17062), .ZN(
        U254_Z_0) );
  OAI22_X1 U3334 ( .A1(n5449), .A2(n17063), .B1(n3402), .B2(n17067), .ZN(
        U253_Z_0) );
  OAI22_X1 U3335 ( .A1(n5478), .A2(n17068), .B1(n3402), .B2(n17072), .ZN(
        U252_Z_0) );
  OAI22_X1 U3336 ( .A1(n5108), .A2(n17073), .B1(n3402), .B2(n17077), .ZN(
        U251_Z_0) );
  OAI22_X1 U3337 ( .A1(n5543), .A2(n17078), .B1(n3402), .B2(n17082), .ZN(
        U250_Z_0) );
  AOI221_X1 U3339 ( .B1(n17006), .B2(n2254), .C1(n16715), .C2(n17010), .A(
        n2055), .ZN(n3404) );
  OAI221_X1 U3340 ( .B1(n3405), .B2(n5818), .C1(n16995), .C2(n2144), .A(n3406), 
        .ZN(n3403) );
  NAND3_X1 U3341 ( .A1(n2131), .A2(n2144), .A3(n5818), .ZN(n3406) );
  AOI221_X1 U3343 ( .B1(n16989), .B2(n2254), .C1(n2198), .C2(n16671), .A(n2732), .ZN(n3407) );
  NOR2_X1 U3344 ( .A1(n1661), .A2(n16993), .ZN(n3405) );
  INV_X1 U3345 ( .A(n2144), .ZN(n1661) );
  NAND4_X1 U3346 ( .A1(n3408), .A2(n3409), .A3(n3410), .A4(n3411), .ZN(n2144)
         );
  AOI222_X1 U3347 ( .A1(n16975), .A2(vis_msp_o[13]), .B1(n16970), .B2(n3267), 
        .C1(n16969), .C2(vis_psp_o[13]), .ZN(n3411) );
  AOI222_X1 U3349 ( .A1(n16984), .A2(vis_r14_o[15]), .B1(n16966), .B2(
        vis_r12_o[15]), .C1(n16987), .C2(vis_r11_o[15]), .ZN(n3410) );
  AOI222_X1 U3352 ( .A1(n16981), .A2(vis_r9_o[15]), .B1(n16963), .B2(
        vis_r10_o[15]), .C1(n16960), .C2(vis_r8_o[15]), .ZN(n3409) );
  AOI22_X1 U3354 ( .A1(n16978), .A2(n1163), .B1(n16956), .B2(n2961), .ZN(n3408) );
  AOI221_X1 U3357 ( .B1(n2872), .B2(n2061), .C1(n2977), .C2(n2057), .A(n3420), 
        .ZN(n48) );
  INV_X1 U3358 ( .A(n3421), .ZN(n3420) );
  AOI221_X1 U3359 ( .B1(n2954), .B2(n2062), .C1(n2871), .C2(n2058), .A(n2873), 
        .ZN(n3421) );
  INV_X1 U3360 ( .A(n3422), .ZN(n2873) );
  OAI211_X1 U3361 ( .C1(n2377), .C2(n3215), .A(n3423), .B(n3424), .ZN(n3422)
         );
  NOR2_X1 U3362 ( .A1(n3214), .A2(n3425), .ZN(n3424) );
  NAND4_X1 U3363 ( .A1(n3215), .A2(n1518), .A3(n3216), .A4(n3426), .ZN(n3423)
         );
  NAND3_X1 U3364 ( .A1(n16837), .A2(n16871), .A3(n195), .ZN(n3426) );
  AOI211_X1 U3365 ( .C1(n2341), .C2(n2358), .A(n2321), .B(n2322), .ZN(n2377)
         );
  INV_X1 U3367 ( .A(n2720), .ZN(n2756) );
  AOI211_X1 U3368 ( .C1(n5102), .C2(n3428), .A(n1712), .B(n728), .ZN(n3427) );
  INV_X1 U3369 ( .A(n605), .ZN(n728) );
  NOR2_X1 U3370 ( .A1(n1210), .A2(n16851), .ZN(n1712) );
  NAND2_X1 U3371 ( .A1(n16842), .A2(n16860), .ZN(n1210) );
  OAI21_X1 U3372 ( .B1(n16839), .B2(n1580), .A(n3429), .ZN(n3428) );
  NAND2_X1 U3373 ( .A1(n2417), .A2(n3269), .ZN(n2954) );
  NAND3_X1 U3374 ( .A1(n827), .A2(n3430), .A3(n3215), .ZN(n3269) );
  INV_X1 U3375 ( .A(n2067), .ZN(n2417) );
  NAND3_X1 U3376 ( .A1(n3243), .A2(n3245), .A3(n3431), .ZN(n2977) );
  NAND3_X1 U3377 ( .A1(n3215), .A2(n3223), .A3(n3432), .ZN(n3431) );
  NAND4_X1 U3378 ( .A1(n3215), .A2(n990), .A3(n3223), .A4(n16841), .ZN(n3245)
         );
  INV_X1 U3379 ( .A(n1964), .ZN(n990) );
  NAND2_X1 U3380 ( .A1(n3285), .A2(n3210), .ZN(n2872) );
  NAND2_X1 U3381 ( .A1(n3433), .A2(n2341), .ZN(n3210) );
  OAI22_X1 U3382 ( .A1(n5595), .A2(n17001), .B1(n3434), .B2(n17004), .ZN(
        U247_Z_0) );
  OAI22_X1 U3385 ( .A1(n4970), .A2(n16996), .B1(n3434), .B2(n16999), .ZN(
        U246_Z_0) );
  OAI22_X1 U3388 ( .A1(n5594), .A2(n17038), .B1(n3434), .B2(n17041), .ZN(
        U245_Z_0) );
  OAI22_X1 U3391 ( .A1(n5593), .A2(n17033), .B1(n3434), .B2(n17036), .ZN(
        U244_Z_0) );
  AND2_X1 U3394 ( .A1(n3440), .A2(n3441), .ZN(n3437) );
  OAI22_X1 U3395 ( .A1(n4960), .A2(n17028), .B1(n3434), .B2(n17031), .ZN(
        U243_Z_0) );
  OAI22_X1 U3398 ( .A1(n5592), .A2(n17023), .B1(n3434), .B2(n17026), .ZN(
        U242_Z_0) );
  OAI22_X1 U3401 ( .A1(n5591), .A2(n17018), .B1(n3434), .B2(n17021), .ZN(
        U241_Z_0) );
  OAI22_X1 U3404 ( .A1(n5590), .A2(n17013), .B1(n3434), .B2(n17016), .ZN(
        U240_Z_0) );
  AND2_X1 U3407 ( .A1(n3444), .A2(n3441), .ZN(n3442) );
  OAI22_X1 U3408 ( .A1(n5589), .A2(n17043), .B1(n3434), .B2(n17046), .ZN(
        U239_Z_0) );
  OAI22_X1 U3411 ( .A1(n5588), .A2(n17048), .B1(n3434), .B2(n17051), .ZN(
        U238_Z_0) );
  OAI22_X1 U3414 ( .A1(n5587), .A2(n17053), .B1(n3434), .B2(n17056), .ZN(
        U237_Z_0) );
  OAI22_X1 U3417 ( .A1(n5586), .A2(n17058), .B1(n3434), .B2(n17061), .ZN(
        U236_Z_0) );
  NOR2_X1 U3420 ( .A1(n3441), .A2(n3444), .ZN(n3445) );
  INV_X1 U3421 ( .A(n3440), .ZN(n3444) );
  OAI22_X1 U3422 ( .A1(n5585), .A2(n17063), .B1(n3434), .B2(n17066), .ZN(
        U235_Z_0) );
  AND2_X1 U3425 ( .A1(n3447), .A2(n3448), .ZN(n3443) );
  OAI22_X1 U3426 ( .A1(n5584), .A2(n17068), .B1(n3434), .B2(n17071), .ZN(
        U234_Z_0) );
  AND2_X1 U3429 ( .A1(n3449), .A2(n3448), .ZN(n3438) );
  OAI22_X1 U3430 ( .A1(n4983), .A2(n17073), .B1(n3434), .B2(n17076), .ZN(
        U233_Z_0) );
  NOR2_X1 U3433 ( .A1(n3448), .A2(n3449), .ZN(n3435) );
  INV_X1 U3434 ( .A(n3447), .ZN(n3449) );
  OAI22_X1 U3435 ( .A1(n5583), .A2(n17078), .B1(n3434), .B2(n17081), .ZN(
        U232_Z_0) );
  AOI221_X1 U3437 ( .B1(n2495), .B2(n16705), .C1(n3450), .C2(n17007), .A(n3451), .ZN(n2103) );
  INV_X1 U3438 ( .A(n3452), .ZN(n3451) );
  AOI211_X1 U3439 ( .C1(n5803), .C2(n3453), .A(n2055), .B(n3454), .ZN(n3452)
         );
  NOR3_X1 U3440 ( .A1(n5803), .A2(n16992), .A3(n1685), .ZN(n3454) );
  OAI22_X1 U3441 ( .A1(n2131), .A2(n1685), .B1(n2501), .B2(n1649), .ZN(n3453)
         );
  INV_X1 U3442 ( .A(n1649), .ZN(n1685) );
  NAND4_X1 U3443 ( .A1(n3455), .A2(n3456), .A3(n3457), .A4(n3458), .ZN(n1649)
         );
  AOI222_X1 U3444 ( .A1(n16975), .A2(vis_msp_o[21]), .B1(n16970), .B2(n3254), 
        .C1(n16969), .C2(vis_psp_o[21]), .ZN(n3458) );
  AOI222_X1 U3446 ( .A1(n16984), .A2(vis_r14_o[23]), .B1(n16964), .B2(
        vis_r12_o[23]), .C1(n16987), .C2(vis_r11_o[23]), .ZN(n3457) );
  AOI222_X1 U3449 ( .A1(n16981), .A2(vis_r9_o[23]), .B1(n16961), .B2(
        vis_r10_o[23]), .C1(n16960), .C2(vis_r8_o[23]), .ZN(n3456) );
  AOI22_X1 U3451 ( .A1(n16978), .A2(n2515), .B1(n16956), .B2(n2713), .ZN(n3455) );
  XOR2_X1 U3455 ( .A(n16990), .B(n3467), .Z(n5803) );
  AOI221_X1 U3456 ( .B1(n2716), .B2(n16683), .C1(n16988), .C2(n3450), .A(n3468), .ZN(n3467) );
  NAND2_X1 U3457 ( .A1(n3469), .A2(n2719), .ZN(n3468) );
  NAND3_X1 U3458 ( .A1(n5254), .A2(n2198), .A3(n16807), .ZN(n3469) );
  INV_X1 U3460 ( .A(n2544), .ZN(n2495) );
  NOR2_X1 U3461 ( .A1(n17011), .A2(n2055), .ZN(n2544) );
  AOI221_X1 U3462 ( .B1(n2749), .B2(n2057), .C1(n2062), .C2(n2074), .A(n3470), 
        .ZN(n44) );
  INV_X1 U3463 ( .A(n3471), .ZN(n3470) );
  AOI221_X1 U3464 ( .B1(n2058), .B2(n2721), .C1(n2720), .C2(n2061), .A(n71), 
        .ZN(n3471) );
  AND4_X1 U3465 ( .A1(n3472), .A2(n3473), .A3(n3211), .A4(n3474), .ZN(n71) );
  NOR3_X1 U3466 ( .A1(n3425), .A2(n3433), .A3(n2074), .ZN(n3474) );
  INV_X1 U3467 ( .A(n3475), .ZN(n3433) );
  NAND2_X1 U3468 ( .A1(n3476), .A2(n3211), .ZN(n2720) );
  NAND2_X1 U3469 ( .A1(n2321), .A2(n3213), .ZN(n3211) );
  NOR2_X1 U3470 ( .A1(n3477), .A2(n3242), .ZN(n2321) );
  INV_X1 U3471 ( .A(n2341), .ZN(n3242) );
  NAND2_X1 U3472 ( .A1(n16830), .A2(n3478), .ZN(n2341) );
  NAND2_X1 U3473 ( .A1(n3472), .A2(n3285), .ZN(n2721) );
  OAI21_X1 U3474 ( .B1(n3213), .B2(n1027), .A(n3475), .ZN(n2749) );
  NOR2_X1 U3477 ( .A1(n3447), .A2(n3448), .ZN(n3439) );
  NAND3_X1 U3478 ( .A1(n17123), .A2(n3479), .A3(n1350), .ZN(n3448) );
  AOI221_X1 U3479 ( .B1(n3480), .B2(n3481), .C1(n1353), .C2(n3482), .A(n3483), 
        .ZN(n1350) );
  OAI21_X1 U3480 ( .B1(n3484), .B2(n5003), .A(n3485), .ZN(n3483) );
  OAI211_X1 U3481 ( .C1(n5162), .C2(n3484), .A(n3486), .B(n3487), .ZN(n3447)
         );
  AOI22_X1 U3482 ( .A1(n3481), .A2(n3488), .B1(n3482), .B2(n3489), .ZN(n3487)
         );
  INV_X1 U3483 ( .A(n3490), .ZN(n3484) );
  NOR2_X1 U3484 ( .A1(n3440), .A2(n3441), .ZN(n3446) );
  NAND3_X1 U3485 ( .A1(n3486), .A2(n3485), .A3(n3491), .ZN(n3441) );
  AOI222_X1 U3486 ( .A1(n3490), .A2(n2731), .B1(n3481), .B2(n3492), .C1(n3482), 
        .C2(n3493), .ZN(n3491) );
  NAND3_X1 U3487 ( .A1(n3486), .A2(n3485), .A3(n3494), .ZN(n3440) );
  AOI222_X1 U3488 ( .A1(n3490), .A2(n1723), .B1(n3481), .B2(n3495), .C1(n3482), 
        .C2(n3496), .ZN(n3494) );
  OAI211_X1 U3489 ( .C1(n16854), .C2(n699), .A(n3497), .B(n3498), .ZN(n3482)
         );
  NAND4_X1 U3490 ( .A1(n611), .A2(n757), .A3(n16839), .A4(n16867), .ZN(n3498)
         );
  INV_X1 U3491 ( .A(n1211), .ZN(n611) );
  NAND2_X1 U3492 ( .A1(n16845), .A2(n16851), .ZN(n1211) );
  NAND4_X1 U3493 ( .A1(n998), .A2(n1262), .A3(n16868), .A4(n16833), .ZN(n3497)
         );
  NAND4_X1 U3495 ( .A1(n3499), .A2(n759), .A3(n3500), .A4(n3501), .ZN(n3481)
         );
  AOI221_X1 U3496 ( .B1(n998), .B2(n16853), .C1(n529), .C2(n16847), .A(n3502), 
        .ZN(n3501) );
  AOI21_X1 U3497 ( .B1(n1868), .B2(n16833), .A(n3503), .ZN(n3500) );
  AOI211_X1 U3498 ( .C1(n918), .C2(n3504), .A(n16866), .B(n16845), .ZN(n3503)
         );
  NAND2_X1 U3499 ( .A1(n16825), .A2(n16806), .ZN(n3504) );
  INV_X1 U3500 ( .A(n723), .ZN(n1868) );
  NAND2_X1 U3501 ( .A1(n483), .A2(n16838), .ZN(n723) );
  NAND2_X1 U3502 ( .A1(n501), .A2(n16855), .ZN(n759) );
  OAI211_X1 U3503 ( .C1(n3505), .C2(n3506), .A(n653), .B(n568), .ZN(n3499) );
  NOR2_X1 U3504 ( .A1(n1086), .A2(n16826), .ZN(n3505) );
  OAI221_X1 U3505 ( .B1(n16869), .B2(n3507), .C1(n1519), .C2(n1580), .A(n3508), 
        .ZN(n3490) );
  NOR2_X1 U3506 ( .A1(n3509), .A2(n3510), .ZN(n3508) );
  NOR3_X1 U3507 ( .A1(n715), .A2(n16845), .A3(n16824), .ZN(n3510) );
  AOI222_X1 U3508 ( .A1(n760), .A2(n16867), .B1(n751), .B2(n16858), .C1(n563), 
        .C2(n16836), .ZN(n3507) );
  INV_X1 U3509 ( .A(n648), .ZN(n751) );
  NAND2_X1 U3510 ( .A1(n16866), .A2(n16856), .ZN(n648) );
  AOI21_X1 U3511 ( .B1(n16859), .B2(n2049), .A(n2631), .ZN(n3485) );
  INV_X1 U3512 ( .A(n1334), .ZN(n2631) );
  NAND2_X1 U3513 ( .A1(n16838), .A2(n16831), .ZN(n1334) );
  INV_X1 U3514 ( .A(n3363), .ZN(n2049) );
  NAND2_X1 U3515 ( .A1(n3430), .A2(n16870), .ZN(n3363) );
  AND3_X1 U3516 ( .A1(n3479), .A2(n713), .A3(n17122), .ZN(n3486) );
  NAND3_X1 U3517 ( .A1(n3511), .A2(n3512), .A3(n3513), .ZN(n3479) );
  NOR4_X1 U3518 ( .A1(n3514), .A2(n3515), .A3(n784), .A4(n3516), .ZN(n3513) );
  NOR4_X1 U3519 ( .A1(n16808), .A2(n556), .A3(n568), .A4(n755), .ZN(n3515) );
  OAI221_X1 U3520 ( .B1(n3517), .B2(n585), .C1(n3518), .C2(n3519), .A(n3520), 
        .ZN(n3514) );
  NAND3_X1 U3521 ( .A1(n909), .A2(n16862), .A3(n1042), .ZN(n3520) );
  AOI211_X1 U3522 ( .C1(n1042), .C2(n827), .A(n16833), .B(n3521), .ZN(n3519)
         );
  NOR3_X1 U3523 ( .A1(n617), .A2(n1086), .A3(n1023), .ZN(n3521) );
  AOI211_X1 U3524 ( .C1(n1605), .C2(n897), .A(n3522), .B(n16829), .ZN(n3518)
         );
  OAI33_X1 U3525 ( .A1(n617), .A2(n1519), .A3(n16805), .B1(n849), .B2(n1104), 
        .B3(n16826), .ZN(n3522) );
  INV_X1 U3526 ( .A(n912), .ZN(n1605) );
  NAND2_X1 U3527 ( .A1(n565), .A2(n16851), .ZN(n912) );
  AOI22_X1 U3528 ( .A1(n812), .A2(n3430), .B1(n1946), .B2(n16824), .ZN(n3517)
         );
  INV_X1 U3529 ( .A(n2689), .ZN(n812) );
  NAND2_X1 U3530 ( .A1(n16680), .A2(n16690), .ZN(n2689) );
  AOI222_X1 U3531 ( .A1(n757), .A2(n3523), .B1(n3524), .B2(n16839), .C1(n563), 
        .C2(n3525), .ZN(n3512) );
  OAI211_X1 U3532 ( .C1(n3526), .C2(n17096), .A(n3527), .B(n3528), .ZN(n3525)
         );
  NAND3_X1 U3533 ( .A1(n566), .A2(n16848), .A3(n997), .ZN(n3527) );
  AOI21_X1 U3534 ( .B1(n1034), .B2(n16680), .A(n1803), .ZN(n3526) );
  OAI22_X1 U3535 ( .A1(n917), .A2(n758), .B1(n3529), .B2(n16821), .ZN(n3524)
         );
  AOI21_X1 U3536 ( .B1(n608), .B2(n16856), .A(n1207), .ZN(n3529) );
  INV_X1 U3537 ( .A(n1027), .ZN(n1207) );
  OAI221_X1 U3538 ( .B1(n16841), .B2(n568), .C1(n16866), .C2(n673), .A(n3530), 
        .ZN(n3523) );
  AOI221_X1 U3539 ( .B1(n3432), .B2(n16826), .C1(n3531), .C2(n16836), .A(n1564), .ZN(n3530) );
  NOR2_X1 U3540 ( .A1(n16845), .A2(n16830), .ZN(n3531) );
  INV_X1 U3541 ( .A(n3429), .ZN(n3432) );
  NAND2_X1 U3542 ( .A1(n16845), .A2(n16849), .ZN(n3429) );
  AOI222_X1 U3543 ( .A1(n506), .A2(n565), .B1(n827), .B2(n785), .C1(n2661), 
        .C2(n3532), .ZN(n3511) );
  INV_X1 U3544 ( .A(n524), .ZN(n785) );
  NAND2_X1 U3545 ( .A1(n16826), .A2(n17096), .ZN(n524) );
  OAI22_X1 U3546 ( .A1(n4948), .A2(n2085), .B1(n3533), .B2(n2087), .ZN(
        U229_Z_0) );
  INV_X1 U3547 ( .A(n2085), .ZN(n2087) );
  AOI222_X1 U3548 ( .A1(n88), .A2(n3534), .B1(n86), .B2(n2077), .C1(n1510), 
        .C2(n84), .ZN(n3533) );
  AOI22_X1 U3549 ( .A1(n2102), .A2(n4947), .B1(n1759), .B2(n1783), .ZN(n1510)
         );
  INV_X1 U3550 ( .A(n3535), .ZN(n1783) );
  OAI221_X1 U3551 ( .B1(n3092), .B2(n2376), .C1(n2375), .C2(n3477), .A(n3536), 
        .ZN(n3535) );
  AOI22_X1 U3552 ( .A1(n3537), .A2(n3538), .B1(n2322), .B2(n1787), .ZN(n3536)
         );
  OAI22_X1 U3553 ( .A1(n1789), .A2(n3539), .B1(n1791), .B2(n2390), .ZN(n3537)
         );
  INV_X1 U3554 ( .A(n2078), .ZN(n2102) );
  OAI211_X1 U3555 ( .C1(n94), .C2(n3540), .A(n3541), .B(n3542), .ZN(n2078) );
  AOI222_X1 U3556 ( .A1(n2125), .A2(vis_apsr_o[3]), .B1(n17008), .B2(n3534), 
        .C1(n16688), .C2(n17009), .ZN(n3542) );
  OAI22_X1 U3557 ( .A1(n16957), .A2(n3543), .B1(n4950), .B2(n3544), .ZN(n2015)
         );
  AOI221_X1 U3558 ( .B1(n1041), .B2(n16690), .C1(n16823), .C2(n3545), .A(n1095), .ZN(n3544) );
  OAI211_X1 U3559 ( .C1(n16829), .C2(n3546), .A(n1233), .B(n1023), .ZN(n3545)
         );
  INV_X1 U3560 ( .A(n1043), .ZN(n1041) );
  NAND2_X1 U3561 ( .A1(n16851), .A2(n16860), .ZN(n1043) );
  OAI21_X1 U3563 ( .B1(n543), .B2(n3547), .A(n1697), .ZN(n2243) );
  NOR2_X1 U3564 ( .A1(n1218), .A2(n532), .ZN(n3547) );
  NAND2_X1 U3565 ( .A1(n16806), .A2(n16855), .ZN(n1218) );
  NAND2_X1 U3567 ( .A1(n914), .A2(n16831), .ZN(n713) );
  NOR3_X1 U3569 ( .A1(n16656), .A2(n16671), .A3(n2168), .ZN(n2125) );
  NAND4_X1 U3570 ( .A1(n2662), .A2(n16868), .A3(n1574), .A4(n1697), .ZN(n2168)
         );
  INV_X1 U3571 ( .A(n606), .ZN(n2662) );
  NAND2_X1 U3572 ( .A1(n16862), .A2(n16856), .ZN(n606) );
  AOI21_X1 U3573 ( .B1(n3548), .B2(n1513), .A(n2055), .ZN(n3541) );
  NAND3_X1 U3575 ( .A1(n16829), .A2(n1697), .A3(n1034), .ZN(n2124) );
  NOR2_X1 U3576 ( .A1(U186_Z_0), .A2(n16993), .ZN(n3548) );
  NAND2_X1 U3578 ( .A1(n3549), .A2(n2501), .ZN(n2127) );
  AOI22_X1 U3579 ( .A1(n1513), .A2(n2126), .B1(n1872), .B2(n16995), .ZN(n3540)
         );
  INV_X1 U3582 ( .A(n1513), .ZN(n1872) );
  OAI221_X1 U3584 ( .B1(n1803), .B2(n515), .C1(n501), .C2(n16829), .A(n16845), 
        .ZN(n3550) );
  INV_X1 U3585 ( .A(n3551), .ZN(n3549) );
  OAI22_X1 U3586 ( .A1(n16957), .A2(n2628), .B1(n4950), .B2(n3552), .ZN(n3551)
         );
  AOI211_X1 U3587 ( .C1(n884), .C2(n16826), .A(n3553), .B(n3554), .ZN(n3552)
         );
  NOR3_X1 U3588 ( .A1(n16826), .A2(n16858), .A3(n1519), .ZN(n3554) );
  OAI21_X1 U3589 ( .B1(n16820), .B2(n818), .A(n3555), .ZN(n3553) );
  INV_X1 U3590 ( .A(n3502), .ZN(n3555) );
  OAI21_X1 U3591 ( .B1(n762), .B2(n3556), .A(n1541), .ZN(n3502) );
  NAND2_X1 U3592 ( .A1(n998), .A2(n16821), .ZN(n3556) );
  INV_X1 U3593 ( .A(n860), .ZN(n998) );
  NAND2_X1 U3594 ( .A1(n16825), .A2(n16845), .ZN(n860) );
  NAND2_X1 U3595 ( .A1(n914), .A2(n16838), .ZN(n818) );
  NOR2_X1 U3596 ( .A1(n532), .A2(n16862), .ZN(n884) );
  INV_X1 U3597 ( .A(n3543), .ZN(n2628) );
  OAI22_X1 U3598 ( .A1(n3557), .A2(n795), .B1(n5100), .B2(n3558), .ZN(n3543)
         );
  AOI22_X1 U3599 ( .A1(n3559), .A2(n16671), .B1(n16810), .B2(n3560), .ZN(n3558) );
  OAI33_X1 U3600 ( .A1(n3561), .A2(n3562), .A3(n3563), .B1(n3564), .B2(n16809), 
        .B3(n3565), .ZN(n3560) );
  AOI221_X1 U3601 ( .B1(n3255), .B2(n1821), .C1(n3348), .C2(n3566), .A(n3567), 
        .ZN(n3565) );
  INV_X1 U3602 ( .A(n2764), .ZN(n3255) );
  OAI22_X1 U3603 ( .A1(n3349), .A2(n1900), .B1(n3256), .B2(n1820), .ZN(n3564)
         );
  INV_X1 U3604 ( .A(n2809), .ZN(n3256) );
  NOR2_X1 U3605 ( .A1(n3346), .A2(n1900), .ZN(n3563) );
  AOI221_X1 U3606 ( .B1(n3251), .B2(n1821), .C1(n3345), .C2(n3566), .A(n3567), 
        .ZN(n3562) );
  INV_X1 U3607 ( .A(n2507), .ZN(n3251) );
  OAI21_X1 U3608 ( .B1(n3252), .B2(n1820), .A(n16809), .ZN(n3561) );
  INV_X1 U3609 ( .A(n2705), .ZN(n3252) );
  OAI33_X1 U3610 ( .A1(n3568), .A2(n3569), .A3(n3570), .B1(n3571), .B2(n16809), 
        .B3(n3572), .ZN(n3559) );
  AOI221_X1 U3611 ( .B1(n3239), .B2(n1821), .C1(n3319), .C2(n3566), .A(n3567), 
        .ZN(n3572) );
  INV_X1 U3612 ( .A(n2585), .ZN(n3239) );
  OAI22_X1 U3613 ( .A1(n3280), .A2(n1900), .B1(n3240), .B2(n1820), .ZN(n3571)
         );
  INV_X1 U3614 ( .A(n3199), .ZN(n3240) );
  NOR2_X1 U3615 ( .A1(n3315), .A2(n1900), .ZN(n3570) );
  AOI221_X1 U3616 ( .B1(n3231), .B2(n1821), .C1(n3314), .C2(n3566), .A(n3567), 
        .ZN(n3569) );
  INV_X1 U3617 ( .A(n3317), .ZN(n3231) );
  OAI21_X1 U3618 ( .B1(n3233), .B2(n1820), .A(n16809), .ZN(n3568) );
  INV_X1 U3619 ( .A(n2531), .ZN(n3233) );
  AOI22_X1 U3620 ( .A1(n3573), .A2(n16671), .B1(n16810), .B2(n3574), .ZN(n3557) );
  OAI33_X1 U3621 ( .A1(n3575), .A2(n3576), .A3(n3577), .B1(n3578), .B2(n16809), 
        .B3(n3579), .ZN(n3574) );
  AOI221_X1 U3622 ( .B1(n3338), .B2(n3566), .C1(n3281), .C2(n1821), .A(n3567), 
        .ZN(n3579) );
  INV_X1 U3623 ( .A(n2271), .ZN(n3281) );
  OAI22_X1 U3624 ( .A1(n3282), .A2(n1820), .B1(n3339), .B2(n1900), .ZN(n3578)
         );
  INV_X1 U3625 ( .A(n2452), .ZN(n3282) );
  NOR2_X1 U3626 ( .A1(n3398), .A2(n1820), .ZN(n3577) );
  INV_X1 U3627 ( .A(n2297), .ZN(n3398) );
  AOI221_X1 U3628 ( .B1(n3278), .B2(n3566), .C1(n2183), .C2(n1821), .A(n3567), 
        .ZN(n3576) );
  INV_X1 U3629 ( .A(n3274), .ZN(n2183) );
  OAI21_X1 U3630 ( .B1(n3341), .B2(n1900), .A(n16809), .ZN(n3575) );
  OAI33_X1 U3631 ( .A1(n3580), .A2(n3581), .A3(n3582), .B1(n3583), .B2(n16809), 
        .B3(n3584), .ZN(n3573) );
  AOI221_X1 U3632 ( .B1(n3261), .B2(n1821), .C1(n3328), .C2(n3566), .A(n3567), 
        .ZN(n3584) );
  INV_X1 U3633 ( .A(n3041), .ZN(n3261) );
  OAI22_X1 U3634 ( .A1(n3329), .A2(n1900), .B1(n3262), .B2(n1820), .ZN(n3583)
         );
  INV_X1 U3635 ( .A(n3155), .ZN(n3262) );
  NOR2_X1 U3636 ( .A1(n3333), .A2(n1900), .ZN(n3582) );
  INV_X1 U3638 ( .A(n3022), .ZN(n3333) );
  AOI221_X1 U3639 ( .B1(n3264), .B2(n1821), .C1(n3332), .C2(n3566), .A(n3567), 
        .ZN(n3581) );
  AND2_X1 U3640 ( .A1(n1821), .A2(n3566), .ZN(n3567) );
  INV_X1 U3643 ( .A(n2856), .ZN(n3264) );
  OAI21_X1 U3644 ( .B1(n3265), .B2(n1820), .A(n16809), .ZN(n3580) );
  NAND4_X1 U3647 ( .A1(n3585), .A2(n3586), .A3(n3587), .A4(n3588), .ZN(n1513)
         );
  AOI222_X1 U3648 ( .A1(n16964), .A2(vis_r12_o[31]), .B1(n16969), .B2(
        vis_psp_o[29]), .C1(n16975), .C2(vis_msp_o[29]), .ZN(n3588) );
  NAND3_X1 U3653 ( .A1(n4978), .A2(n5036), .A3(n3593), .ZN(n2182) );
  AOI222_X1 U3654 ( .A1(n16961), .A2(vis_r10_o[31]), .B1(n16987), .B2(
        vis_r11_o[31]), .C1(n16984), .C2(vis_r14_o[31]), .ZN(n3587) );
  NOR2_X1 U3657 ( .A1(n2184), .A2(n3597), .ZN(n3593) );
  NAND3_X1 U3661 ( .A1(n4978), .A2(n3480), .A3(n3598), .ZN(n2191) );
  AOI222_X1 U3662 ( .A1(n16970), .A2(n3400), .B1(n16960), .B2(vis_r8_o[31]), 
        .C1(n16981), .C2(vis_r9_o[31]), .ZN(n3586) );
  NAND2_X1 U3664 ( .A1(n3598), .A2(n3592), .ZN(n2637) );
  NAND3_X1 U3667 ( .A1(n4978), .A2(n5036), .A3(n3598), .ZN(n2190) );
  NOR3_X1 U3668 ( .A1(n3492), .A2(n4959), .A3(n2184), .ZN(n3598) );
  NAND2_X1 U3670 ( .A1(n16957), .A2(n3601), .ZN(n2184) );
  AOI22_X1 U3672 ( .A1(n16976), .A2(n867), .B1(n16956), .B2(n874), .ZN(n3585)
         );
  NOR4_X1 U3676 ( .A1(n727), .A2(n3602), .A3(n3603), .A4(n3604), .ZN(n3601) );
  OAI221_X1 U3677 ( .B1(n989), .B2(n3221), .C1(n16806), .C2(n1086), .A(n3605), 
        .ZN(n3604) );
  OAI21_X1 U3678 ( .B1(n991), .B2(n527), .A(n16845), .ZN(n3605) );
  INV_X1 U3679 ( .A(n1300), .ZN(n3221) );
  NOR2_X1 U3680 ( .A1(n16839), .A2(n16848), .ZN(n1300) );
  OAI33_X1 U3681 ( .A1(n715), .A2(n16871), .A3(n604), .B1(n3597), .B2(n4978), 
        .B3(n5036), .ZN(n3603) );
  NAND2_X1 U3682 ( .A1(n3492), .A2(n3495), .ZN(n3597) );
  NOR3_X1 U3683 ( .A1(n994), .A2(n16836), .A3(n16826), .ZN(n3602) );
  INV_X1 U3684 ( .A(n1946), .ZN(n994) );
  NOR2_X1 U3685 ( .A1(n1234), .A2(n16848), .ZN(n1946) );
  INV_X1 U3686 ( .A(n891), .ZN(n727) );
  OAI21_X1 U3687 ( .B1(n16821), .B2(n1177), .A(n3606), .ZN(n2222) );
  NAND3_X1 U3688 ( .A1(n3430), .A2(n16871), .A3(n1034), .ZN(n3606) );
  NAND4_X1 U3689 ( .A1(n597), .A2(n1805), .A3(n991), .A4(n16856), .ZN(n1177)
         );
  INV_X1 U3690 ( .A(U186_Z_0), .ZN(n94) );
  INV_X1 U3691 ( .A(n28), .ZN(n2077) );
  AOI221_X1 U3692 ( .B1(n2061), .B2(n2067), .C1(n2057), .C2(n2072), .A(n3607), 
        .ZN(n28) );
  INV_X1 U3693 ( .A(n3608), .ZN(n3607) );
  AOI221_X1 U3694 ( .B1(n2069), .B2(n2062), .C1(n2074), .C2(n2058), .A(n2076), 
        .ZN(n3608) );
  NAND4_X1 U3697 ( .A1(n3216), .A2(n3092), .A3(n3610), .A4(n3611), .ZN(n3209)
         );
  AOI222_X1 U3698 ( .A1(n3532), .A2(n3612), .B1(n3613), .B2(n1564), .C1(n3614), 
        .C2(n2062), .ZN(n3611) );
  OAI21_X1 U3699 ( .B1(n3615), .B2(n16859), .A(n1233), .ZN(n3614) );
  AOI21_X1 U3700 ( .B1(n5227), .B2(n5102), .A(n16842), .ZN(n3615) );
  NOR2_X1 U3701 ( .A1(n3616), .A2(n16839), .ZN(n3613) );
  OAI21_X1 U3702 ( .B1(n5227), .B2(n3616), .A(n3617), .ZN(n3612) );
  NAND3_X1 U3703 ( .A1(n2061), .A2(n3223), .A3(n5227), .ZN(n3617) );
  AOI22_X1 U3704 ( .A1(n3223), .A2(n2057), .B1(n2058), .B2(n5102), .ZN(n3616)
         );
  INV_X1 U3706 ( .A(n917), .ZN(n3532) );
  NAND2_X1 U3707 ( .A1(n16845), .A2(n16862), .ZN(n917) );
  NAND4_X1 U3708 ( .A1(n2058), .A2(n16847), .A3(n16858), .A4(n16867), .ZN(
        n3610) );
  INV_X1 U3709 ( .A(n3473), .ZN(n3609) );
  OAI211_X1 U3710 ( .C1(n16862), .C2(n1104), .A(n3215), .B(n3618), .ZN(n3473)
         );
  NOR2_X1 U3711 ( .A1(n3619), .A2(n3620), .ZN(n3618) );
  NOR3_X1 U3712 ( .A1(n673), .A2(n16868), .A3(n16854), .ZN(n3620) );
  INV_X1 U3713 ( .A(n3216), .ZN(n3619) );
  NAND2_X1 U3714 ( .A1(hresp_i), .A2(n2882), .ZN(n3216) );
  OR3_X1 U3715 ( .A1(n2359), .A2(n2322), .A3(n2323), .ZN(n2376) );
  AOI21_X1 U3716 ( .B1(n3539), .B2(n2390), .A(n2389), .ZN(n2323) );
  INV_X1 U3717 ( .A(n3477), .ZN(n2359) );
  NAND3_X1 U3718 ( .A1(n3621), .A2(n3622), .A3(n3623), .ZN(n2058) );
  AOI221_X1 U3719 ( .B1(hrdata_i[15]), .B2(n2879), .C1(n2922), .C2(n3624), .A(
        n3625), .ZN(n3623) );
  OAI22_X1 U3720 ( .A1(n2981), .A2(n282), .B1(n5505), .B2(n16685), .ZN(n3625)
         );
  INV_X1 U3722 ( .A(n1791), .ZN(n3624) );
  OAI22_X1 U3723 ( .A1(n16789), .A2(n2384), .B1(n2337), .B2(n2354), .ZN(n1791)
         );
  OAI221_X1 U3724 ( .B1(n3346), .B2(n16950), .C1(n3348), .C2(n16953), .A(n3626), .ZN(n2354) );
  AOI22_X1 U3725 ( .A1(n16947), .A2(n2764), .B1(n16942), .B2(n2705), .ZN(n3626) );
  NAND3_X1 U3726 ( .A1(n3627), .A2(n3628), .A3(n3629), .ZN(n2705) );
  AOI221_X1 U3727 ( .B1(n16941), .B2(vis_r2_o[22]), .C1(n16938), .C2(
        vis_r0_o[22]), .A(n3634), .ZN(n3629) );
  OAI22_X1 U3728 ( .A1(n5050), .A2(n16935), .B1(n5436), .B2(n16932), .ZN(n3634) );
  AOI22_X1 U3730 ( .A1(n16929), .A2(vis_r5_o[22]), .B1(n16926), .B2(
        vis_r4_o[22]), .ZN(n3628) );
  AOI22_X1 U3731 ( .A1(n16923), .A2(vis_r6_o[22]), .B1(n16920), .B2(
        vis_r1_o[22]), .ZN(n3627) );
  NAND3_X1 U3734 ( .A1(n3645), .A2(n3646), .A3(n3647), .ZN(n2764) );
  AOI221_X1 U3735 ( .B1(n16941), .B2(vis_r2_o[20]), .C1(n16938), .C2(
        vis_r0_o[20]), .A(n3650), .ZN(n3647) );
  OAI22_X1 U3736 ( .A1(n5613), .A2(n16935), .B1(n5605), .B2(n16932), .ZN(n3650) );
  AOI22_X1 U3738 ( .A1(n16929), .A2(vis_r5_o[20]), .B1(n16926), .B2(
        vis_r4_o[20]), .ZN(n3646) );
  AOI22_X1 U3739 ( .A1(n16923), .A2(vis_r6_o[20]), .B1(n16920), .B2(
        vis_r1_o[20]), .ZN(n3645) );
  INV_X1 U3742 ( .A(n2787), .ZN(n3348) );
  NAND3_X1 U3743 ( .A1(n3655), .A2(n3656), .A3(n3657), .ZN(n2787) );
  AOI221_X1 U3744 ( .B1(n16941), .B2(vis_r2_o[19]), .C1(n16938), .C2(
        vis_r0_o[19]), .A(n3660), .ZN(n3657) );
  OAI22_X1 U3745 ( .A1(n5090), .A2(n16935), .B1(n5438), .B2(n16932), .ZN(n3660) );
  AOI22_X1 U3747 ( .A1(n16929), .A2(vis_r5_o[19]), .B1(n16926), .B2(
        vis_r4_o[19]), .ZN(n3656) );
  AOI22_X1 U3748 ( .A1(n16923), .A2(vis_r6_o[19]), .B1(n16920), .B2(
        vis_r1_o[19]), .ZN(n3655) );
  INV_X1 U3751 ( .A(n2738), .ZN(n3346) );
  NAND3_X1 U3752 ( .A1(n3665), .A2(n3666), .A3(n3667), .ZN(n2738) );
  AOI221_X1 U3753 ( .B1(n16941), .B2(vis_r2_o[21]), .C1(n16938), .C2(
        vis_r0_o[21]), .A(n3670), .ZN(n3667) );
  OAI22_X1 U3754 ( .A1(n5117), .A2(n16935), .B1(n5437), .B2(n16932), .ZN(n3670) );
  AOI22_X1 U3756 ( .A1(n16929), .A2(vis_r5_o[21]), .B1(n16926), .B2(
        vis_r4_o[21]), .ZN(n3666) );
  AOI22_X1 U3757 ( .A1(n16923), .A2(vis_r6_o[21]), .B1(n16920), .B2(
        vis_r1_o[21]), .ZN(n3665) );
  OAI221_X1 U3760 ( .B1(n3349), .B2(n16950), .C1(n3332), .C2(n16953), .A(n3675), .ZN(n2384) );
  AOI22_X1 U3761 ( .A1(n16947), .A2(n2856), .B1(n16942), .B2(n2809), .ZN(n3675) );
  NAND3_X1 U3762 ( .A1(n3676), .A2(n3677), .A3(n3678), .ZN(n2809) );
  AOI221_X1 U3763 ( .B1(n16941), .B2(vis_r2_o[18]), .C1(n16938), .C2(
        vis_r0_o[18]), .A(n3681), .ZN(n3678) );
  OAI22_X1 U3764 ( .A1(n5064), .A2(n16935), .B1(n5439), .B2(n16932), .ZN(n3681) );
  AOI22_X1 U3766 ( .A1(n16929), .A2(vis_r5_o[18]), .B1(n16926), .B2(
        vis_r4_o[18]), .ZN(n3677) );
  AOI22_X1 U3767 ( .A1(n16923), .A2(vis_r6_o[18]), .B1(n16920), .B2(
        vis_r1_o[18]), .ZN(n3676) );
  NAND3_X1 U3770 ( .A1(n3686), .A2(n3687), .A3(n3688), .ZN(n2856) );
  AOI221_X1 U3771 ( .B1(n16941), .B2(vis_r2_o[16]), .C1(n16938), .C2(
        vis_r0_o[16]), .A(n3691), .ZN(n3688) );
  OAI22_X1 U3772 ( .A1(n5071), .A2(n16935), .B1(n5441), .B2(n16932), .ZN(n3691) );
  AOI22_X1 U3774 ( .A1(n16929), .A2(vis_r5_o[16]), .B1(n16926), .B2(
        vis_r4_o[16]), .ZN(n3687) );
  AOI22_X1 U3775 ( .A1(n16923), .A2(vis_r6_o[16]), .B1(n16920), .B2(
        vis_r1_o[16]), .ZN(n3686) );
  INV_X1 U3778 ( .A(n3267), .ZN(n3332) );
  NAND3_X1 U3779 ( .A1(n3696), .A2(n3697), .A3(n3698), .ZN(n3267) );
  AOI221_X1 U3780 ( .B1(n16941), .B2(vis_r2_o[15]), .C1(n16938), .C2(
        vis_r0_o[15]), .A(n3701), .ZN(n3698) );
  OAI22_X1 U3781 ( .A1(n5110), .A2(n16935), .B1(n5449), .B2(n16932), .ZN(n3701) );
  AOI22_X1 U3783 ( .A1(n16929), .A2(vis_r5_o[15]), .B1(n16926), .B2(
        vis_r4_o[15]), .ZN(n3697) );
  AOI22_X1 U3784 ( .A1(n16923), .A2(vis_r6_o[15]), .B1(n16920), .B2(
        vis_r1_o[15]), .ZN(n3696) );
  INV_X1 U3787 ( .A(n2833), .ZN(n3349) );
  NAND3_X1 U3788 ( .A1(n3706), .A2(n3707), .A3(n3708), .ZN(n2833) );
  AOI221_X1 U3789 ( .B1(n16941), .B2(vis_r2_o[17]), .C1(n16938), .C2(
        vis_r0_o[17]), .A(n3711), .ZN(n3708) );
  OAI22_X1 U3790 ( .A1(n5085), .A2(n16935), .B1(n5440), .B2(n16932), .ZN(n3711) );
  AOI22_X1 U3792 ( .A1(n16929), .A2(vis_r5_o[17]), .B1(n16926), .B2(
        vis_r4_o[17]), .ZN(n3707) );
  AOI22_X1 U3793 ( .A1(n16923), .A2(vis_r6_o[17]), .B1(n16920), .B2(
        vis_r1_o[17]), .ZN(n3706) );
  AOI221_X1 U3796 ( .B1(n2895), .B2(n416), .C1(n2882), .C2(n3716), .A(n2897), 
        .ZN(n3622) );
  INV_X1 U3797 ( .A(n3247), .ZN(n2897) );
  NAND4_X1 U3798 ( .A1(n4905), .A2(n3717), .A3(n2882), .A4(n5017), .ZN(n3247)
         );
  OAI221_X1 U3799 ( .B1(n5150), .B2(n2898), .C1(n5156), .C2(n2899), .A(n3718), 
        .ZN(n3716) );
  AOI22_X1 U3800 ( .A1(n1897), .A2(n3719), .B1(n1893), .B2(n3720), .ZN(n3718)
         );
  INV_X1 U3801 ( .A(n424), .ZN(n416) );
  NAND2_X1 U3802 ( .A1(n2905), .A2(n3721), .ZN(n424) );
  NAND3_X1 U3803 ( .A1(n2908), .A2(n1372), .A3(n2907), .ZN(n3721) );
  NOR3_X1 U3804 ( .A1(n3066), .A2(n1067), .A3(n1066), .ZN(n2905) );
  NOR3_X1 U3805 ( .A1(n3722), .A2(n2907), .A3(n1370), .ZN(n1067) );
  INV_X1 U3806 ( .A(n1372), .ZN(n1370) );
  OAI21_X1 U3807 ( .B1(n3723), .B2(n209), .A(n3724), .ZN(n1372) );
  OAI221_X1 U3808 ( .B1(n3725), .B2(n1371), .C1(n2907), .C2(n3722), .A(n3726), 
        .ZN(n3724) );
  OAI21_X1 U3809 ( .B1(n3727), .B2(n3728), .A(n1368), .ZN(n3726) );
  OAI22_X1 U3810 ( .A1(n3722), .A2(n3729), .B1(n5098), .B2(n3730), .ZN(n1368)
         );
  INV_X1 U3811 ( .A(n3725), .ZN(n3728) );
  INV_X1 U3812 ( .A(n3727), .ZN(n1371) );
  AOI22_X1 U3813 ( .A1(n3731), .A2(n2903), .B1(n3732), .B2(n3723), .ZN(n3727)
         );
  NOR2_X1 U3814 ( .A1(n3733), .A2(n1369), .ZN(n3725) );
  OAI22_X1 U3815 ( .A1(n3734), .A2(n3722), .B1(n5097), .B2(n3730), .ZN(n1369)
         );
  INV_X1 U3816 ( .A(n1373), .ZN(n3733) );
  AOI22_X1 U3817 ( .A1(n2903), .A2(n4826), .B1(n5503), .B2(n3723), .ZN(n1373)
         );
  INV_X1 U3818 ( .A(n2903), .ZN(n3723) );
  OAI21_X1 U3819 ( .B1(n4802), .B2(n3735), .A(n1053), .ZN(n2903) );
  AOI22_X1 U3820 ( .A1(n3736), .A2(n4826), .B1(n4961), .B2(n3732), .ZN(n3735)
         );
  AOI21_X1 U3821 ( .B1(n5504), .B2(n3731), .A(n5503), .ZN(n3736) );
  AND2_X1 U3822 ( .A1(n3730), .A2(n3737), .ZN(n2907) );
  INV_X1 U3823 ( .A(n3730), .ZN(n3722) );
  OAI21_X1 U3824 ( .B1(n3738), .B2(n3739), .A(n203), .ZN(n3730) );
  OAI21_X1 U3826 ( .B1(n3729), .B2(n3740), .A(n3737), .ZN(n3739) );
  NAND3_X1 U3827 ( .A1(n2911), .A2(n2909), .A3(n3741), .ZN(n3737) );
  AOI22_X1 U3828 ( .A1(n3729), .A2(n3740), .B1(n3734), .B2(n2929), .ZN(n3738)
         );
  AOI22_X1 U3829 ( .A1(n3742), .A2(n2908), .B1(n3743), .B2(n2911), .ZN(n3734)
         );
  OAI22_X1 U3830 ( .A1(n2908), .A2(n3744), .B1(n3745), .B2(n2911), .ZN(n3729)
         );
  INV_X1 U3831 ( .A(n2911), .ZN(n2908) );
  OAI21_X1 U3832 ( .B1(n3746), .B2(n2997), .A(n3747), .ZN(n2911) );
  OAI221_X1 U3833 ( .B1(n3748), .B2(n3745), .C1(n2993), .C2(n3749), .A(n3750), 
        .ZN(n3747) );
  OAI21_X1 U3834 ( .B1(n3751), .B2(n3752), .A(n3744), .ZN(n3750) );
  OAI22_X1 U3835 ( .A1(n2993), .A2(n3753), .B1(n3754), .B2(n2909), .ZN(n3744)
         );
  INV_X1 U3836 ( .A(n3748), .ZN(n3752) );
  INV_X1 U3837 ( .A(n3745), .ZN(n3751) );
  OAI22_X1 U3838 ( .A1(n3755), .A2(n2910), .B1(n3073), .B2(n3756), .ZN(n3745)
         );
  NOR2_X1 U3839 ( .A1(n3757), .A2(n3743), .ZN(n3748) );
  OAI22_X1 U3840 ( .A1(n3758), .A2(n2909), .B1(n3759), .B2(n2993), .ZN(n3743)
         );
  INV_X1 U3841 ( .A(n2909), .ZN(n2993) );
  NAND3_X1 U3843 ( .A1(n3764), .A2(n3759), .A3(n3765), .ZN(n3763) );
  AOI21_X1 U3844 ( .B1(n3766), .B2(n3754), .A(n3741), .ZN(n3765) );
  INV_X1 U3845 ( .A(n3749), .ZN(n3741) );
  INV_X1 U3846 ( .A(n3753), .ZN(n3766) );
  AOI22_X1 U3847 ( .A1(n2995), .A2(n3767), .B1(n3768), .B2(n3086), .ZN(n3759)
         );
  INV_X1 U3848 ( .A(n3758), .ZN(n3764) );
  INV_X1 U3849 ( .A(n2994), .ZN(n3761) );
  NAND2_X1 U3850 ( .A1(n3749), .A2(n3753), .ZN(n3760) );
  OAI22_X1 U3851 ( .A1(n3086), .A2(n3769), .B1(n3770), .B2(n2995), .ZN(n3753)
         );
  INV_X1 U3852 ( .A(n2995), .ZN(n3086) );
  NAND2_X1 U3853 ( .A1(n3771), .A2(n2995), .ZN(n3749) );
  OAI21_X1 U3854 ( .B1(n3771), .B2(n3772), .A(n3774), .ZN(n2995) );
  OAI21_X1 U3855 ( .B1(n244), .B2(n3775), .A(n3087), .ZN(n3774) );
  AOI22_X1 U3856 ( .A1(n3776), .A2(n3770), .B1(n3777), .B2(n3768), .ZN(n3772)
         );
  AOI22_X1 U3857 ( .A1(n3087), .A2(n5151), .B1(n1885), .B2(n3778), .ZN(n3768)
         );
  AOI21_X1 U3858 ( .B1(n3779), .B2(n3769), .A(n3767), .ZN(n3777) );
  AOI22_X1 U3859 ( .A1(n3088), .A2(n5154), .B1(n3780), .B2(n5152), .ZN(n3767)
         );
  INV_X1 U3860 ( .A(n3770), .ZN(n3779) );
  OAI22_X1 U3861 ( .A1(n5150), .A2(n3778), .B1(n5521), .B2(n3087), .ZN(n3770)
         );
  INV_X1 U3862 ( .A(n3778), .ZN(n3087) );
  NOR3_X1 U3863 ( .A1(n4795), .A2(n4749), .A3(n3781), .ZN(n3778) );
  AOI211_X1 U3864 ( .C1(n3782), .C2(n3783), .A(n244), .B(n3775), .ZN(n3781) );
  NAND2_X1 U3866 ( .A1(n3784), .A2(n5150), .ZN(n3783) );
  OAI211_X1 U3867 ( .C1(n3784), .C2(n5150), .A(n5151), .B(n4753), .ZN(n3782)
         );
  INV_X1 U3868 ( .A(n3769), .ZN(n3776) );
  OAI22_X1 U3869 ( .A1(n5155), .A2(n3780), .B1(n5153), .B2(n3088), .ZN(n3769)
         );
  AOI21_X1 U3870 ( .B1(n3785), .B2(n3786), .A(n3780), .ZN(n3771) );
  INV_X1 U3871 ( .A(n3088), .ZN(n3780) );
  OAI211_X1 U3872 ( .C1(n3787), .C2(n3788), .A(n2916), .B(n2914), .ZN(n3088)
         );
  NAND2_X1 U3875 ( .A1(n3785), .A2(n3786), .ZN(n3788) );
  AOI22_X1 U3876 ( .A1(n3789), .A2(n5154), .B1(n5155), .B2(n3790), .ZN(n3787)
         );
  AOI21_X1 U3877 ( .B1(n5153), .B2(n3791), .A(n5152), .ZN(n3789) );
  OAI222_X1 U3878 ( .A1(n3792), .A2(n3085), .B1(n3793), .B2(n3794), .C1(n3795), 
        .C2(n2994), .ZN(n3754) );
  OAI221_X1 U3879 ( .B1(n2932), .B2(n3085), .C1(n3796), .C2(n2994), .A(n3797), 
        .ZN(n3758) );
  NAND3_X1 U3880 ( .A1(n3798), .A2(n2994), .A3(n5158), .ZN(n3797) );
  NAND2_X1 U3881 ( .A1(n2994), .A2(n3794), .ZN(n3085) );
  NAND3_X1 U3882 ( .A1(n3799), .A2(n3800), .A3(n3801), .ZN(n2994) );
  OAI21_X1 U3883 ( .B1(n5578), .B2(n5011), .A(n3802), .ZN(n3801) );
  NAND3_X1 U3884 ( .A1(n3762), .A2(n3795), .A3(n3803), .ZN(n3800) );
  NAND2_X1 U3885 ( .A1(n3794), .A2(n3804), .ZN(n3762) );
  OAI21_X1 U3886 ( .B1(n3803), .B2(n3795), .A(n3805), .ZN(n3799) );
  OAI22_X1 U3887 ( .A1(n3793), .A2(n3794), .B1(n3792), .B2(n3804), .ZN(n3805)
         );
  INV_X1 U3888 ( .A(n3806), .ZN(n3804) );
  OAI22_X1 U3889 ( .A1(n5156), .A2(n3084), .B1(n5522), .B2(n3802), .ZN(n3795)
         );
  INV_X1 U3890 ( .A(n3807), .ZN(n3803) );
  OAI221_X1 U3891 ( .B1(n5158), .B2(n3794), .C1(n5160), .C2(n3798), .A(n3796), 
        .ZN(n3807) );
  AOI22_X1 U3892 ( .A1(n3802), .A2(n5157), .B1(n3084), .B2(n5518), .ZN(n3796)
         );
  INV_X1 U3893 ( .A(n3084), .ZN(n3802) );
  AOI211_X1 U3894 ( .C1(n3808), .C2(n3809), .A(n4796), .B(n4747), .ZN(n3084)
         );
  NOR2_X1 U3895 ( .A1(n5578), .A2(n5011), .ZN(n3809) );
  INV_X1 U3896 ( .A(n3810), .ZN(n3808) );
  AOI22_X1 U3897 ( .A1(n3811), .A2(n5157), .B1(n5156), .B2(n3812), .ZN(n3810)
         );
  AOI21_X1 U3898 ( .B1(n5522), .B2(n3813), .A(n5518), .ZN(n3811) );
  INV_X1 U3899 ( .A(n3798), .ZN(n3794) );
  AOI211_X1 U3900 ( .C1(n3814), .C2(n3806), .A(n5537), .B(n4748), .ZN(n3798)
         );
  NOR2_X1 U3901 ( .A1(n5570), .A2(n5572), .ZN(n3806) );
  OAI22_X1 U3902 ( .A1(n3815), .A2(n2932), .B1(n3792), .B2(n5159), .ZN(n3814)
         );
  OAI21_X1 U3903 ( .B1(n3793), .B2(n5161), .A(n2888), .ZN(n3815) );
  INV_X1 U3905 ( .A(n3742), .ZN(n3757) );
  AOI22_X1 U3906 ( .A1(n3816), .A2(n3073), .B1(n2910), .B2(n3817), .ZN(n3742)
         );
  INV_X1 U3907 ( .A(n2910), .ZN(n3073) );
  NAND2_X1 U3908 ( .A1(n3076), .A2(n2910), .ZN(n2997) );
  OAI21_X1 U3909 ( .B1(n2996), .B2(n3818), .A(n3819), .ZN(n2910) );
  OAI221_X1 U3910 ( .B1(n3820), .B2(n3756), .C1(n3821), .C2(n3746), .A(n3822), 
        .ZN(n3819) );
  OAI22_X1 U3911 ( .A1(n3823), .A2(n3755), .B1(n3824), .B2(n3816), .ZN(n3822)
         );
  OAI221_X1 U3912 ( .B1(n2933), .B2(n3080), .C1(n3825), .C2(n3079), .A(n3826), 
        .ZN(n3816) );
  NAND3_X1 U3913 ( .A1(n3079), .A2(n1896), .A3(n3827), .ZN(n3826) );
  INV_X1 U3914 ( .A(n3828), .ZN(n3825) );
  INV_X1 U3915 ( .A(n3817), .ZN(n3824) );
  OAI22_X1 U3916 ( .A1(n3829), .A2(n3821), .B1(n3830), .B2(n3076), .ZN(n3817)
         );
  INV_X1 U3917 ( .A(n3756), .ZN(n3823) );
  OAI22_X1 U3918 ( .A1(n3831), .A2(n3821), .B1(n3832), .B2(n3076), .ZN(n3756)
         );
  INV_X1 U3919 ( .A(n3076), .ZN(n3821) );
  INV_X1 U3920 ( .A(n3755), .ZN(n3820) );
  OAI222_X1 U3921 ( .A1(n3833), .A2(n3080), .B1(n3834), .B2(n3835), .C1(n3836), 
        .C2(n3079), .ZN(n3755) );
  NAND2_X1 U3922 ( .A1(n3079), .A2(n3835), .ZN(n3080) );
  INV_X1 U3923 ( .A(n3079), .ZN(n2996) );
  NAND3_X1 U3924 ( .A1(n3837), .A2(n3838), .A3(n3839), .ZN(n3079) );
  OAI21_X1 U3925 ( .B1(n5535), .B2(n5534), .A(n3840), .ZN(n3839) );
  NAND3_X1 U3926 ( .A1(n3818), .A2(n3836), .A3(n3841), .ZN(n3838) );
  NAND2_X1 U3927 ( .A1(n3842), .A2(n3835), .ZN(n3818) );
  OAI21_X1 U3928 ( .B1(n3841), .B2(n3836), .A(n3843), .ZN(n3837) );
  OAI22_X1 U3929 ( .A1(n3834), .A2(n3835), .B1(n3833), .B2(n3842), .ZN(n3843)
         );
  OAI22_X1 U3930 ( .A1(n5547), .A2(n3078), .B1(n5549), .B2(n3840), .ZN(n3836)
         );
  AOI221_X1 U3931 ( .B1(n4752), .B2(n3827), .C1(n2933), .C2(n3835), .A(n3828), 
        .ZN(n3841) );
  OAI22_X1 U3932 ( .A1(n3078), .A2(n2901), .B1(n3840), .B2(n2951), .ZN(n3828)
         );
  INV_X1 U3933 ( .A(n3078), .ZN(n3840) );
  AOI211_X1 U3934 ( .C1(n3844), .C2(n3845), .A(n5540), .B(n5005), .ZN(n3078)
         );
  NOR2_X1 U3935 ( .A1(n5535), .A2(n5534), .ZN(n3845) );
  OAI22_X1 U3936 ( .A1(n3846), .A2(n2901), .B1(n3719), .B2(n5549), .ZN(n3844)
         );
  OAI21_X1 U3939 ( .B1(n3847), .B2(n5547), .A(n2951), .ZN(n3846) );
  INV_X1 U3941 ( .A(n3835), .ZN(n3827) );
  OAI211_X1 U3942 ( .C1(n3848), .C2(n3842), .A(n3238), .B(n217), .ZN(n3835) );
  NAND2_X1 U3944 ( .A1(n220), .A2(n3107), .ZN(n3842) );
  AOI22_X1 U3947 ( .A1(n3849), .A2(n5552), .B1(n5553), .B2(n3834), .ZN(n3848)
         );
  AOI21_X1 U3949 ( .B1(n5551), .B2(n3833), .A(n1896), .ZN(n3849) );
  OAI21_X1 U3951 ( .B1(n3850), .B2(n3851), .A(n3852), .ZN(n3076) );
  OAI21_X1 U3952 ( .B1(n5533), .B2(n3010), .A(n3853), .ZN(n3852) );
  AOI22_X1 U3954 ( .A1(n3854), .A2(n3830), .B1(n3832), .B2(n3855), .ZN(n3851)
         );
  AOI22_X1 U3955 ( .A1(n3853), .A2(n5046), .B1(n3077), .B2(n5519), .ZN(n3830)
         );
  AOI21_X1 U3956 ( .B1(n3831), .B2(n3856), .A(n3829), .ZN(n3854) );
  AOI22_X1 U3957 ( .A1(n3072), .A2(n5009), .B1(n3857), .B2(n5053), .ZN(n3829)
         );
  INV_X1 U3958 ( .A(n3832), .ZN(n3856) );
  OAI22_X1 U3959 ( .A1(n5023), .A2(n3077), .B1(n5523), .B2(n3853), .ZN(n3832)
         );
  INV_X1 U3960 ( .A(n3853), .ZN(n3077) );
  NAND3_X1 U3961 ( .A1(n223), .A2(n3060), .A3(n3858), .ZN(n3853) );
  OAI211_X1 U3962 ( .C1(n3859), .C2(n3860), .A(n3861), .B(n4799), .ZN(n3858)
         );
  NOR2_X1 U3964 ( .A1(n5523), .A2(n3720), .ZN(n3860) );
  AOI211_X1 U3965 ( .C1(n5523), .C2(n3720), .A(n2902), .B(n5519), .ZN(n3859)
         );
  INV_X1 U3969 ( .A(n3855), .ZN(n3831) );
  OAI22_X1 U3970 ( .A1(n3857), .A2(n3862), .B1(n3863), .B2(n3072), .ZN(n3855)
         );
  INV_X1 U3971 ( .A(n3072), .ZN(n3857) );
  INV_X1 U3972 ( .A(n3746), .ZN(n3850) );
  OAI21_X1 U3973 ( .B1(n5530), .B2(n4797), .A(n3072), .ZN(n3746) );
  OAI211_X1 U3974 ( .C1(n3864), .C2(n3865), .A(n2953), .B(n228), .ZN(n3072) );
  OR2_X1 U3977 ( .A1(n5530), .A2(n4797), .ZN(n3865) );
  AOI22_X1 U3978 ( .A1(n3866), .A2(n5009), .B1(n5010), .B2(n3863), .ZN(n3864)
         );
  AOI21_X1 U3979 ( .B1(n5008), .B2(n3862), .A(n5053), .ZN(n3866) );
  AOI22_X1 U3980 ( .A1(n2913), .A2(n3786), .B1(n2915), .B2(n3785), .ZN(n3621)
         );
  INV_X1 U3983 ( .A(n3011), .ZN(n2913) );
  NAND2_X1 U3985 ( .A1(n3214), .A2(n3538), .ZN(n2723) );
  INV_X1 U3986 ( .A(n3243), .ZN(n3214) );
  NAND2_X1 U3987 ( .A1(n2340), .A2(n3213), .ZN(n3243) );
  INV_X1 U3988 ( .A(n2390), .ZN(n2340) );
  NAND3_X1 U3989 ( .A1(n3867), .A2(n1774), .A3(n1773), .ZN(n2390) );
  INV_X1 U3990 ( .A(n1780), .ZN(n1773) );
  NAND2_X1 U3991 ( .A1(n3868), .A2(n3869), .ZN(n2062) );
  AOI221_X1 U3992 ( .B1(n2915), .B2(n231), .C1(hrdata_i[7]), .C2(n2879), .A(
        n3870), .ZN(n3869) );
  OAI22_X1 U3993 ( .A1(n5530), .A2(n3011), .B1(n3871), .B2(n2926), .ZN(n3870)
         );
  AOI221_X1 U3994 ( .B1(n1887), .B2(n3784), .C1(n1890), .C2(n3812), .A(n3872), 
        .ZN(n3871) );
  OAI22_X1 U3995 ( .A1(n5523), .A2(n2886), .B1(n5549), .B2(n2885), .ZN(n3872)
         );
  INV_X1 U3999 ( .A(n2948), .ZN(n2915) );
  NOR4_X1 U4001 ( .A1(n3874), .A2(n3875), .A3(n1110), .A4(n5502), .ZN(n252) );
  INV_X1 U4002 ( .A(n3876), .ZN(n3868) );
  OAI222_X1 U4003 ( .A1(n298), .A2(n2981), .B1(n1789), .B2(n2998), .C1(n16685), 
        .C2(n5520), .ZN(n3876) );
  OAI22_X1 U4004 ( .A1(n2337), .A2(n2386), .B1(n16788), .B2(n2338), .ZN(n1789)
         );
  OAI221_X1 U4005 ( .B1(n3329), .B2(n16950), .C1(n3314), .C2(n16953), .A(n3877), .ZN(n2338) );
  AOI22_X1 U4006 ( .A1(n16947), .A2(n3317), .B1(n16942), .B2(n3155), .ZN(n3877) );
  NAND3_X1 U4007 ( .A1(n3878), .A2(n3879), .A3(n3880), .ZN(n3155) );
  AOI221_X1 U4008 ( .B1(n16941), .B2(vis_r2_o[10]), .C1(n16938), .C2(
        vis_r0_o[10]), .A(n3883), .ZN(n3880) );
  OAI22_X1 U4009 ( .A1(n5146), .A2(n16935), .B1(n5445), .B2(n16932), .ZN(n3883) );
  AOI22_X1 U4011 ( .A1(n16929), .A2(vis_r5_o[10]), .B1(n16926), .B2(
        vis_r4_o[10]), .ZN(n3879) );
  AOI22_X1 U4012 ( .A1(n16923), .A2(vis_r6_o[10]), .B1(n16920), .B2(
        vis_r1_o[10]), .ZN(n3878) );
  NAND3_X1 U4015 ( .A1(n3888), .A2(n3889), .A3(n3890), .ZN(n3317) );
  AOI221_X1 U4016 ( .B1(n16941), .B2(vis_r2_o[8]), .C1(n16938), .C2(
        vis_r0_o[8]), .A(n3893), .ZN(n3890) );
  OAI22_X1 U4017 ( .A1(n5137), .A2(n16935), .B1(n5448), .B2(n16932), .ZN(n3893) );
  AOI22_X1 U4019 ( .A1(n16929), .A2(vis_r5_o[8]), .B1(n16926), .B2(vis_r4_o[8]), .ZN(n3889) );
  AOI22_X1 U4020 ( .A1(n16923), .A2(vis_r6_o[8]), .B1(n16920), .B2(vis_r1_o[8]), .ZN(n3888) );
  INV_X1 U4023 ( .A(n2209), .ZN(n3314) );
  NAND3_X1 U4024 ( .A1(n3898), .A2(n3899), .A3(n3900), .ZN(n2209) );
  AOI221_X1 U4025 ( .B1(n16940), .B2(vis_r2_o[7]), .C1(n16937), .C2(
        vis_r0_o[7]), .A(n3903), .ZN(n3900) );
  OAI22_X1 U4026 ( .A1(n5020), .A2(n16934), .B1(n5423), .B2(n16931), .ZN(n3903) );
  AOI22_X1 U4029 ( .A1(n16928), .A2(vis_r5_o[7]), .B1(n16925), .B2(vis_r4_o[7]), .ZN(n3899) );
  AOI22_X1 U4030 ( .A1(n16922), .A2(vis_r6_o[7]), .B1(n16919), .B2(vis_r1_o[7]), .ZN(n3898) );
  INV_X1 U4033 ( .A(n3237), .ZN(n3329) );
  NAND3_X1 U4034 ( .A1(n3908), .A2(n3909), .A3(n3910), .ZN(n3237) );
  AOI221_X1 U4035 ( .B1(n16940), .B2(vis_r2_o[9]), .C1(n16937), .C2(
        vis_r0_o[9]), .A(n3913), .ZN(n3910) );
  OAI22_X1 U4036 ( .A1(n5143), .A2(n16934), .B1(n5447), .B2(n16931), .ZN(n3913) );
  AOI22_X1 U4038 ( .A1(n16928), .A2(vis_r5_o[9]), .B1(n16925), .B2(vis_r4_o[9]), .ZN(n3909) );
  AOI22_X1 U4039 ( .A1(n16922), .A2(vis_r6_o[9]), .B1(n16919), .B2(vis_r1_o[9]), .ZN(n3908) );
  OAI221_X1 U4042 ( .B1(n3265), .B2(n3279), .C1(n3328), .C2(n16953), .A(n3918), 
        .ZN(n2386) );
  AOI22_X1 U4043 ( .A1(n16947), .A2(n3041), .B1(n3275), .B2(n3022), .ZN(n3918)
         );
  NAND3_X1 U4044 ( .A1(n3919), .A2(n3920), .A3(n3921), .ZN(n3022) );
  AOI221_X1 U4045 ( .B1(n16940), .B2(vis_r2_o[13]), .C1(n16937), .C2(
        vis_r0_o[13]), .A(n3924), .ZN(n3921) );
  OAI22_X1 U4046 ( .A1(n5134), .A2(n16934), .B1(n5443), .B2(n16931), .ZN(n3924) );
  AOI22_X1 U4048 ( .A1(n16928), .A2(vis_r5_o[13]), .B1(n16925), .B2(
        vis_r4_o[13]), .ZN(n3920) );
  AOI22_X1 U4049 ( .A1(n16922), .A2(vis_r6_o[13]), .B1(n16919), .B2(
        vis_r1_o[13]), .ZN(n3919) );
  NAND3_X1 U4052 ( .A1(n3929), .A2(n3930), .A3(n3931), .ZN(n3041) );
  AOI221_X1 U4053 ( .B1(n16940), .B2(vis_r2_o[12]), .C1(n16937), .C2(
        vis_r0_o[12]), .A(n3934), .ZN(n3931) );
  OAI22_X1 U4054 ( .A1(n5129), .A2(n16934), .B1(n5444), .B2(n16931), .ZN(n3934) );
  AOI22_X1 U4056 ( .A1(n16928), .A2(vis_r5_o[12]), .B1(n16925), .B2(
        vis_r4_o[12]), .ZN(n3930) );
  AOI22_X1 U4057 ( .A1(n16922), .A2(vis_r6_o[12]), .B1(n16919), .B2(
        vis_r1_o[12]), .ZN(n3929) );
  INV_X1 U4060 ( .A(n3134), .ZN(n3328) );
  NAND3_X1 U4061 ( .A1(n3939), .A2(n3940), .A3(n3941), .ZN(n3134) );
  AOI221_X1 U4062 ( .B1(n16940), .B2(vis_r2_o[11]), .C1(n16937), .C2(
        vis_r0_o[11]), .A(n3944), .ZN(n3941) );
  OAI22_X1 U4063 ( .A1(n5565), .A2(n16934), .B1(n5557), .B2(n16931), .ZN(n3944) );
  AOI22_X1 U4065 ( .A1(n16928), .A2(vis_r5_o[11]), .B1(n16925), .B2(
        vis_r4_o[11]), .ZN(n3940) );
  AOI22_X1 U4066 ( .A1(n16922), .A2(vis_r6_o[11]), .B1(n16919), .B2(
        vis_r1_o[11]), .ZN(n3939) );
  INV_X1 U4069 ( .A(n2964), .ZN(n3265) );
  NAND3_X1 U4070 ( .A1(n3949), .A2(n3950), .A3(n3951), .ZN(n2964) );
  AOI221_X1 U4071 ( .B1(n16940), .B2(vis_r2_o[14]), .C1(n16937), .C2(
        vis_r0_o[14]), .A(n3954), .ZN(n3951) );
  OAI22_X1 U4072 ( .A1(n5105), .A2(n16934), .B1(n5442), .B2(n16931), .ZN(n3954) );
  AOI22_X1 U4074 ( .A1(n16928), .A2(vis_r5_o[14]), .B1(n16925), .B2(
        vis_r4_o[14]), .ZN(n3950) );
  AOI22_X1 U4075 ( .A1(n16922), .A2(vis_r6_o[14]), .B1(n16919), .B2(
        vis_r1_o[14]), .ZN(n3949) );
  OAI21_X1 U4078 ( .B1(n2389), .B2(n3475), .A(n3285), .ZN(n2069) );
  NAND2_X1 U4079 ( .A1(n3215), .A2(n1574), .ZN(n3285) );
  NAND2_X1 U4080 ( .A1(n2358), .A2(n3213), .ZN(n3475) );
  INV_X1 U4081 ( .A(n3539), .ZN(n2358) );
  NAND3_X1 U4082 ( .A1(n1780), .A2(n3867), .A3(n1790), .ZN(n3539) );
  OAI21_X1 U4083 ( .B1(n3215), .B2(n3477), .A(n3476), .ZN(n2072) );
  OAI21_X1 U4084 ( .B1(n16869), .B2(n3959), .A(n3215), .ZN(n3476) );
  AOI21_X1 U4085 ( .B1(n16826), .B2(n16842), .A(n760), .ZN(n3959) );
  NAND3_X1 U4086 ( .A1(n3867), .A2(n1774), .A3(n1780), .ZN(n3477) );
  OAI211_X1 U4088 ( .C1(n2998), .C2(n2375), .A(n2919), .B(n3960), .ZN(n2057)
         );
  AOI222_X1 U4089 ( .A1(hrdata_i[31]), .A2(n2879), .B1(n2882), .B2(n3961), 
        .C1(n2895), .C2(n1066), .ZN(n3960) );
  NAND2_X1 U4092 ( .A1(n3963), .A2(n3964), .ZN(n3961) );
  AOI222_X1 U4093 ( .A1(n1887), .A2(n3791), .B1(n3965), .B2(n1189), .C1(n1191), 
        .C2(n3740), .ZN(n3964) );
  NOR2_X1 U4095 ( .A1(n5504), .A2(n2930), .ZN(n3965) );
  AOI222_X1 U4096 ( .A1(n1893), .A2(n3862), .B1(n1890), .B2(n3792), .C1(n1897), 
        .C2(n3833), .ZN(n3963) );
  INV_X1 U4097 ( .A(n2885), .ZN(n1897) );
  INV_X1 U4098 ( .A(n2886), .ZN(n1893) );
  AND2_X1 U4099 ( .A1(n3003), .A2(n3966), .ZN(n2919) );
  NAND3_X1 U4100 ( .A1(n3318), .A2(n5502), .A3(n3967), .ZN(n3966) );
  NOR3_X1 U4101 ( .A1(n5096), .A2(n4905), .A3(n5017), .ZN(n3967) );
  NOR2_X1 U4102 ( .A1(n2926), .A2(n5149), .ZN(n3318) );
  NAND2_X1 U4103 ( .A1(n2882), .A2(n14), .ZN(n3003) );
  NOR3_X1 U4104 ( .A1(n2930), .A2(n5502), .A3(n3875), .ZN(n14) );
  OAI22_X1 U4105 ( .A1(n2313), .A2(n3968), .B1(n1786), .B2(n3969), .ZN(n2375)
         );
  INV_X1 U4106 ( .A(n3968), .ZN(n3969) );
  INV_X1 U4107 ( .A(n3970), .ZN(n1786) );
  OAI22_X1 U4108 ( .A1(n16789), .A2(n2369), .B1(n2337), .B2(n2334), .ZN(n3970)
         );
  OAI221_X1 U4109 ( .B1(n3315), .B2(n16950), .C1(n3319), .C2(n16953), .A(n3971), .ZN(n2334) );
  AOI22_X1 U4110 ( .A1(n16947), .A2(n2585), .B1(n16942), .B2(n2531), .ZN(n3971) );
  NAND3_X1 U4111 ( .A1(n3972), .A2(n3973), .A3(n3974), .ZN(n2531) );
  AOI221_X1 U4112 ( .B1(n16940), .B2(vis_r2_o[6]), .C1(n16937), .C2(
        vis_r0_o[6]), .A(n3977), .ZN(n3974) );
  OAI22_X1 U4113 ( .A1(n5043), .A2(n16934), .B1(n5432), .B2(n16931), .ZN(n3977) );
  AOI22_X1 U4116 ( .A1(n16928), .A2(vis_r5_o[6]), .B1(n16925), .B2(vis_r4_o[6]), .ZN(n3973) );
  AOI22_X1 U4117 ( .A1(n16922), .A2(vis_r6_o[6]), .B1(n16919), .B2(vis_r1_o[6]), .ZN(n3972) );
  NAND3_X1 U4120 ( .A1(n3982), .A2(n3983), .A3(n3984), .ZN(n2585) );
  AOI221_X1 U4121 ( .B1(n16940), .B2(vis_r2_o[4]), .C1(n16937), .C2(
        vis_r0_o[4]), .A(n3987), .ZN(n3984) );
  OAI22_X1 U4122 ( .A1(n5123), .A2(n16934), .B1(n5434), .B2(n16931), .ZN(n3987) );
  AOI22_X1 U4125 ( .A1(n16928), .A2(vis_r5_o[4]), .B1(n16925), .B2(vis_r4_o[4]), .ZN(n3983) );
  AOI22_X1 U4126 ( .A1(n16922), .A2(vis_r6_o[4]), .B1(n16919), .B2(vis_r1_o[4]), .ZN(n3982) );
  INV_X1 U4129 ( .A(n2612), .ZN(n3319) );
  NAND3_X1 U4130 ( .A1(n3992), .A2(n3993), .A3(n3994), .ZN(n2612) );
  AOI221_X1 U4131 ( .B1(n16940), .B2(vis_r2_o[3]), .C1(n16937), .C2(
        vis_r0_o[3]), .A(n3997), .ZN(n3994) );
  OAI22_X1 U4132 ( .A1(n5030), .A2(n16934), .B1(n5435), .B2(n16931), .ZN(n3997) );
  AOI22_X1 U4135 ( .A1(n16928), .A2(vis_r5_o[3]), .B1(n16925), .B2(vis_r4_o[3]), .ZN(n3993) );
  AOI22_X1 U4136 ( .A1(n16922), .A2(vis_r6_o[3]), .B1(n16919), .B2(vis_r1_o[3]), .ZN(n3992) );
  INV_X1 U4139 ( .A(n2562), .ZN(n3315) );
  NAND3_X1 U4140 ( .A1(n4002), .A2(n4003), .A3(n4004), .ZN(n2562) );
  AOI221_X1 U4141 ( .B1(n16940), .B2(vis_r2_o[5]), .C1(n16937), .C2(
        vis_r0_o[5]), .A(n4007), .ZN(n4004) );
  OAI22_X1 U4142 ( .A1(n5093), .A2(n16934), .B1(n5433), .B2(n16931), .ZN(n4007) );
  AOI22_X1 U4145 ( .A1(n16928), .A2(vis_r5_o[5]), .B1(n16925), .B2(vis_r4_o[5]), .ZN(n4003) );
  AOI22_X1 U4146 ( .A1(n16922), .A2(vis_r6_o[5]), .B1(n16919), .B2(vis_r1_o[5]), .ZN(n4002) );
  OAI221_X1 U4149 ( .B1(n3280), .B2(n16950), .C1(n3278), .C2(n16953), .A(n4012), .ZN(n2369) );
  AOI22_X1 U4150 ( .A1(n16947), .A2(n3274), .B1(n16942), .B2(n3199), .ZN(n4012) );
  NAND3_X1 U4151 ( .A1(n4013), .A2(n4014), .A3(n4015), .ZN(n3199) );
  AOI221_X1 U4152 ( .B1(n16940), .B2(vis_r2_o[2]), .C1(n16937), .C2(
        vis_r0_o[2]), .A(n4018), .ZN(n4015) );
  OAI22_X1 U4153 ( .A1(n5058), .A2(n16934), .B1(n5446), .B2(n16931), .ZN(n4018) );
  AOI22_X1 U4156 ( .A1(n16928), .A2(vis_r5_o[2]), .B1(n16925), .B2(vis_r4_o[2]), .ZN(n4014) );
  AOI22_X1 U4157 ( .A1(n16922), .A2(vis_r6_o[2]), .B1(n16919), .B2(vis_r1_o[2]), .ZN(n4013) );
  NAND3_X1 U4160 ( .A1(n4023), .A2(n4024), .A3(n4025), .ZN(n3274) );
  AOI221_X1 U4161 ( .B1(n16939), .B2(vis_r2_o[0]), .C1(n16936), .C2(
        vis_r0_o[0]), .A(n4028), .ZN(n4025) );
  OAI22_X1 U4162 ( .A1(n5038), .A2(n16933), .B1(n5425), .B2(n16930), .ZN(n4028) );
  AOI22_X1 U4165 ( .A1(n16927), .A2(vis_r5_o[0]), .B1(n16924), .B2(vis_r4_o[0]), .ZN(n4024) );
  AOI22_X1 U4166 ( .A1(n16921), .A2(vis_r6_o[0]), .B1(n16918), .B2(vis_r1_o[0]), .ZN(n4023) );
  INV_X1 U4169 ( .A(n3400), .ZN(n3278) );
  INV_X1 U4170 ( .A(n2639), .ZN(n3280) );
  NAND3_X1 U4171 ( .A1(n4033), .A2(n4034), .A3(n4035), .ZN(n2639) );
  AOI221_X1 U4172 ( .B1(n16939), .B2(vis_r2_o[1]), .C1(n16936), .C2(
        vis_r0_o[1]), .A(n4038), .ZN(n4035) );
  OAI22_X1 U4173 ( .A1(n4985), .A2(n16933), .B1(n5424), .B2(n16930), .ZN(n4038) );
  AOI22_X1 U4176 ( .A1(n16927), .A2(vis_r5_o[1]), .B1(n16924), .B2(vis_r4_o[1]), .ZN(n4034) );
  AOI22_X1 U4177 ( .A1(n16921), .A2(vis_r6_o[1]), .B1(n16918), .B2(vis_r1_o[1]), .ZN(n4033) );
  AOI22_X1 U4180 ( .A1(n3118), .A2(n2940), .B1(n16951), .B2(n2941), .ZN(n3968)
         );
  NOR2_X1 U4181 ( .A1(n3120), .A2(n16851), .ZN(n2941) );
  INV_X1 U4182 ( .A(n3091), .ZN(n2940) );
  OAI211_X1 U4183 ( .C1(n3120), .C2(n16789), .A(n3119), .B(n16848), .ZN(n3091)
         );
  NAND2_X1 U4184 ( .A1(n3120), .A2(n16789), .ZN(n3119) );
  INV_X1 U4185 ( .A(n3343), .ZN(n3120) );
  NAND2_X1 U4186 ( .A1(n3538), .A2(n3478), .ZN(n3343) );
  NAND4_X1 U4187 ( .A1(n3118), .A2(n2337), .A3(n1780), .A4(n1774), .ZN(n3478)
         );
  INV_X1 U4188 ( .A(n3092), .ZN(n2313) );
  NAND3_X1 U4189 ( .A1(n3400), .A2(n1759), .A3(n4043), .ZN(n3092) );
  OAI21_X1 U4190 ( .B1(n16830), .B2(n1086), .A(n1784), .ZN(n4043) );
  NAND3_X1 U4191 ( .A1(n4044), .A2(n4045), .A3(n4046), .ZN(n3400) );
  AOI221_X1 U4192 ( .B1(n16939), .B2(vis_r2_o[31]), .C1(n16936), .C2(
        vis_r0_o[31]), .A(n4049), .ZN(n4046) );
  OAI22_X1 U4193 ( .A1(n4962), .A2(n16933), .B1(n5421), .B2(n16930), .ZN(n4049) );
  AOI22_X1 U4195 ( .A1(n16927), .A2(vis_r5_o[31]), .B1(n16924), .B2(
        vis_r4_o[31]), .ZN(n4045) );
  AOI22_X1 U4196 ( .A1(n16921), .A2(vis_r6_o[31]), .B1(n16918), .B2(
        vis_r1_o[31]), .ZN(n4044) );
  OAI21_X1 U4199 ( .B1(n3213), .B2(n1027), .A(n3472), .ZN(n2067) );
  NAND2_X1 U4200 ( .A1(n2322), .A2(n3213), .ZN(n3472) );
  NOR2_X1 U4201 ( .A1(n3217), .A2(n2389), .ZN(n2322) );
  INV_X1 U4202 ( .A(n3538), .ZN(n2389) );
  NAND2_X1 U4203 ( .A1(n16834), .A2(n918), .ZN(n3538) );
  NAND2_X1 U4205 ( .A1(n1793), .A2(n16849), .ZN(n3867) );
  OAI21_X1 U4206 ( .B1(n4054), .B2(n1519), .A(n4055), .ZN(n1793) );
  NAND4_X1 U4207 ( .A1(n563), .A2(n16833), .A3(n4056), .A4(n4057), .ZN(n4055)
         );
  NOR3_X1 U4208 ( .A1(n16656), .A2(n16671), .A3(n795), .ZN(n4057) );
  INV_X1 U4209 ( .A(n3566), .ZN(n4056) );
  NOR3_X1 U4211 ( .A1(n1794), .A2(n4058), .A3(n1795), .ZN(n4054) );
  NOR2_X1 U4212 ( .A1(n1774), .A2(n1780), .ZN(n1777) );
  OAI21_X1 U4213 ( .B1(n16830), .B2(n4059), .A(n4060), .ZN(n1780) );
  OAI21_X1 U4214 ( .B1(n4061), .B2(n1763), .A(n16831), .ZN(n4060) );
  AND3_X1 U4215 ( .A1(n4062), .A2(n4063), .A3(n4064), .ZN(n1763) );
  AOI21_X1 U4216 ( .B1(n4062), .B2(n4063), .A(n4064), .ZN(n4061) );
  INV_X1 U4217 ( .A(n4064), .ZN(n4059) );
  AOI22_X1 U4218 ( .A1(n16671), .A2(n563), .B1(n4065), .B2(n529), .ZN(n4064)
         );
  INV_X1 U4219 ( .A(n1790), .ZN(n1774) );
  AOI22_X1 U4220 ( .A1(n16833), .A2(n4063), .B1(n16828), .B2(n4066), .ZN(n1790) );
  XNOR2_X1 U4221 ( .A(n4063), .B(n4062), .ZN(n4066) );
  AND2_X1 U4222 ( .A1(n4067), .A2(n4068), .ZN(n4062) );
  AOI22_X1 U4223 ( .A1(n795), .A2(n563), .B1(n4069), .B2(n529), .ZN(n4063) );
  NAND2_X1 U4225 ( .A1(n195), .A2(n16842), .ZN(n1027) );
  NAND2_X1 U4227 ( .A1(n624), .A2(n616), .ZN(n4070) );
  OAI221_X1 U4228 ( .B1(n16685), .B2(n262), .C1(n2981), .C2(n264), .A(n4071), 
        .ZN(n2061) );
  AOI222_X1 U4229 ( .A1(n1787), .A2(n2922), .B1(n2882), .B2(n4072), .C1(
        hrdata_i[23]), .C2(n2879), .ZN(n4071) );
  AND3_X1 U4232 ( .A1(n4905), .A2(n5096), .A3(n1189), .ZN(n1111) );
  NOR2_X1 U4233 ( .A1(n4073), .A2(n3875), .ZN(n1189) );
  OAI221_X1 U4234 ( .B1(n5551), .B2(n2885), .C1(n5008), .C2(n2886), .A(n4074), 
        .ZN(n4072) );
  AOI222_X1 U4235 ( .A1(n1890), .A2(n3793), .B1(n1191), .B2(n3731), .C1(n1887), 
        .C2(n3790), .ZN(n4074) );
  INV_X1 U4237 ( .A(n2898), .ZN(n1887) );
  NAND3_X1 U4238 ( .A1(n4073), .A2(n3875), .A3(n1188), .ZN(n2898) );
  INV_X1 U4239 ( .A(n2930), .ZN(n1188) );
  NAND3_X1 U4240 ( .A1(n3874), .A2(n251), .A3(n5149), .ZN(n2930) );
  AND3_X1 U4242 ( .A1(n5017), .A2(n4073), .A3(n4075), .ZN(n1191) );
  INV_X1 U4244 ( .A(n2899), .ZN(n1890) );
  NAND3_X1 U4245 ( .A1(n4905), .A2(n5149), .A3(n4076), .ZN(n2899) );
  NOR3_X1 U4246 ( .A1(n5502), .A2(n5017), .A3(n5096), .ZN(n4076) );
  NAND3_X1 U4247 ( .A1(n3875), .A2(n251), .A3(n3717), .ZN(n2886) );
  NAND3_X1 U4248 ( .A1(n3717), .A2(n3875), .A3(n4905), .ZN(n2885) );
  OAI211_X1 U4251 ( .C1(n16845), .C2(n526), .A(n1233), .B(n3546), .ZN(n4077)
         );
  NAND2_X1 U4252 ( .A1(n16806), .A2(n16866), .ZN(n3546) );
  INV_X1 U4253 ( .A(n2346), .ZN(n1787) );
  OAI22_X1 U4254 ( .A1(n16789), .A2(n2356), .B1(n2337), .B2(n3117), .ZN(n2346)
         );
  OAI221_X1 U4255 ( .B1(n3341), .B2(n16950), .C1(n3338), .C2(n16953), .A(n4078), .ZN(n3117) );
  AOI22_X1 U4256 ( .A1(n16947), .A2(n2271), .B1(n16942), .B2(n2297), .ZN(n4078) );
  NAND3_X1 U4257 ( .A1(n4079), .A2(n4080), .A3(n4081), .ZN(n2297) );
  AOI221_X1 U4258 ( .B1(n16939), .B2(vis_r2_o[30]), .C1(n16936), .C2(
        vis_r0_o[30]), .A(n4084), .ZN(n4081) );
  OAI22_X1 U4259 ( .A1(n5082), .A2(n16933), .B1(n5426), .B2(n16930), .ZN(n4084) );
  AOI22_X1 U4261 ( .A1(n16927), .A2(vis_r5_o[30]), .B1(n16924), .B2(
        vis_r4_o[30]), .ZN(n4080) );
  AOI22_X1 U4262 ( .A1(n16921), .A2(vis_r6_o[30]), .B1(n16918), .B2(
        vis_r1_o[30]), .ZN(n4079) );
  NAND3_X1 U4265 ( .A1(n4089), .A2(n4090), .A3(n4091), .ZN(n2271) );
  AOI221_X1 U4266 ( .B1(n16939), .B2(vis_r2_o[28]), .C1(n16936), .C2(
        vis_r0_o[28]), .A(n4094), .ZN(n4091) );
  OAI22_X1 U4267 ( .A1(n4996), .A2(n16933), .B1(n5422), .B2(n16930), .ZN(n4094) );
  AOI22_X1 U4269 ( .A1(n16927), .A2(vis_r5_o[28]), .B1(n16924), .B2(
        vis_r4_o[28]), .ZN(n4090) );
  AOI22_X1 U4270 ( .A1(n16921), .A2(vis_r6_o[28]), .B1(n16918), .B2(
        vis_r1_o[28]), .ZN(n4089) );
  INV_X1 U4273 ( .A(n2433), .ZN(n3338) );
  NAND3_X1 U4274 ( .A1(n4099), .A2(n4100), .A3(n4101), .ZN(n2433) );
  AOI221_X1 U4275 ( .B1(n16939), .B2(vis_r2_o[27]), .C1(n16936), .C2(
        vis_r0_o[27]), .A(n4104), .ZN(n4101) );
  OAI22_X1 U4276 ( .A1(n5113), .A2(n16933), .B1(n5428), .B2(n16930), .ZN(n4104) );
  AOI22_X1 U4278 ( .A1(n16927), .A2(vis_r5_o[27]), .B1(n16924), .B2(
        vis_r4_o[27]), .ZN(n4100) );
  AOI22_X1 U4279 ( .A1(n16921), .A2(vis_r6_o[27]), .B1(n16918), .B2(
        vis_r1_o[27]), .ZN(n4099) );
  INV_X1 U4282 ( .A(n2402), .ZN(n3341) );
  NAND3_X1 U4283 ( .A1(n4109), .A2(n4110), .A3(n4111), .ZN(n2402) );
  AOI221_X1 U4284 ( .B1(n16939), .B2(vis_r2_o[29]), .C1(n16936), .C2(
        vis_r0_o[29]), .A(n4114), .ZN(n4111) );
  OAI22_X1 U4285 ( .A1(n5077), .A2(n16933), .B1(n5427), .B2(n16930), .ZN(n4114) );
  AOI22_X1 U4287 ( .A1(n16927), .A2(vis_r5_o[29]), .B1(n16924), .B2(
        vis_r4_o[29]), .ZN(n4110) );
  AOI22_X1 U4288 ( .A1(n16921), .A2(vis_r6_o[29]), .B1(n16918), .B2(
        vis_r1_o[29]), .ZN(n4109) );
  OAI221_X1 U4292 ( .B1(n3339), .B2(n16948), .C1(n3345), .C2(n16951), .A(n4119), .ZN(n2356) );
  AOI22_X1 U4293 ( .A1(n16945), .A2(n2507), .B1(n16942), .B2(n2452), .ZN(n4119) );
  NAND3_X1 U4294 ( .A1(n4120), .A2(n4121), .A3(n4122), .ZN(n2452) );
  AOI221_X1 U4295 ( .B1(n16939), .B2(vis_r2_o[26]), .C1(n16936), .C2(
        vis_r0_o[26]), .A(n4125), .ZN(n4122) );
  OAI22_X1 U4296 ( .A1(n4991), .A2(n16933), .B1(n5429), .B2(n16930), .ZN(n4125) );
  AOI22_X1 U4298 ( .A1(n16927), .A2(vis_r5_o[26]), .B1(n16924), .B2(
        vis_r4_o[26]), .ZN(n4121) );
  AOI22_X1 U4299 ( .A1(n16921), .A2(vis_r6_o[26]), .B1(n16918), .B2(
        vis_r1_o[26]), .ZN(n4120) );
  NAND2_X1 U4303 ( .A1(n4130), .A2(n4131), .ZN(n3279) );
  NAND3_X1 U4304 ( .A1(n4132), .A2(n4133), .A3(n4134), .ZN(n2507) );
  AOI221_X1 U4305 ( .B1(n16939), .B2(vis_r2_o[24]), .C1(n16936), .C2(
        vis_r0_o[24]), .A(n4137), .ZN(n4134) );
  OAI22_X1 U4306 ( .A1(n4972), .A2(n16933), .B1(n5431), .B2(n16930), .ZN(n4137) );
  AOI22_X1 U4308 ( .A1(n16927), .A2(vis_r5_o[24]), .B1(n16924), .B2(
        vis_r4_o[24]), .ZN(n4133) );
  AOI22_X1 U4309 ( .A1(n16921), .A2(vis_r6_o[24]), .B1(n16918), .B2(
        vis_r1_o[24]), .ZN(n4132) );
  NAND2_X1 U4313 ( .A1(n4131), .A2(n4142), .ZN(n3277) );
  INV_X1 U4316 ( .A(n3254), .ZN(n3345) );
  NAND3_X1 U4317 ( .A1(n4143), .A2(n4144), .A3(n4145), .ZN(n3254) );
  AOI221_X1 U4318 ( .B1(n16939), .B2(vis_r2_o[23]), .C1(n16936), .C2(
        vis_r0_o[23]), .A(n4148), .ZN(n4145) );
  OAI22_X1 U4319 ( .A1(n4960), .A2(n16933), .B1(n5585), .B2(n16930), .ZN(n4148) );
  AOI22_X1 U4321 ( .A1(n16927), .A2(vis_r5_o[23]), .B1(n16924), .B2(
        vis_r4_o[23]), .ZN(n4144) );
  AOI22_X1 U4322 ( .A1(n16921), .A2(vis_r6_o[23]), .B1(n16918), .B2(
        vis_r1_o[23]), .ZN(n4143) );
  INV_X1 U4327 ( .A(n4130), .ZN(n4142) );
  AOI221_X1 U4328 ( .B1(n4153), .B2(n4154), .C1(n16833), .C2(n4155), .A(n4067), 
        .ZN(n4130) );
  INV_X1 U4329 ( .A(n4153), .ZN(n4155) );
  AND2_X1 U4330 ( .A1(n4131), .A2(n16830), .ZN(n4154) );
  INV_X1 U4331 ( .A(n2484), .ZN(n3339) );
  NAND3_X1 U4332 ( .A1(n4156), .A2(n4157), .A3(n4158), .ZN(n2484) );
  AOI221_X1 U4333 ( .B1(n16939), .B2(vis_r2_o[25]), .C1(n16936), .C2(
        vis_r0_o[25]), .A(n4161), .ZN(n4158) );
  OAI22_X1 U4334 ( .A1(n5014), .A2(n16933), .B1(n5430), .B2(n16930), .ZN(n4161) );
  NOR3_X1 U4337 ( .A1(n5036), .A2(n4978), .A3(n3495), .ZN(n4162) );
  NOR3_X1 U4341 ( .A1(n3488), .A2(n3495), .A3(n3492), .ZN(n4163) );
  AOI22_X1 U4342 ( .A1(n16927), .A2(vis_r5_o[25]), .B1(n16924), .B2(
        vis_r4_o[25]), .ZN(n4157) );
  AOI22_X1 U4346 ( .A1(n16921), .A2(vis_r6_o[25]), .B1(n16918), .B2(
        vis_r1_o[25]), .ZN(n4156) );
  NOR2_X1 U4349 ( .A1(n3480), .A2(n4978), .ZN(n3592) );
  NOR2_X1 U4356 ( .A1(n4067), .A2(n16833), .ZN(n4168) );
  NOR2_X1 U4357 ( .A1(n4131), .A2(n4153), .ZN(n4067) );
  OAI22_X1 U4358 ( .A1(n5027), .A2(n1234), .B1(n4169), .B2(n1519), .ZN(n4153)
         );
  OAI22_X1 U4359 ( .A1(n5120), .A2(n1234), .B1(n4170), .B2(n1519), .ZN(n4131)
         );
  AOI22_X1 U4360 ( .A1(n16656), .A2(n563), .B1(n4171), .B2(n529), .ZN(n4068)
         );
  NAND2_X1 U4361 ( .A1(n316), .A2(n2882), .ZN(n2981) );
  AND3_X1 U4363 ( .A1(n5502), .A2(n3875), .A3(n4075), .ZN(n316) );
  NOR3_X1 U4364 ( .A1(n5149), .A2(n5096), .A3(n251), .ZN(n4075) );
  NAND4_X1 U4368 ( .A1(n5502), .A2(n5096), .A3(n5149), .A4(n3875), .ZN(n261)
         );
  OAI211_X1 U4371 ( .C1(n16845), .C2(n1964), .A(n4173), .B(n4174), .ZN(n4172)
         );
  AOI21_X1 U4372 ( .B1(n1262), .B2(n16869), .A(n17096), .ZN(n4174) );
  INV_X1 U4373 ( .A(n616), .ZN(n1262) );
  NAND3_X1 U4375 ( .A1(n16845), .A2(n16864), .A3(n757), .ZN(n4173) );
  INV_X1 U4376 ( .A(n624), .ZN(n757) );
  NAND2_X1 U4377 ( .A1(n16680), .A2(n16871), .ZN(n624) );
  NAND2_X1 U4378 ( .A1(n526), .A2(n16838), .ZN(n1964) );
  AOI21_X1 U4380 ( .B1(n84), .B2(n1508), .A(n17127), .ZN(n2085) );
  AOI21_X1 U4382 ( .B1(n4175), .B2(n16871), .A(n3516), .ZN(n1508) );
  NOR2_X1 U4383 ( .A1(n758), .A2(n1519), .ZN(n3516) );
  OR4_X1 U4384 ( .A1(n1801), .A2(n1803), .A3(n4176), .A4(n4177), .ZN(n4175) );
  OAI222_X1 U4385 ( .A1(n16864), .A2(n1579), .B1(n849), .B2(n16858), .C1(n653), 
        .C2(n1104), .ZN(n4177) );
  OAI21_X1 U4386 ( .B1(n4178), .B2(n16824), .A(n1230), .ZN(n4176) );
  NAND2_X1 U4387 ( .A1(n16866), .A2(n16851), .ZN(n1230) );
  NOR2_X1 U4388 ( .A1(n16864), .A2(n16834), .ZN(n1803) );
  AND3_X1 U4389 ( .A1(n4178), .A2(n16829), .A3(n4179), .ZN(n1801) );
  INV_X1 U4390 ( .A(n1606), .ZN(n4178) );
  NOR2_X1 U4391 ( .A1(n16842), .A2(n1086), .ZN(n1606) );
  NOR2_X1 U4392 ( .A1(n88), .A2(n86), .ZN(n84) );
  NOR2_X1 U4393 ( .A1(n499), .A2(n1040), .ZN(n86) );
  NOR3_X1 U4394 ( .A1(n16671), .A2(n1348), .A3(n16656), .ZN(n88) );
  INV_X1 U4396 ( .A(n2027), .ZN(n1348) );
  OAI21_X1 U4397 ( .B1(n16851), .B2(n891), .A(n4180), .ZN(n2027) );
  NAND3_X1 U4398 ( .A1(n566), .A2(n16862), .A3(n563), .ZN(n4180) );
  NOR2_X1 U4399 ( .A1(n851), .A2(n16834), .ZN(n566) );
  NAND2_X1 U4400 ( .A1(n760), .A2(n17096), .ZN(n891) );
  OAI22_X1 U4401 ( .A1(n4956), .A2(n4181), .B1(n4182), .B2(n1096), .ZN(
        U227_Z_0) );
  NOR4_X1 U4403 ( .A1(n4183), .A2(n17092), .A3(rxev_i), .A4(txev_o), .ZN(n4182) );
  OAI21_X1 U4405 ( .B1(n5168), .B2(n4184), .A(n1314), .ZN(n4183) );
  NOR2_X1 U4407 ( .A1(n1092), .A2(n605), .ZN(n1125) );
  NAND2_X1 U4408 ( .A1(n16851), .A2(n16855), .ZN(n605) );
  NAND2_X1 U4409 ( .A1(n997), .A2(n527), .ZN(n1092) );
  NOR4_X1 U4410 ( .A1(n4185), .A2(n4186), .A3(n4187), .A4(n4188), .ZN(n4184)
         );
  INV_X1 U4411 ( .A(n4189), .ZN(n4188) );
  AOI222_X1 U4412 ( .A1(n4965), .A2(n11928), .B1(n5526), .B2(n4893), .C1(n5005), .C2(n11929), .ZN(n4189) );
  AOI21_X1 U4413 ( .B1(n1318), .B2(n17092), .A(n4190), .ZN(n11929) );
  AOI21_X1 U4414 ( .B1(n1310), .B2(irq_i[0]), .A(n4191), .ZN(n4190) );
  AOI22_X1 U4415 ( .A1(n1316), .A2(n5005), .B1(hwdata_o[0]), .B2(n4192), .ZN(
        n4191) );
  NAND2_X1 U4416 ( .A1(hwdata_o[0]), .A2(n1124), .ZN(n1316) );
  AOI21_X1 U4420 ( .B1(n1392), .B2(n17092), .A(n4193), .ZN(n4893) );
  AOI21_X1 U4421 ( .B1(irq_i[3]), .B2(n5525), .A(n4194), .ZN(n4193) );
  AOI22_X1 U4422 ( .A1(n1390), .A2(n5526), .B1(hwdata_o[3]), .B2(n4192), .ZN(
        n4194) );
  NAND2_X1 U4423 ( .A1(hwdata_o[3]), .A2(n1124), .ZN(n1390) );
  AOI21_X1 U4426 ( .B1(n4965), .B2(n4195), .A(n1429), .ZN(n11928) );
  NOR2_X1 U4427 ( .A1(n200), .A2(n183), .ZN(n1429) );
  NAND2_X1 U4428 ( .A1(n1343), .A2(n186), .ZN(n183) );
  AOI21_X1 U4429 ( .B1(n4964), .B2(nmi_i), .A(n1428), .ZN(n4195) );
  NOR2_X1 U4430 ( .A1(n1187), .A2(n3962), .ZN(n1428) );
  OAI221_X1 U4431 ( .B1(n1012), .B2(n3066), .C1(n3238), .C2(n4196), .A(n4197), 
        .ZN(n4187) );
  OAI21_X1 U4432 ( .B1(n4198), .B2(n4199), .A(n1124), .ZN(n4197) );
  NAND4_X1 U4433 ( .A1(n19), .A2(n1190), .A3(n4200), .A4(n4201), .ZN(n4199) );
  NOR3_X1 U4434 ( .A1(hwdata_o[30]), .A2(hwdata_o[19]), .A3(hwdata_o[21]), 
        .ZN(n4201) );
  NAND4_X1 U4437 ( .A1(n4204), .A2(n4205), .A3(n4206), .A4(n4207), .ZN(n21) );
  AOI221_X1 U4438 ( .B1(n16917), .B2(vis_r4_o[21]), .C1(n16914), .C2(
        vis_r5_o[21]), .A(n4210), .ZN(n4207) );
  OAI222_X1 U4439 ( .A1(n4765), .A2(n16910), .B1(n5185), .B2(n16907), .C1(
        n5466), .C2(n16904), .ZN(n4210) );
  AOI221_X1 U4442 ( .B1(n16901), .B2(vis_psp_o[19]), .C1(n16898), .C2(
        vis_r10_o[21]), .A(n4216), .ZN(n4206) );
  OAI22_X1 U4443 ( .A1(n5622), .A2(n16896), .B1(n5623), .B2(n16892), .ZN(n4216) );
  AOI221_X1 U4446 ( .B1(n16890), .B2(vis_r9_o[21]), .C1(n16887), .C2(
        vis_r12_o[21]), .A(n4221), .ZN(n4205) );
  OAI22_X1 U4447 ( .A1(n5115), .A2(n16884), .B1(n5408), .B2(n16881), .ZN(n4221) );
  AOI221_X1 U4450 ( .B1(n4224), .B2(vis_r0_o[21]), .C1(n16878), .C2(
        vis_r3_o[21]), .A(n4227), .ZN(n4204) );
  OAI22_X1 U4451 ( .A1(n5117), .A2(n16876), .B1(n5321), .B2(n16873), .ZN(n4227) );
  NAND4_X1 U4456 ( .A1(n4230), .A2(n4231), .A3(n4232), .A4(n4233), .ZN(n22) );
  AOI221_X1 U4457 ( .B1(n16917), .B2(vis_r4_o[19]), .C1(n16914), .C2(
        vis_r5_o[19]), .A(n4234), .ZN(n4233) );
  OAI222_X1 U4458 ( .A1(n4767), .A2(n16909), .B1(n5186), .B2(n16906), .C1(
        n5467), .C2(n16903), .ZN(n4234) );
  AOI221_X1 U4461 ( .B1(n16900), .B2(vis_psp_o[17]), .C1(n16897), .C2(
        vis_r10_o[19]), .A(n4235), .ZN(n4232) );
  OAI22_X1 U4462 ( .A1(n5636), .A2(n16896), .B1(n5637), .B2(n16892), .ZN(n4235) );
  AOI221_X1 U4465 ( .B1(n16889), .B2(vis_r9_o[19]), .C1(n16886), .C2(
        vis_r12_o[19]), .A(n4236), .ZN(n4231) );
  OAI22_X1 U4466 ( .A1(n5088), .A2(n16883), .B1(n5409), .B2(n16881), .ZN(n4236) );
  AOI221_X1 U4469 ( .B1(n4224), .B2(vis_r0_o[19]), .C1(n16877), .C2(
        vis_r3_o[19]), .A(n4238), .ZN(n4230) );
  OAI22_X1 U4470 ( .A1(n5090), .A2(n16876), .B1(n5322), .B2(n16873), .ZN(n4238) );
  INV_X1 U4475 ( .A(n18), .ZN(n4200) );
  NAND3_X1 U4476 ( .A1(n1187), .A2(n1115), .A3(n4241), .ZN(n18) );
  NOR3_X1 U4477 ( .A1(hwdata_o[25]), .A2(hwdata_o[28]), .A3(hwdata_o[27]), 
        .ZN(n4241) );
  AOI222_X1 U4479 ( .A1(n2257), .A2(n16786), .B1(n2246), .B2(n4240), .C1(n2427), .C2(n4203), .ZN(n208) );
  AOI222_X1 U4482 ( .A1(n3287), .A2(n4240), .B1(n2248), .B2(n4203), .C1(n2028), 
        .C2(n16786), .ZN(n201) );
  NAND4_X1 U4483 ( .A1(n4242), .A2(n4243), .A3(n4244), .A4(n4245), .ZN(n2248)
         );
  AOI221_X1 U4484 ( .B1(n16917), .B2(vis_r4_o[25]), .C1(n16914), .C2(
        vis_r5_o[25]), .A(n4246), .ZN(n4245) );
  OAI222_X1 U4485 ( .A1(n4763), .A2(n16909), .B1(n5178), .B2(n16906), .C1(
        n5459), .C2(n16903), .ZN(n4246) );
  AOI221_X1 U4488 ( .B1(n16900), .B2(vis_psp_o[23]), .C1(n16898), .C2(
        vis_r10_o[25]), .A(n4247), .ZN(n4244) );
  OAI22_X1 U4489 ( .A1(n5291), .A2(n16896), .B1(n5015), .B2(n16893), .ZN(n4247) );
  AOI221_X1 U4492 ( .B1(n16889), .B2(vis_r9_o[25]), .C1(n16887), .C2(
        vis_r12_o[25]), .A(n4248), .ZN(n4243) );
  OAI22_X1 U4493 ( .A1(n5012), .A2(n16883), .B1(n5401), .B2(n16882), .ZN(n4248) );
  AOI221_X1 U4496 ( .B1(n16880), .B2(vis_r0_o[25]), .C1(n16878), .C2(
        vis_r3_o[25]), .A(n4250), .ZN(n4242) );
  OAI22_X1 U4497 ( .A1(n5014), .A2(n16875), .B1(n5314), .B2(n16874), .ZN(n4250) );
  NAND4_X1 U4501 ( .A1(n4251), .A2(n4252), .A3(n4253), .A4(n4254), .ZN(n2249)
         );
  AOI221_X1 U4502 ( .B1(n16917), .B2(vis_r4_o[18]), .C1(n16914), .C2(
        vis_r5_o[18]), .A(n4255), .ZN(n4254) );
  OAI222_X1 U4503 ( .A1(n4768), .A2(n16909), .B1(n5187), .B2(n16906), .C1(
        n5468), .C2(n16903), .ZN(n4255) );
  AOI221_X1 U4506 ( .B1(n16900), .B2(vis_psp_o[16]), .C1(n16898), .C2(
        vis_r10_o[18]), .A(n4256), .ZN(n4253) );
  OAI22_X1 U4507 ( .A1(n5297), .A2(n16896), .B1(n5065), .B2(n16893), .ZN(n4256) );
  AOI221_X1 U4510 ( .B1(n16889), .B2(vis_r9_o[18]), .C1(n16887), .C2(
        vis_r12_o[18]), .A(n4257), .ZN(n4252) );
  OAI22_X1 U4511 ( .A1(n5062), .A2(n16883), .B1(n5410), .B2(n16882), .ZN(n4257) );
  AOI221_X1 U4514 ( .B1(n16880), .B2(vis_r0_o[18]), .C1(n16878), .C2(
        vis_r3_o[18]), .A(n4259), .ZN(n4251) );
  OAI22_X1 U4515 ( .A1(n5064), .A2(n16875), .B1(n5323), .B2(n16874), .ZN(n4259) );
  NAND2_X1 U4518 ( .A1(n253), .A2(hwdata_o[31]), .ZN(n1187) );
  AOI222_X1 U4520 ( .A1(n2196), .A2(n16786), .B1(n2254), .B2(n4240), .C1(n3534), .C2(n4203), .ZN(n4260) );
  INV_X1 U4521 ( .A(n13), .ZN(n1190) );
  NOR2_X1 U4522 ( .A1(n5007), .A2(n4261), .ZN(n13) );
  NAND4_X1 U4524 ( .A1(n4262), .A2(n4263), .A3(n4264), .A4(n4265), .ZN(n2251)
         );
  AOI221_X1 U4525 ( .B1(n16917), .B2(vis_r4_o[22]), .C1(n16914), .C2(
        vis_r5_o[22]), .A(n4266), .ZN(n4265) );
  OAI222_X1 U4526 ( .A1(n4764), .A2(n16909), .B1(n5184), .B2(n16906), .C1(
        n5465), .C2(n16903), .ZN(n4266) );
  AOI221_X1 U4529 ( .B1(n16900), .B2(vis_psp_o[20]), .C1(n16897), .C2(
        vis_r10_o[22]), .A(n4267), .ZN(n4264) );
  OAI22_X1 U4530 ( .A1(n5296), .A2(n16895), .B1(n5051), .B2(n16893), .ZN(n4267) );
  AOI221_X1 U4533 ( .B1(n16889), .B2(vis_r9_o[22]), .C1(n16886), .C2(
        vis_r12_o[22]), .A(n4268), .ZN(n4263) );
  OAI22_X1 U4534 ( .A1(n5048), .A2(n16883), .B1(n5407), .B2(n16882), .ZN(n4268) );
  AOI221_X1 U4537 ( .B1(n16880), .B2(vis_r0_o[22]), .C1(n16877), .C2(
        vis_r3_o[22]), .A(n4270), .ZN(n4262) );
  OAI22_X1 U4538 ( .A1(n5050), .A2(n16875), .B1(n5320), .B2(n16874), .ZN(n4270) );
  NAND4_X1 U4541 ( .A1(n1112), .A2(n1118), .A3(n1117), .A4(n4271), .ZN(n4198)
         );
  NOR3_X1 U4542 ( .A1(hwdata_o[24]), .A2(hwdata_o[29]), .A3(hwdata_o[26]), 
        .ZN(n4271) );
  AOI222_X1 U4545 ( .A1(n2556), .A2(n16786), .B1(n2259), .B2(n4240), .C1(n1755), .C2(n4203), .ZN(n4272) );
  AOI222_X1 U4547 ( .A1(n1354), .A2(n16786), .B1(n2261), .B2(n4240), .C1(n2496), .C2(n4203), .ZN(n25) );
  NAND4_X1 U4549 ( .A1(n4273), .A2(n4274), .A3(n4275), .A4(n4276), .ZN(n20) );
  AOI221_X1 U4550 ( .B1(n16917), .B2(vis_r4_o[20]), .C1(n16914), .C2(
        vis_r5_o[20]), .A(n4277), .ZN(n4276) );
  OAI222_X1 U4551 ( .A1(n4766), .A2(n16909), .B1(n5612), .B2(n16906), .C1(
        n5604), .C2(n16903), .ZN(n4277) );
  AOI221_X1 U4554 ( .B1(n16900), .B2(vis_psp_o[18]), .C1(n16898), .C2(
        vis_r10_o[20]), .A(n4278), .ZN(n4275) );
  OAI22_X1 U4555 ( .A1(n5615), .A2(n16895), .B1(n5616), .B2(n16893), .ZN(n4278) );
  AOI221_X1 U4558 ( .B1(n16889), .B2(vis_r9_o[20]), .C1(n16887), .C2(
        vis_r12_o[20]), .A(n4279), .ZN(n4274) );
  OAI22_X1 U4559 ( .A1(n5603), .A2(n16883), .B1(n5606), .B2(n16882), .ZN(n4279) );
  AOI221_X1 U4562 ( .B1(n16880), .B2(vis_r0_o[20]), .C1(n16878), .C2(
        vis_r3_o[20]), .A(n4281), .ZN(n4273) );
  OAI22_X1 U4563 ( .A1(n5613), .A2(n16875), .B1(n5609), .B2(n16874), .ZN(n4281) );
  NAND4_X1 U4567 ( .A1(n4282), .A2(n4283), .A3(n4284), .A4(n4285), .ZN(n17) );
  AOI221_X1 U4568 ( .B1(n16917), .B2(vis_r4_o[16]), .C1(n16914), .C2(
        vis_r5_o[16]), .A(n4286), .ZN(n4285) );
  OAI222_X1 U4569 ( .A1(n4770), .A2(n16909), .B1(n5189), .B2(n16906), .C1(
        n5470), .C2(n16903), .ZN(n4286) );
  AOI221_X1 U4572 ( .B1(n16900), .B2(vis_psp_o[14]), .C1(n16898), .C2(
        vis_r10_o[16]), .A(n4287), .ZN(n4284) );
  OAI22_X1 U4573 ( .A1(n5299), .A2(n16895), .B1(n5072), .B2(n16893), .ZN(n4287) );
  AOI221_X1 U4576 ( .B1(n16889), .B2(vis_r9_o[16]), .C1(n16887), .C2(
        vis_r12_o[16]), .A(n4288), .ZN(n4283) );
  OAI22_X1 U4577 ( .A1(n5069), .A2(n16883), .B1(n5412), .B2(n16882), .ZN(n4288) );
  AOI221_X1 U4580 ( .B1(n16880), .B2(vis_r0_o[16]), .C1(n16878), .C2(
        vis_r3_o[16]), .A(n4290), .ZN(n4282) );
  OAI22_X1 U4581 ( .A1(n5071), .A2(n16875), .B1(n5325), .B2(n16874), .ZN(n4290) );
  NAND4_X1 U4585 ( .A1(n4291), .A2(n4292), .A3(n4293), .A4(n4294), .ZN(n2258)
         );
  AOI221_X1 U4586 ( .B1(n16917), .B2(vis_r4_o[17]), .C1(n16914), .C2(
        vis_r5_o[17]), .A(n4295), .ZN(n4294) );
  OAI222_X1 U4587 ( .A1(n4769), .A2(n16909), .B1(n5188), .B2(n16906), .C1(
        n5469), .C2(n16903), .ZN(n4295) );
  AOI221_X1 U4590 ( .B1(n16900), .B2(vis_psp_o[15]), .C1(n16898), .C2(
        vis_r10_o[17]), .A(n4296), .ZN(n4293) );
  OAI22_X1 U4591 ( .A1(n5298), .A2(n16895), .B1(n5086), .B2(n16893), .ZN(n4296) );
  AOI221_X1 U4594 ( .B1(n16889), .B2(vis_r9_o[17]), .C1(n16887), .C2(
        vis_r12_o[17]), .A(n4297), .ZN(n4292) );
  OAI22_X1 U4595 ( .A1(n5083), .A2(n16883), .B1(n5411), .B2(n16882), .ZN(n4297) );
  AOI221_X1 U4598 ( .B1(n16880), .B2(vis_r0_o[17]), .C1(n16878), .C2(
        vis_r3_o[17]), .A(n4299), .ZN(n4291) );
  OAI22_X1 U4599 ( .A1(n5085), .A2(n16875), .B1(n5324), .B2(n16874), .ZN(n4299) );
  INV_X1 U4602 ( .A(n4894), .ZN(n4196) );
  AOI21_X1 U4603 ( .B1(n1398), .B2(n17092), .A(n4300), .ZN(n4894) );
  AOI21_X1 U4604 ( .B1(irq_i[2]), .B2(n5527), .A(n4301), .ZN(n4300) );
  AOI22_X1 U4605 ( .A1(n1396), .A2(n5528), .B1(hwdata_o[2]), .B2(n4192), .ZN(
        n4301) );
  NAND2_X1 U4606 ( .A1(hwdata_o[2]), .A2(n1124), .ZN(n1396) );
  INV_X1 U4611 ( .A(n4302), .ZN(n1012) );
  OAI221_X1 U4612 ( .B1(n4303), .B2(n4304), .C1(n559), .C2(n4305), .A(n4306), 
        .ZN(n4302) );
  OAI21_X1 U4613 ( .B1(n1866), .B2(n4307), .A(n5228), .ZN(n4306) );
  OAI33_X1 U4614 ( .A1(n4179), .A2(n16802), .A3(n4308), .B1(n4309), .B2(n585), 
        .B3(n532), .ZN(n4307) );
  OR2_X1 U4615 ( .A1(n1856), .A2(n918), .ZN(n4309) );
  NAND2_X1 U4616 ( .A1(n16825), .A2(n16842), .ZN(n1856) );
  NAND2_X1 U4617 ( .A1(n1574), .A2(n16690), .ZN(n4179) );
  OAI211_X1 U4618 ( .C1(n559), .C2(n4310), .A(n4311), .B(n4312), .ZN(n1866) );
  NOR2_X1 U4619 ( .A1(n1839), .A2(n4313), .ZN(n4312) );
  NOR4_X1 U4620 ( .A1(n4314), .A2(n532), .A3(n1469), .A4(n604), .ZN(n4313) );
  AOI21_X1 U4621 ( .B1(n781), .B2(n659), .A(n669), .ZN(n1469) );
  NAND2_X1 U4623 ( .A1(n760), .A2(n466), .ZN(n4314) );
  INV_X1 U4624 ( .A(n2658), .ZN(n1839) );
  OAI21_X1 U4625 ( .B1(n667), .B2(n991), .A(n909), .ZN(n2658) );
  INV_X1 U4626 ( .A(n1541), .ZN(n909) );
  NAND2_X1 U4627 ( .A1(n16806), .A2(n16808), .ZN(n1541) );
  NAND3_X1 U4628 ( .A1(n4315), .A2(n16826), .A3(n4316), .ZN(n4311) );
  INV_X1 U4629 ( .A(n4308), .ZN(n4316) );
  NAND3_X1 U4630 ( .A1(n592), .A2(n1094), .A3(n501), .ZN(n4308) );
  OAI21_X1 U4631 ( .B1(n16725), .B2(n603), .A(n2673), .ZN(n4315) );
  NOR2_X1 U4632 ( .A1(n602), .A2(n475), .ZN(n2673) );
  OAI21_X1 U4633 ( .B1(n16802), .B2(n16659), .A(n711), .ZN(n602) );
  NAND2_X1 U4634 ( .A1(n16804), .A2(n16725), .ZN(n711) );
  NAND2_X1 U4635 ( .A1(n4974), .A2(n16802), .ZN(n603) );
  INV_X1 U4636 ( .A(n930), .ZN(n559) );
  NAND2_X1 U4637 ( .A1(n17096), .A2(n16808), .ZN(n4304) );
  AOI22_X1 U4639 ( .A1(n5167), .A2(n4317), .B1(n5228), .B2(n1063), .ZN(n4303)
         );
  NAND2_X1 U4640 ( .A1(n1040), .A2(n1343), .ZN(n4317) );
  INV_X1 U4641 ( .A(n181), .ZN(n1343) );
  INV_X1 U4642 ( .A(n1058), .ZN(n1040) );
  NAND4_X1 U4643 ( .A1(n4318), .A2(n1860), .A3(n4319), .A4(n4320), .ZN(n1058)
         );
  AOI22_X1 U4644 ( .A1(n1173), .A2(n16862), .B1(n528), .B2(n529), .ZN(n4320)
         );
  INV_X1 U4645 ( .A(n692), .ZN(n528) );
  AND3_X1 U4646 ( .A1(n563), .A2(n16829), .A3(n1034), .ZN(n1173) );
  NOR2_X1 U4647 ( .A1(n16826), .A2(n16839), .ZN(n1034) );
  NAND4_X1 U4648 ( .A1(n809), .A2(n760), .A3(n16821), .A4(n16856), .ZN(n4319)
         );
  INV_X1 U4649 ( .A(n1473), .ZN(n1860) );
  NOR3_X1 U4650 ( .A1(n745), .A2(n5165), .A3(n641), .ZN(n1473) );
  INV_X1 U4651 ( .A(n4321), .ZN(n4186) );
  AOI221_X1 U4652 ( .B1(n11971), .B2(n5572), .C1(n4900), .C2(n4749), .A(n4322), 
        .ZN(n4321) );
  INV_X1 U4653 ( .A(n4323), .ZN(n4322) );
  AOI222_X1 U4654 ( .A1(n5011), .A2(n11957), .B1(n11939), .B2(n5534), .C1(
        n11945), .C2(n5533), .ZN(n4323) );
  AOI21_X1 U4655 ( .B1(n1419), .B2(n17092), .A(n4324), .ZN(n11945) );
  AOI21_X1 U4656 ( .B1(n1411), .B2(irq_i[5]), .A(n4325), .ZN(n4324) );
  AOI22_X1 U4657 ( .A1(n1416), .A2(n5533), .B1(hwdata_o[5]), .B2(n4192), .ZN(
        n4325) );
  NAND2_X1 U4658 ( .A1(hwdata_o[5]), .A2(n1124), .ZN(n1416) );
  AOI21_X1 U4662 ( .B1(n1453), .B2(n17092), .A(n4326), .ZN(n11939) );
  AOI21_X1 U4663 ( .B1(n1447), .B2(irq_i[1]), .A(n4327), .ZN(n4326) );
  AOI22_X1 U4664 ( .A1(n1452), .A2(n5534), .B1(hwdata_o[1]), .B2(n4192), .ZN(
        n4327) );
  NAND2_X1 U4665 ( .A1(hwdata_o[1]), .A2(n1124), .ZN(n1452) );
  NOR2_X1 U4669 ( .A1(n4328), .A2(n1128), .ZN(n11957) );
  NOR2_X1 U4670 ( .A1(n200), .A2(n4329), .ZN(n1128) );
  AOI221_X1 U4671 ( .B1(hwdata_o[9]), .B2(n1124), .C1(n5580), .C2(irq_i[9]), 
        .A(n4330), .ZN(n4328) );
  AOI21_X1 U4672 ( .B1(hwdata_o[9]), .B2(n4192), .A(n5011), .ZN(n4330) );
  AOI21_X1 U4673 ( .B1(n1446), .B2(n17092), .A(n4331), .ZN(n4900) );
  INV_X1 U4674 ( .A(n4332), .ZN(n4331) );
  OAI221_X1 U4675 ( .B1(n240), .B2(n1385), .C1(n1444), .C2(n4333), .A(n4334), 
        .ZN(n4332) );
  OAI21_X1 U4676 ( .B1(n240), .B2(n4335), .A(n3089), .ZN(n4334) );
  INV_X1 U4679 ( .A(irq_i[12]), .ZN(n1444) );
  NOR2_X1 U4680 ( .A1(n4336), .A2(n1432), .ZN(n11971) );
  NOR2_X1 U4681 ( .A1(n200), .A2(n4337), .ZN(n1432) );
  AOI221_X1 U4682 ( .B1(hwdata_o[11]), .B2(n1124), .C1(n4338), .C2(irq_i[11]), 
        .A(n4339), .ZN(n4336) );
  AOI21_X1 U4683 ( .B1(hwdata_o[11]), .B2(n4192), .A(n5572), .ZN(n4339) );
  NAND4_X1 U4685 ( .A1(n4340), .A2(n4341), .A3(n4342), .A4(n4343), .ZN(n4185)
         );
  AOI21_X1 U4686 ( .B1(n4748), .B2(n4344), .A(n4345), .ZN(n4343) );
  OAI33_X1 U4687 ( .A1(n202), .A2(n205), .A3(n209), .B1(n1053), .B2(n1050), 
        .B3(n930), .ZN(n4345) );
  OAI211_X1 U4688 ( .C1(n4346), .C2(n4347), .A(n181), .B(n1045), .ZN(n930) );
  NAND4_X1 U4690 ( .A1(vis_ipsr_o[1]), .A2(n176), .A3(n4348), .A4(n170), .ZN(
        n181) );
  AOI22_X1 U4691 ( .A1(n4349), .A2(n3732), .B1(n1355), .B2(n4350), .ZN(n4347)
         );
  OR2_X1 U4692 ( .A1(n4350), .A2(n1355), .ZN(n4349) );
  NOR4_X1 U4693 ( .A1(n4351), .A2(n4352), .A3(n4353), .A4(n4354), .ZN(n1355)
         );
  OAI221_X1 U4694 ( .B1(n5153), .B2(n1456), .C1(n5098), .C2(n199), .A(n4355), 
        .ZN(n4354) );
  AOI222_X1 U4695 ( .A1(n1378), .A2(n3791), .B1(n1386), .B2(n4356), .C1(n1404), 
        .C2(n3862), .ZN(n4355) );
  OAI221_X1 U4699 ( .B1(n5023), .B2(n1415), .C1(n5547), .C2(n1451), .A(n4357), 
        .ZN(n4353) );
  AOI222_X1 U4700 ( .A1(n1122), .A2(n3793), .B1(n4358), .B2(n3732), .C1(n1430), 
        .C2(n3792), .ZN(n4357) );
  OAI221_X1 U4704 ( .B1(n5522), .B2(n1441), .C1(n5523), .C2(n1423), .A(n4359), 
        .ZN(n4352) );
  AOI22_X1 U4705 ( .A1(n1318), .A2(n3847), .B1(n1392), .B2(n3833), .ZN(n4359)
         );
  INV_X1 U4707 ( .A(n1391), .ZN(n1392) );
  OAI221_X1 U4709 ( .B1(n5551), .B2(n1397), .C1(n4961), .C2(n207), .A(n4360), 
        .ZN(n4351) );
  AOI222_X1 U4710 ( .A1(n1410), .A2(n3863), .B1(n1446), .B2(n3784), .C1(n1126), 
        .C2(n3813), .ZN(n4360) );
  INV_X1 U4712 ( .A(n4329), .ZN(n1126) );
  INV_X1 U4714 ( .A(n1445), .ZN(n1446) );
  NAND2_X1 U4716 ( .A1(n5503), .A2(n4361), .ZN(n4350) );
  NAND4_X1 U4717 ( .A1(n1362), .A2(n1363), .A3(n1365), .A4(n1367), .ZN(n4361)
         );
  AOI221_X1 U4718 ( .B1(n2931), .B2(n1404), .C1(n2888), .C2(n1122), .A(n4362), 
        .ZN(n1367) );
  OAI22_X1 U4719 ( .A1(n4337), .A2(n5160), .B1(n1384), .B2(n5151), .ZN(n4362)
         );
  INV_X1 U4722 ( .A(n4363), .ZN(n1365) );
  OAI221_X1 U4723 ( .B1(n5152), .B2(n1456), .C1(n1445), .C2(n1885), .A(n4364), 
        .ZN(n4363) );
  AOI222_X1 U4724 ( .A1(n1378), .A2(n2927), .B1(n4365), .B2(n2929), .C1(n4366), 
        .C2(n2889), .ZN(n4364) );
  AOI221_X1 U4729 ( .B1(n4367), .B2(n1410), .C1(n2902), .C2(n1419), .A(n4368), 
        .ZN(n1363) );
  OAI222_X1 U4730 ( .A1(n1423), .A2(n5519), .B1(n1441), .B2(n5518), .C1(n4329), 
        .C2(n5157), .ZN(n4368) );
  INV_X1 U4731 ( .A(n1415), .ZN(n1419) );
  AOI221_X1 U4734 ( .B1(n1398), .B2(n4752), .C1(n2951), .C2(n1318), .A(n4369), 
        .ZN(n1362) );
  OAI22_X1 U4735 ( .A1(n1451), .A2(n5550), .B1(n1391), .B2(n5552), .ZN(n4369)
         );
  INV_X1 U4737 ( .A(n1358), .ZN(n4346) );
  NAND4_X1 U4738 ( .A1(n4370), .A2(n4371), .A3(n4372), .A4(n4373), .ZN(n1358)
         );
  NOR4_X1 U4739 ( .A1(n4374), .A2(n1453), .A3(n4366), .A4(n4365), .ZN(n4373)
         );
  INV_X1 U4740 ( .A(n199), .ZN(n4365) );
  NAND2_X1 U4741 ( .A1(n4375), .A2(n4376), .ZN(n199) );
  INV_X1 U4742 ( .A(n207), .ZN(n4366) );
  NAND2_X1 U4743 ( .A1(n4377), .A2(n4376), .ZN(n207) );
  INV_X1 U4744 ( .A(n1451), .ZN(n1453) );
  NAND2_X1 U4745 ( .A1(n4378), .A2(n4379), .ZN(n1451) );
  NAND2_X1 U4746 ( .A1(n1391), .A2(n1415), .ZN(n4374) );
  NAND2_X1 U4747 ( .A1(n4379), .A2(n4375), .ZN(n1415) );
  NAND2_X1 U4748 ( .A1(n4380), .A2(n4378), .ZN(n1391) );
  NOR4_X1 U4749 ( .A1(n4381), .A2(n1410), .A3(n1318), .A4(n1398), .ZN(n4372)
         );
  INV_X1 U4750 ( .A(n1397), .ZN(n1398) );
  NAND2_X1 U4751 ( .A1(n4382), .A2(n4380), .ZN(n1397) );
  INV_X1 U4752 ( .A(n1315), .ZN(n1318) );
  NAND2_X1 U4753 ( .A1(n4382), .A2(n4379), .ZN(n1315) );
  NAND2_X1 U4754 ( .A1(n4329), .A2(n1423), .ZN(n4381) );
  NAND2_X1 U4755 ( .A1(n4383), .A2(n4378), .ZN(n4329) );
  NOR3_X1 U4756 ( .A1(n4384), .A2(n1378), .A3(n1122), .ZN(n4371) );
  INV_X1 U4757 ( .A(n1436), .ZN(n1122) );
  NAND2_X1 U4758 ( .A1(n4385), .A2(n4382), .ZN(n1436) );
  NAND3_X1 U4759 ( .A1(n1445), .A2(n1441), .A3(n1456), .ZN(n4384) );
  NAND2_X1 U4760 ( .A1(n4383), .A2(n4382), .ZN(n1441) );
  NAND2_X1 U4761 ( .A1(n4383), .A2(n4377), .ZN(n1445) );
  NOR4_X1 U4762 ( .A1(n1404), .A2(n1386), .A3(n1430), .A4(n4358), .ZN(n4370)
         );
  INV_X1 U4763 ( .A(n1052), .ZN(n4358) );
  NAND2_X1 U4764 ( .A1(n4378), .A2(n4376), .ZN(n1052) );
  NOR4_X1 U4765 ( .A1(n170), .A2(n191), .A3(vis_ipsr_o[4]), .A4(vis_ipsr_o[5]), 
        .ZN(n4376) );
  INV_X1 U4766 ( .A(n4337), .ZN(n1430) );
  NAND2_X1 U4767 ( .A1(n4385), .A2(n4378), .ZN(n4337) );
  NOR2_X1 U4768 ( .A1(n186), .A2(vis_ipsr_o[2]), .ZN(n4378) );
  AND2_X1 U4769 ( .A1(n4305), .A2(n4310), .ZN(n1050) );
  NAND3_X1 U4770 ( .A1(n827), .A2(n914), .A3(n542), .ZN(n4310) );
  NOR2_X1 U4771 ( .A1(n16842), .A2(n16856), .ZN(n542) );
  INV_X1 U4772 ( .A(n762), .ZN(n914) );
  NAND2_X1 U4773 ( .A1(n16806), .A2(n16870), .ZN(n762) );
  NAND4_X1 U4775 ( .A1(n563), .A2(n16823), .A3(n16819), .A4(n3509), .ZN(n4305)
         );
  INV_X1 U4776 ( .A(n1088), .ZN(n3509) );
  NAND3_X1 U4777 ( .A1(n991), .A2(n1574), .A3(n16862), .ZN(n1088) );
  NAND2_X1 U4781 ( .A1(n16845), .A2(n16694), .ZN(n1234) );
  AOI222_X1 U4784 ( .A1(n2578), .A2(n16786), .B1(n2247), .B2(n4240), .C1(n89), 
        .C2(n4203), .ZN(n205) );
  INV_X1 U4785 ( .A(n1123), .ZN(n4344) );
  AOI221_X1 U4786 ( .B1(hwdata_o[10]), .B2(n1124), .C1(irq_i[10]), .C2(n5061), 
        .A(n4386), .ZN(n1123) );
  AOI21_X1 U4787 ( .B1(hwdata_o[10]), .B2(n4192), .A(n4748), .ZN(n4386) );
  AOI222_X1 U4788 ( .A1(n4898), .A2(n5532), .B1(n4899), .B2(n5530), .C1(n4747), 
        .C2(n4387), .ZN(n4342) );
  INV_X1 U4789 ( .A(n1121), .ZN(n4387) );
  AOI221_X1 U4790 ( .B1(hwdata_o[8]), .B2(n1124), .C1(irq_i[8]), .C2(n5582), 
        .A(n4388), .ZN(n1121) );
  AOI21_X1 U4791 ( .B1(hwdata_o[8]), .B2(n4192), .A(n4747), .ZN(n4388) );
  AOI21_X1 U4792 ( .B1(n1404), .B2(n17093), .A(n4389), .ZN(n4899) );
  AOI21_X1 U4793 ( .B1(irq_i[7]), .B2(n5529), .A(n4390), .ZN(n4389) );
  AOI22_X1 U4794 ( .A1(n1403), .A2(n5530), .B1(hwdata_o[7]), .B2(n4192), .ZN(
        n4390) );
  NAND2_X1 U4795 ( .A1(hwdata_o[7]), .A2(n1124), .ZN(n1403) );
  INV_X1 U4798 ( .A(n1402), .ZN(n1404) );
  NAND2_X1 U4799 ( .A1(n4380), .A2(n4375), .ZN(n1402) );
  AOI21_X1 U4800 ( .B1(n1410), .B2(n17093), .A(n4391), .ZN(n4898) );
  AOI21_X1 U4801 ( .B1(irq_i[6]), .B2(n5531), .A(n4392), .ZN(n4391) );
  AOI22_X1 U4802 ( .A1(n1409), .A2(n5532), .B1(hwdata_o[6]), .B2(n4192), .ZN(
        n4392) );
  NAND2_X1 U4803 ( .A1(hwdata_o[6]), .A2(n1124), .ZN(n1409) );
  INV_X1 U4806 ( .A(n1408), .ZN(n1410) );
  NAND2_X1 U4807 ( .A1(n4380), .A2(n4377), .ZN(n1408) );
  AND2_X1 U4808 ( .A1(n4393), .A2(vis_ipsr_o[1]), .ZN(n4380) );
  AOI222_X1 U4809 ( .A1(n5047), .A2(n4896), .B1(n4901), .B2(n4750), .C1(n4897), 
        .C2(n3775), .ZN(n4341) );
  AOI21_X1 U4810 ( .B1(n1386), .B2(n17093), .A(n4394), .ZN(n4897) );
  AOI221_X1 U4811 ( .B1(hwdata_o[13]), .B2(n1124), .C1(irq_i[13]), .C2(n5118), 
        .A(n4395), .ZN(n4394) );
  AOI21_X1 U4812 ( .B1(hwdata_o[13]), .B2(n4192), .A(n3775), .ZN(n4395) );
  INV_X1 U4814 ( .A(n1384), .ZN(n1386) );
  NAND2_X1 U4815 ( .A1(n4383), .A2(n4375), .ZN(n1384) );
  AND2_X1 U4816 ( .A1(n4396), .A2(n191), .ZN(n4383) );
  AOI21_X1 U4817 ( .B1(n1425), .B2(n17093), .A(n4397), .ZN(n4901) );
  AOI21_X1 U4818 ( .B1(irq_i[4]), .B2(n5524), .A(n4398), .ZN(n4397) );
  AOI22_X1 U4819 ( .A1(hwdata_o[4]), .A2(n4192), .B1(n1424), .B2(n4750), .ZN(
        n4398) );
  NAND2_X1 U4820 ( .A1(hwdata_o[4]), .A2(n1124), .ZN(n1424) );
  INV_X1 U4823 ( .A(n1423), .ZN(n1425) );
  NAND2_X1 U4824 ( .A1(n4379), .A2(n4377), .ZN(n1423) );
  AND2_X1 U4825 ( .A1(n4393), .A2(n191), .ZN(n4379) );
  NOR3_X1 U4826 ( .A1(vis_ipsr_o[3]), .A2(vis_ipsr_o[5]), .A3(n165), .ZN(n4393) );
  AOI21_X1 U4827 ( .B1(n1459), .B2(n17092), .A(n4399), .ZN(n4896) );
  AOI221_X1 U4828 ( .B1(n1124), .B2(hwdata_o[14]), .C1(irq_i[14]), .C2(n5619), 
        .A(n4400), .ZN(n4399) );
  AOI21_X1 U4829 ( .B1(hwdata_o[14]), .B2(n4192), .A(n5047), .ZN(n4400) );
  NAND4_X1 U4832 ( .A1(n4402), .A2(n4403), .A3(n4404), .A4(n4405), .ZN(n2253)
         );
  AOI221_X1 U4833 ( .B1(n16917), .B2(vis_r4_o[14]), .C1(n16914), .C2(
        vis_r5_o[14]), .A(n4406), .ZN(n4405) );
  OAI222_X1 U4834 ( .A1(n4850), .A2(n16909), .B1(n5190), .B2(n16906), .C1(
        n5471), .C2(n16903), .ZN(n4406) );
  AOI221_X1 U4837 ( .B1(n16900), .B2(vis_psp_o[12]), .C1(n16898), .C2(
        vis_r10_o[14]), .A(n4407), .ZN(n4404) );
  OAI22_X1 U4838 ( .A1(n5300), .A2(n16895), .B1(n5106), .B2(n16893), .ZN(n4407) );
  AOI221_X1 U4841 ( .B1(n16889), .B2(vis_r9_o[14]), .C1(n16887), .C2(
        vis_r12_o[14]), .A(n4408), .ZN(n4403) );
  OAI22_X1 U4842 ( .A1(n5103), .A2(n16883), .B1(n5413), .B2(n16882), .ZN(n4408) );
  AOI221_X1 U4845 ( .B1(n16880), .B2(vis_r0_o[14]), .C1(n16878), .C2(
        vis_r3_o[14]), .A(n4410), .ZN(n4402) );
  OAI22_X1 U4846 ( .A1(n5105), .A2(n16875), .B1(n5326), .B2(n16874), .ZN(n4410) );
  NAND4_X1 U4849 ( .A1(n4411), .A2(n4412), .A3(n4413), .A4(n4414), .ZN(n2250)
         );
  AOI222_X1 U4850 ( .A1(n16652), .A2(vis_r14_o[6]), .B1(n16911), .B2(n1152), 
        .C1(n16651), .C2(vis_msp_o[4]), .ZN(n4414) );
  AOI22_X1 U4854 ( .A1(n16902), .A2(vis_psp_o[4]), .B1(n16897), .B2(
        vis_r10_o[6]), .ZN(n4413) );
  AOI222_X1 U4857 ( .A1(n16886), .A2(vis_r12_o[6]), .B1(n16648), .B2(
        vis_r8_o[6]), .C1(n16891), .C2(vis_r9_o[6]), .ZN(n4412) );
  AOI21_X1 U4861 ( .B1(n16650), .B2(vis_r11_o[6]), .A(n1794), .ZN(n4411) );
  NAND2_X1 U4862 ( .A1(n4420), .A2(n4421), .ZN(n1794) );
  AOI221_X1 U4863 ( .B1(n16917), .B2(vis_r4_o[6]), .C1(n16914), .C2(
        vis_r5_o[6]), .A(n4422), .ZN(n4421) );
  OAI22_X1 U4864 ( .A1(n5461), .A2(n16905), .B1(n5180), .B2(n16908), .ZN(n4422) );
  AOI221_X1 U4867 ( .B1(n16877), .B2(vis_r3_o[6]), .C1(n16649), .C2(
        vis_r7_o[6]), .A(n4426), .ZN(n4420) );
  OAI22_X1 U4868 ( .A1(n5485), .A2(n4427), .B1(n5041), .B2(n16885), .ZN(n4426)
         );
  INV_X1 U4872 ( .A(n1456), .ZN(n1459) );
  NAND2_X1 U4873 ( .A1(n4385), .A2(n4377), .ZN(n1456) );
  NOR2_X1 U4874 ( .A1(n176), .A2(vis_ipsr_o[0]), .ZN(n4377) );
  AOI22_X1 U4875 ( .A1(n5024), .A2(n4895), .B1(n4988), .B2(n204), .ZN(n4340)
         );
  OAI21_X1 U4876 ( .B1(n24), .B2(n202), .A(n4428), .ZN(n204) );
  OR4_X1 U4877 ( .A1(n259), .A2(n260), .A3(n5516), .A4(n4833), .ZN(n4428) );
  NAND4_X1 U4879 ( .A1(n4429), .A2(n4430), .A3(n4431), .A4(n4432), .ZN(n259)
         );
  NOR4_X1 U4880 ( .A1(n4433), .A2(sub_2068_A_4_), .A3(sub_2068_A_6_), .A4(
        sub_2068_A_5_), .ZN(n4432) );
  NAND3_X1 U4881 ( .A1(n296), .A2(n294), .A3(n298), .ZN(n4433) );
  NOR4_X1 U4885 ( .A1(n4434), .A2(sub_2068_A_20_), .A3(sub_2068_A_22_), .A4(
        sub_2068_A_21_), .ZN(n4431) );
  NAND3_X1 U4886 ( .A1(n308), .A2(n306), .A3(n264), .ZN(n4434) );
  NOR4_X1 U4890 ( .A1(n4435), .A2(sub_2068_A_15_), .A3(sub_2068_A_17_), .A4(
        sub_2068_A_16_), .ZN(n4430) );
  NAND3_X1 U4891 ( .A1(n274), .A2(n310), .A3(n276), .ZN(n4435) );
  NOR3_X1 U4895 ( .A1(n4436), .A2(sub_2068_A_11_), .A3(sub_2068_A_10_), .ZN(
        n4429) );
  NAND3_X1 U4896 ( .A1(n286), .A2(n284), .A3(n288), .ZN(n4436) );
  OR2_X1 U4900 ( .A1(n3962), .A2(n5007), .ZN(n202) );
  NAND3_X1 U4901 ( .A1(n5017), .A2(n251), .A3(n3717), .ZN(n3962) );
  NOR3_X1 U4902 ( .A1(n5502), .A2(n5149), .A3(n3874), .ZN(n3717) );
  AOI222_X1 U4904 ( .A1(n3145), .A2(n4240), .B1(n2260), .B2(n4203), .C1(n3177), 
        .C2(n16786), .ZN(n24) );
  NAND4_X1 U4905 ( .A1(n4437), .A2(n4438), .A3(n4439), .A4(n4440), .ZN(n2260)
         );
  AOI221_X1 U4906 ( .B1(n16916), .B2(vis_r4_o[26]), .C1(n16913), .C2(
        vis_r5_o[26]), .A(n4441), .ZN(n4440) );
  OAI222_X1 U4907 ( .A1(n4762), .A2(n16909), .B1(n5177), .B2(n16906), .C1(
        n5458), .C2(n16903), .ZN(n4441) );
  AOI221_X1 U4910 ( .B1(n16900), .B2(vis_psp_o[24]), .C1(n16898), .C2(
        vis_r10_o[26]), .A(n4442), .ZN(n4439) );
  OAI22_X1 U4911 ( .A1(n5290), .A2(n16895), .B1(n4992), .B2(n16893), .ZN(n4442) );
  AOI221_X1 U4914 ( .B1(n16889), .B2(vis_r9_o[26]), .C1(n16887), .C2(
        vis_r12_o[26]), .A(n4443), .ZN(n4438) );
  OAI22_X1 U4915 ( .A1(n4989), .A2(n16883), .B1(n5400), .B2(n16882), .ZN(n4443) );
  AOI221_X1 U4918 ( .B1(n16880), .B2(vis_r0_o[26]), .C1(n16878), .C2(
        vis_r3_o[26]), .A(n4445), .ZN(n4437) );
  OAI22_X1 U4919 ( .A1(n4991), .A2(n16875), .B1(n5313), .B2(n16874), .ZN(n4445) );
  INV_X1 U4923 ( .A(n1670), .ZN(n1614) );
  AOI21_X1 U4924 ( .B1(n1378), .B2(n17092), .A(n4446), .ZN(n4895) );
  AOI221_X1 U4925 ( .B1(n1124), .B2(hwdata_o[15]), .C1(irq_i[15]), .C2(n5620), 
        .A(n4447), .ZN(n4446) );
  AOI21_X1 U4926 ( .B1(hwdata_o[15]), .B2(n4192), .A(n5024), .ZN(n4447) );
  NAND3_X1 U4928 ( .A1(n1385), .A2(n253), .A3(n3873), .ZN(n4335) );
  NAND4_X1 U4931 ( .A1(n4448), .A2(n4449), .A3(n4450), .A4(n4451), .ZN(n2254)
         );
  AOI221_X1 U4932 ( .B1(n16916), .B2(vis_r4_o[15]), .C1(n16913), .C2(
        vis_r5_o[15]), .A(n4452), .ZN(n4451) );
  OAI222_X1 U4933 ( .A1(n4827), .A2(n16909), .B1(n5197), .B2(n16906), .C1(
        n5478), .C2(n16903), .ZN(n4452) );
  AOI221_X1 U4936 ( .B1(n16900), .B2(vis_psp_o[13]), .C1(n16898), .C2(
        vis_r10_o[15]), .A(n4453), .ZN(n4450) );
  OAI22_X1 U4937 ( .A1(n5632), .A2(n16895), .B1(n5633), .B2(n16893), .ZN(n4453) );
  AOI221_X1 U4940 ( .B1(n16889), .B2(vis_r9_o[15]), .C1(n16887), .C2(
        vis_r12_o[15]), .A(n4454), .ZN(n4449) );
  OAI22_X1 U4941 ( .A1(n5108), .A2(n16883), .B1(n5420), .B2(n16882), .ZN(n4454) );
  AOI221_X1 U4944 ( .B1(n16880), .B2(vis_r0_o[15]), .C1(n16878), .C2(
        vis_r3_o[15]), .A(n4456), .ZN(n4448) );
  OAI22_X1 U4945 ( .A1(n5110), .A2(n16875), .B1(n5333), .B2(n16874), .ZN(n4456) );
  NAND3_X1 U4949 ( .A1(n4905), .A2(n253), .A3(n3873), .ZN(n1385) );
  NOR4_X1 U4950 ( .A1(n3874), .A2(n1110), .A3(n5502), .A4(n5017), .ZN(n3873)
         );
  INV_X1 U4956 ( .A(n568), .ZN(n760) );
  INV_X1 U4957 ( .A(n813), .ZN(n809) );
  NAND2_X1 U4958 ( .A1(n608), .A2(n16831), .ZN(n813) );
  AND2_X1 U4959 ( .A1(n4385), .A2(n4375), .ZN(n1378) );
  NOR2_X1 U4960 ( .A1(n186), .A2(n176), .ZN(n4375) );
  AND2_X1 U4963 ( .A1(n4396), .A2(vis_ipsr_o[1]), .ZN(n4385) );
  NOR3_X1 U4964 ( .A1(n170), .A2(vis_ipsr_o[5]), .A3(n165), .ZN(n4396) );
  NOR4_X1 U4966 ( .A1(n4457), .A2(n1784), .A3(n16850), .A4(n1583), .ZN(n4181)
         );
  NOR3_X1 U4967 ( .A1(n16871), .A2(n16821), .A3(n604), .ZN(n1583) );
  NAND2_X1 U4968 ( .A1(n1097), .A2(n2661), .ZN(n4457) );
  INV_X1 U4969 ( .A(n849), .ZN(n2661) );
  INV_X1 U4970 ( .A(n989), .ZN(n1097) );
  NAND2_X1 U4971 ( .A1(n997), .A2(n16834), .ZN(n989) );
  NAND4_X1 U4974 ( .A1(n4458), .A2(n4459), .A3(n4460), .A4(n4461), .ZN(n2261)
         );
  AOI221_X1 U4975 ( .B1(n16916), .B2(vis_r4_o[8]), .C1(n16913), .C2(
        vis_r5_o[8]), .A(n4462), .ZN(n4461) );
  OAI222_X1 U4976 ( .A1(n4851), .A2(n16910), .B1(n5196), .B2(n16907), .C1(
        n5477), .C2(n16904), .ZN(n4462) );
  AOI221_X1 U4979 ( .B1(n16901), .B2(vis_psp_o[6]), .C1(n16898), .C2(
        vis_r10_o[8]), .A(n4463), .ZN(n4460) );
  OAI22_X1 U4980 ( .A1(n5304), .A2(n16895), .B1(n5138), .B2(n16893), .ZN(n4463) );
  AOI221_X1 U4983 ( .B1(n16890), .B2(vis_r9_o[8]), .C1(n16887), .C2(
        vis_r12_o[8]), .A(n4464), .ZN(n4459) );
  OAI22_X1 U4984 ( .A1(n5135), .A2(n16884), .B1(n5419), .B2(n16882), .ZN(n4464) );
  AOI221_X1 U4987 ( .B1(n16880), .B2(vis_r0_o[8]), .C1(n16878), .C2(
        vis_r3_o[8]), .A(n4466), .ZN(n4458) );
  OAI22_X1 U4988 ( .A1(n5137), .A2(n16875), .B1(n5332), .B2(n16874), .ZN(n4466) );
  NAND4_X1 U4991 ( .A1(n4170), .A2(n4467), .A3(n4468), .A4(n4469), .ZN(n1354)
         );
  AOI221_X1 U4992 ( .B1(n16897), .B2(vis_r10_o[0]), .C1(n16648), .C2(
        vis_r8_o[0]), .A(n4472), .ZN(n4469) );
  OAI22_X1 U4993 ( .A1(n5288), .A2(n16895), .B1(n5101), .B2(n4211), .ZN(n4472)
         );
  AOI22_X1 U4996 ( .A1(n16891), .A2(vis_r9_o[0]), .B1(n16886), .B2(
        vis_r12_o[0]), .ZN(n4468) );
  NAND2_X1 U4999 ( .A1(n16650), .A2(vis_r11_o[0]), .ZN(n4467) );
  AND2_X1 U5001 ( .A1(n4474), .A2(n4475), .ZN(n4170) );
  AOI221_X1 U5002 ( .B1(n16916), .B2(vis_r4_o[0]), .C1(n16913), .C2(
        vis_r5_o[0]), .A(n4476), .ZN(n4475) );
  OAI22_X1 U5003 ( .A1(n5454), .A2(n16905), .B1(n5173), .B2(n16908), .ZN(n4476) );
  AOI221_X1 U5006 ( .B1(n16877), .B2(vis_r3_o[0]), .C1(n16649), .C2(
        vis_r7_o[0]), .A(n4479), .ZN(n4474) );
  OAI22_X1 U5007 ( .A1(n5040), .A2(n4427), .B1(n5039), .B2(n16885), .ZN(n4479)
         );
  NAND4_X1 U5012 ( .A1(n4169), .A2(n4480), .A3(n4481), .A4(n4482), .ZN(n2028)
         );
  AOI221_X1 U5013 ( .B1(n16897), .B2(vis_r10_o[1]), .C1(n16648), .C2(
        vis_r8_o[1]), .A(n4484), .ZN(n4482) );
  OAI22_X1 U5014 ( .A1(n5287), .A2(n16895), .B1(n5255), .B2(n4211), .ZN(n4484)
         );
  AOI22_X1 U5017 ( .A1(n16891), .A2(vis_r9_o[1]), .B1(n16886), .B2(
        vis_r12_o[1]), .ZN(n4481) );
  NAND2_X1 U5020 ( .A1(n16650), .A2(vis_r11_o[1]), .ZN(n4480) );
  AND2_X1 U5022 ( .A1(n4486), .A2(n4487), .ZN(n4169) );
  AOI221_X1 U5023 ( .B1(n16916), .B2(vis_r4_o[1]), .C1(n16913), .C2(
        vis_r5_o[1]), .A(n4488), .ZN(n4487) );
  OAI22_X1 U5024 ( .A1(n5453), .A2(n16905), .B1(n5172), .B2(n16908), .ZN(n4488) );
  AOI221_X1 U5027 ( .B1(n16877), .B2(vis_r3_o[1]), .C1(n16649), .C2(
        vis_r7_o[1]), .A(n4491), .ZN(n4486) );
  OAI22_X1 U5028 ( .A1(n4987), .A2(n4427), .B1(n4986), .B2(n16885), .ZN(n4491)
         );
  NAND4_X1 U5031 ( .A1(n4492), .A2(n4493), .A3(n4494), .A4(n4495), .ZN(n3287)
         );
  AOI221_X1 U5032 ( .B1(n16916), .B2(vis_r4_o[9]), .C1(n16913), .C2(
        vis_r5_o[9]), .A(n4496), .ZN(n4495) );
  OAI222_X1 U5033 ( .A1(n5140), .A2(n16910), .B1(n5195), .B2(n16907), .C1(
        n5476), .C2(n16904), .ZN(n4496) );
  AOI221_X1 U5036 ( .B1(n16901), .B2(vis_psp_o[7]), .C1(n16898), .C2(
        vis_r10_o[9]), .A(n4497), .ZN(n4494) );
  OAI22_X1 U5037 ( .A1(n5575), .A2(n16895), .B1(n5576), .B2(n16893), .ZN(n4497) );
  AOI221_X1 U5040 ( .B1(n16890), .B2(vis_r9_o[9]), .C1(n16887), .C2(
        vis_r12_o[9]), .A(n4498), .ZN(n4493) );
  OAI22_X1 U5041 ( .A1(n5141), .A2(n16884), .B1(n5418), .B2(n16882), .ZN(n4498) );
  AOI221_X1 U5044 ( .B1(n16880), .B2(vis_r0_o[9]), .C1(n16878), .C2(
        vis_r3_o[9]), .A(n4500), .ZN(n4492) );
  OAI22_X1 U5045 ( .A1(n5143), .A2(n16875), .B1(n5331), .B2(n16874), .ZN(n4500) );
  NAND4_X1 U5050 ( .A1(n4501), .A2(n4502), .A3(n4503), .A4(n4504), .ZN(n3145)
         );
  AOI221_X1 U5051 ( .B1(n16916), .B2(vis_r4_o[10]), .C1(n16913), .C2(
        vis_r5_o[10]), .A(n4505), .ZN(n4504) );
  OAI222_X1 U5052 ( .A1(n4771), .A2(n16910), .B1(n5193), .B2(n16907), .C1(
        n5474), .C2(n16904), .ZN(n4505) );
  AOI221_X1 U5055 ( .B1(n16901), .B2(vis_psp_o[8]), .C1(n16899), .C2(
        vis_r10_o[10]), .A(n4506), .ZN(n4503) );
  OAI22_X1 U5056 ( .A1(n5302), .A2(n16894), .B1(n5147), .B2(n16892), .ZN(n4506) );
  AOI221_X1 U5059 ( .B1(n16890), .B2(vis_r9_o[10]), .C1(n16888), .C2(
        vis_r12_o[10]), .A(n4507), .ZN(n4502) );
  OAI22_X1 U5060 ( .A1(n5144), .A2(n16884), .B1(n5416), .B2(n16881), .ZN(n4507) );
  AOI221_X1 U5063 ( .B1(n16880), .B2(vis_r0_o[10]), .C1(n16879), .C2(
        vis_r3_o[10]), .A(n4509), .ZN(n4501) );
  OAI22_X1 U5064 ( .A1(n5146), .A2(n16876), .B1(n5329), .B2(n16873), .ZN(n4509) );
  NAND4_X1 U5067 ( .A1(n4510), .A2(n4511), .A3(n4512), .A4(n4513), .ZN(n3177)
         );
  AOI222_X1 U5068 ( .A1(n16652), .A2(vis_r14_o[2]), .B1(n16911), .B2(n2620), 
        .C1(n16651), .C2(vis_msp_o[0]), .ZN(n4513) );
  AOI22_X1 U5072 ( .A1(n16902), .A2(vis_psp_o[0]), .B1(n16897), .B2(
        vis_r10_o[2]), .ZN(n4512) );
  AOI222_X1 U5075 ( .A1(n16886), .A2(vis_r12_o[2]), .B1(n16648), .B2(
        vis_r8_o[2]), .C1(n16891), .C2(vis_r9_o[2]), .ZN(n4511) );
  AOI21_X1 U5079 ( .B1(n16650), .B2(vis_r11_o[2]), .A(n4171), .ZN(n4510) );
  NAND2_X1 U5080 ( .A1(n4514), .A2(n4515), .ZN(n4171) );
  AOI221_X1 U5081 ( .B1(n16916), .B2(vis_r4_o[2]), .C1(n16913), .C2(
        vis_r5_o[2]), .A(n4516), .ZN(n4515) );
  OAI22_X1 U5082 ( .A1(n5475), .A2(n16905), .B1(n5194), .B2(n16908), .ZN(n4516) );
  AOI221_X1 U5085 ( .B1(n16877), .B2(vis_r3_o[2]), .C1(n16649), .C2(
        vis_r7_o[2]), .A(n4519), .ZN(n4514) );
  OAI22_X1 U5086 ( .A1(n5499), .A2(n4427), .B1(n5056), .B2(n16885), .ZN(n4519)
         );
  NAND4_X1 U5092 ( .A1(n4520), .A2(n4521), .A3(n4522), .A4(n4523), .ZN(n2246)
         );
  AOI221_X1 U5093 ( .B1(n16916), .B2(vis_r4_o[11]), .C1(n16913), .C2(
        vis_r5_o[11]), .A(n4524), .ZN(n4523) );
  OAI222_X1 U5094 ( .A1(n4831), .A2(n16910), .B1(n5564), .B2(n16907), .C1(
        n5556), .C2(n16904), .ZN(n4524) );
  AOI221_X1 U5097 ( .B1(n16901), .B2(vis_psp_o[9]), .C1(n16899), .C2(
        vis_r10_o[11]), .A(n4525), .ZN(n4522) );
  OAI22_X1 U5098 ( .A1(n5567), .A2(n16894), .B1(n5568), .B2(n16892), .ZN(n4525) );
  AOI221_X1 U5101 ( .B1(n16890), .B2(vis_r9_o[11]), .C1(n16888), .C2(
        vis_r12_o[11]), .A(n4526), .ZN(n4521) );
  OAI22_X1 U5102 ( .A1(n5555), .A2(n16884), .B1(n5558), .B2(n16881), .ZN(n4526) );
  AOI221_X1 U5105 ( .B1(n16880), .B2(vis_r0_o[11]), .C1(n16879), .C2(
        vis_r3_o[11]), .A(n4528), .ZN(n4520) );
  OAI22_X1 U5106 ( .A1(n5565), .A2(n16876), .B1(n5561), .B2(n16873), .ZN(n4528) );
  NAND4_X1 U5109 ( .A1(n4529), .A2(n4530), .A3(n4531), .A4(n4532), .ZN(n2257)
         );
  AOI222_X1 U5110 ( .A1(n16652), .A2(vis_r14_o[3]), .B1(n16911), .B2(n2593), 
        .C1(n16651), .C2(vis_msp_o[1]), .ZN(n4532) );
  AOI22_X1 U5114 ( .A1(n16902), .A2(vis_psp_o[1]), .B1(n16897), .B2(
        vis_r10_o[3]), .ZN(n4531) );
  AOI222_X1 U5117 ( .A1(n16886), .A2(vis_r12_o[3]), .B1(n16648), .B2(
        vis_r8_o[3]), .C1(n16891), .C2(vis_r9_o[3]), .ZN(n4530) );
  AOI21_X1 U5121 ( .B1(n16650), .B2(vis_r11_o[3]), .A(n4069), .ZN(n4529) );
  NAND2_X1 U5122 ( .A1(n4533), .A2(n4534), .ZN(n4069) );
  AOI221_X1 U5123 ( .B1(n16916), .B2(vis_r4_o[3]), .C1(n16913), .C2(
        vis_r5_o[3]), .A(n4535), .ZN(n4534) );
  OAI22_X1 U5124 ( .A1(n5464), .A2(n16905), .B1(n5183), .B2(n16908), .ZN(n4535) );
  AOI221_X1 U5127 ( .B1(n16877), .B2(vis_r3_o[3]), .C1(n16649), .C2(
        vis_r7_o[3]), .A(n4538), .ZN(n4533) );
  OAI22_X1 U5128 ( .A1(n5488), .A2(n4427), .B1(n5028), .B2(n16885), .ZN(n4538)
         );
  NAND4_X1 U5134 ( .A1(n4539), .A2(n4540), .A3(n4541), .A4(n4542), .ZN(n2247)
         );
  AOI221_X1 U5135 ( .B1(n16916), .B2(vis_r4_o[12]), .C1(n16913), .C2(
        vis_r5_o[12]), .A(n4543), .ZN(n4542) );
  OAI222_X1 U5136 ( .A1(n4830), .A2(n16910), .B1(n5192), .B2(n16907), .C1(
        n5473), .C2(n16904), .ZN(n4543) );
  AOI221_X1 U5139 ( .B1(n16901), .B2(vis_psp_o[10]), .C1(n16899), .C2(
        vis_r10_o[12]), .A(n4544), .ZN(n4541) );
  OAI22_X1 U5140 ( .A1(n5301), .A2(n16894), .B1(n5130), .B2(n16892), .ZN(n4544) );
  AOI221_X1 U5143 ( .B1(n16890), .B2(vis_r9_o[12]), .C1(n16888), .C2(
        vis_r12_o[12]), .A(n4545), .ZN(n4540) );
  OAI22_X1 U5144 ( .A1(n5127), .A2(n16884), .B1(n5415), .B2(n16881), .ZN(n4545) );
  AOI221_X1 U5147 ( .B1(n4224), .B2(vis_r0_o[12]), .C1(n16879), .C2(
        vis_r3_o[12]), .A(n4547), .ZN(n4539) );
  OAI22_X1 U5148 ( .A1(n5129), .A2(n16876), .B1(n5328), .B2(n16873), .ZN(n4547) );
  NAND4_X1 U5151 ( .A1(n4548), .A2(n4549), .A3(n4550), .A4(n4551), .ZN(n2578)
         );
  AOI222_X1 U5152 ( .A1(n16652), .A2(vis_r14_o[4]), .B1(n16911), .B2(n2570), 
        .C1(n16651), .C2(vis_msp_o[2]), .ZN(n4551) );
  AOI22_X1 U5156 ( .A1(n16902), .A2(vis_psp_o[2]), .B1(n16897), .B2(
        vis_r10_o[4]), .ZN(n4550) );
  AOI222_X1 U5159 ( .A1(n16886), .A2(vis_r12_o[4]), .B1(n16648), .B2(
        vis_r8_o[4]), .C1(n16891), .C2(vis_r9_o[4]), .ZN(n4549) );
  AOI21_X1 U5163 ( .B1(n16650), .B2(vis_r11_o[4]), .A(n4065), .ZN(n4548) );
  NAND2_X1 U5164 ( .A1(n4552), .A2(n4553), .ZN(n4065) );
  AOI221_X1 U5165 ( .B1(n16915), .B2(vis_r4_o[4]), .C1(n16912), .C2(
        vis_r5_o[4]), .A(n4554), .ZN(n4553) );
  OAI22_X1 U5166 ( .A1(n5463), .A2(n16905), .B1(n5182), .B2(n16908), .ZN(n4554) );
  AOI221_X1 U5169 ( .B1(n16877), .B2(vis_r3_o[4]), .C1(n16649), .C2(
        vis_r7_o[4]), .A(n4557), .ZN(n4552) );
  OAI22_X1 U5170 ( .A1(n5487), .A2(n4427), .B1(n5121), .B2(n16885), .ZN(n4557)
         );
  NAND4_X1 U5176 ( .A1(n4558), .A2(n4559), .A3(n4560), .A4(n4561), .ZN(n2259)
         );
  AOI221_X1 U5177 ( .B1(n16915), .B2(vis_r4_o[13]), .C1(n16912), .C2(
        vis_r5_o[13]), .A(n4562), .ZN(n4561) );
  OAI222_X1 U5178 ( .A1(n4832), .A2(n16910), .B1(n5191), .B2(n16907), .C1(
        n5472), .C2(n16904), .ZN(n4562) );
  AOI221_X1 U5181 ( .B1(n16901), .B2(vis_psp_o[11]), .C1(n16899), .C2(
        vis_r10_o[13]), .A(n4563), .ZN(n4560) );
  OAI22_X1 U5182 ( .A1(n5597), .A2(n16894), .B1(n5598), .B2(n16892), .ZN(n4563) );
  AOI221_X1 U5185 ( .B1(n16890), .B2(vis_r9_o[13]), .C1(n16888), .C2(
        vis_r12_o[13]), .A(n4564), .ZN(n4559) );
  OAI22_X1 U5186 ( .A1(n5132), .A2(n16884), .B1(n5414), .B2(n16881), .ZN(n4564) );
  AOI221_X1 U5189 ( .B1(n4224), .B2(vis_r0_o[13]), .C1(n16879), .C2(
        vis_r3_o[13]), .A(n4566), .ZN(n4558) );
  OAI22_X1 U5190 ( .A1(n5134), .A2(n16876), .B1(n5327), .B2(n16873), .ZN(n4566) );
  INV_X1 U5193 ( .A(n16786), .ZN(n4401) );
  NOR3_X1 U5194 ( .A1(n1670), .A2(n5167), .A3(n1612), .ZN(n4239) );
  AOI21_X1 U5195 ( .B1(n3362), .B2(n4567), .A(n1612), .ZN(n1670) );
  OAI21_X1 U5196 ( .B1(n16856), .B2(n632), .A(n556), .ZN(n4567) );
  NAND2_X1 U5197 ( .A1(n16834), .A2(n16856), .ZN(n556) );
  INV_X1 U5198 ( .A(n604), .ZN(n632) );
  NAND2_X1 U5199 ( .A1(n16834), .A2(n16860), .ZN(n604) );
  NAND2_X1 U5200 ( .A1(n16837), .A2(n16855), .ZN(n3362) );
  NAND4_X1 U5201 ( .A1(n4568), .A2(n4569), .A3(n4570), .A4(n4571), .ZN(n2556)
         );
  AOI222_X1 U5202 ( .A1(n16652), .A2(vis_r14_o[5]), .B1(n16911), .B2(n2539), 
        .C1(n16651), .C2(vis_msp_o[3]), .ZN(n4571) );
  AOI22_X1 U5206 ( .A1(n16902), .A2(vis_psp_o[3]), .B1(n16897), .B2(
        vis_r10_o[5]), .ZN(n4570) );
  AOI222_X1 U5209 ( .A1(n16886), .A2(vis_r12_o[5]), .B1(n16648), .B2(
        vis_r8_o[5]), .C1(n16891), .C2(vis_r9_o[5]), .ZN(n4569) );
  AOI21_X1 U5213 ( .B1(n16650), .B2(vis_r11_o[5]), .A(n4058), .ZN(n4568) );
  NAND2_X1 U5214 ( .A1(n4572), .A2(n4573), .ZN(n4058) );
  AOI221_X1 U5215 ( .B1(n16915), .B2(vis_r4_o[5]), .C1(n16912), .C2(
        vis_r5_o[5]), .A(n4574), .ZN(n4573) );
  OAI22_X1 U5216 ( .A1(n5462), .A2(n16905), .B1(n5181), .B2(n16908), .ZN(n4574) );
  AOI221_X1 U5219 ( .B1(n16877), .B2(vis_r3_o[5]), .C1(n16649), .C2(
        vis_r7_o[5]), .A(n4577), .ZN(n4572) );
  OAI22_X1 U5220 ( .A1(n5486), .A2(n4427), .B1(n5091), .B2(n16885), .ZN(n4577)
         );
  NAND4_X1 U5226 ( .A1(n4578), .A2(n4579), .A3(n4580), .A4(n4581), .ZN(n2196)
         );
  AOI222_X1 U5227 ( .A1(n16652), .A2(vis_r14_o[7]), .B1(n16911), .B2(n2221), 
        .C1(n16651), .C2(vis_msp_o[5]), .ZN(n4581) );
  AOI22_X1 U5234 ( .A1(n16902), .A2(vis_psp_o[5]), .B1(n16897), .B2(
        vis_r10_o[7]), .ZN(n4580) );
  AOI222_X1 U5237 ( .A1(n16886), .A2(vis_r12_o[7]), .B1(n16648), .B2(
        vis_r8_o[7]), .C1(n16891), .C2(vis_r9_o[7]), .ZN(n4579) );
  AOI21_X1 U5242 ( .B1(n16650), .B2(vis_r11_o[7]), .A(n1795), .ZN(n4578) );
  NAND2_X1 U5243 ( .A1(n4582), .A2(n4583), .ZN(n1795) );
  AOI221_X1 U5244 ( .B1(n16915), .B2(vis_r4_o[7]), .C1(n16912), .C2(
        vis_r5_o[7]), .A(n4584), .ZN(n4583) );
  OAI22_X1 U5245 ( .A1(n5452), .A2(n16905), .B1(n5171), .B2(n16908), .ZN(n4584) );
  AOI221_X1 U5248 ( .B1(n16877), .B2(vis_r3_o[7]), .C1(n16649), .C2(
        vis_r7_o[7]), .A(n4587), .ZN(n4582) );
  OAI22_X1 U5249 ( .A1(n5022), .A2(n4427), .B1(n5021), .B2(n16885), .ZN(n4587)
         );
  NAND3_X1 U5258 ( .A1(n16839), .A2(n16859), .A3(n3430), .ZN(n4589) );
  NAND2_X1 U5259 ( .A1(n1805), .A2(n1094), .ZN(n4588) );
  INV_X1 U5260 ( .A(n1023), .ZN(n1094) );
  NAND2_X1 U5261 ( .A1(n16854), .A2(n16867), .ZN(n1023) );
  NAND2_X1 U5262 ( .A1(n16845), .A2(n16838), .ZN(n1603) );
  NAND4_X1 U5264 ( .A1(n4591), .A2(n4592), .A3(n4593), .A4(n4594), .ZN(n3450)
         );
  AOI221_X1 U5265 ( .B1(n16915), .B2(vis_r4_o[23]), .C1(n16912), .C2(
        vis_r5_o[23]), .A(n4595), .ZN(n4594) );
  OAI222_X1 U5266 ( .A1(n4772), .A2(n16910), .B1(n5592), .B2(n16907), .C1(
        n5584), .C2(n16904), .ZN(n4595) );
  AOI221_X1 U5269 ( .B1(n16901), .B2(vis_psp_o[21]), .C1(n16899), .C2(
        vis_r10_o[23]), .A(n4596), .ZN(n4593) );
  OAI22_X1 U5270 ( .A1(n5594), .A2(n16894), .B1(n4970), .B2(n16892), .ZN(n4596) );
  AOI221_X1 U5273 ( .B1(n16890), .B2(vis_r9_o[23]), .C1(n16888), .C2(
        vis_r12_o[23]), .A(n4597), .ZN(n4592) );
  OAI22_X1 U5274 ( .A1(n4983), .A2(n16884), .B1(n5586), .B2(n16881), .ZN(n4597) );
  AOI221_X1 U5277 ( .B1(n4224), .B2(vis_r0_o[23]), .C1(n16879), .C2(
        vis_r3_o[23]), .A(n4599), .ZN(n4591) );
  OAI22_X1 U5278 ( .A1(n4960), .A2(n16876), .B1(n5589), .B2(n16873), .ZN(n4599) );
  OAI22_X1 U5281 ( .A1(n2461), .A2(n4600), .B1(n2462), .B2(n89), .ZN(U189_Z_0)
         );
  INV_X1 U5282 ( .A(n89), .ZN(n4600) );
  NAND4_X1 U5283 ( .A1(n4601), .A2(n4602), .A3(n4603), .A4(n4604), .ZN(n89) );
  AOI221_X1 U5284 ( .B1(n16915), .B2(vis_r4_o[28]), .C1(n16912), .C2(
        vis_r5_o[28]), .A(n4605), .ZN(n4604) );
  OAI222_X1 U5285 ( .A1(n5626), .A2(n16910), .B1(n5170), .B2(n16907), .C1(
        n5451), .C2(n16904), .ZN(n4605) );
  AOI221_X1 U5288 ( .B1(n16901), .B2(vis_psp_o[26]), .C1(n16899), .C2(
        vis_r10_o[28]), .A(n4606), .ZN(n4603) );
  OAI22_X1 U5289 ( .A1(n5285), .A2(n16894), .B1(n4994), .B2(n16892), .ZN(n4606) );
  AOI221_X1 U5292 ( .B1(n16890), .B2(vis_r9_o[28]), .C1(n16888), .C2(
        vis_r12_o[28]), .A(n4607), .ZN(n4602) );
  OAI22_X1 U5293 ( .A1(n4997), .A2(n16884), .B1(n5393), .B2(n16881), .ZN(n4607) );
  AOI221_X1 U5296 ( .B1(n4224), .B2(vis_r0_o[28]), .C1(n16879), .C2(
        vis_r3_o[28]), .A(n4609), .ZN(n4601) );
  OAI22_X1 U5297 ( .A1(n4996), .A2(n16876), .B1(n5306), .B2(n16873), .ZN(n4609) );
  INV_X1 U5301 ( .A(n3534), .ZN(n4610) );
  NAND4_X1 U5302 ( .A1(n4611), .A2(n4612), .A3(n4613), .A4(n4614), .ZN(n3534)
         );
  AOI221_X1 U5303 ( .B1(n16915), .B2(vis_r4_o[31]), .C1(n16912), .C2(
        vis_r5_o[31]), .A(n4615), .ZN(n4614) );
  OAI222_X1 U5304 ( .A1(n4774), .A2(n16910), .B1(n5169), .B2(n16907), .C1(
        n5450), .C2(n16904), .ZN(n4615) );
  AOI221_X1 U5307 ( .B1(n16902), .B2(vis_psp_o[29]), .C1(n16899), .C2(
        vis_r10_o[31]), .A(n4616), .ZN(n4613) );
  OAI22_X1 U5308 ( .A1(n5284), .A2(n16894), .B1(n4969), .B2(n16892), .ZN(n4616) );
  AOI221_X1 U5311 ( .B1(n16890), .B2(vis_r9_o[31]), .C1(n16888), .C2(
        vis_r12_o[31]), .A(n4617), .ZN(n4612) );
  OAI22_X1 U5312 ( .A1(n4981), .A2(n16884), .B1(n5392), .B2(n16881), .ZN(n4617) );
  AOI221_X1 U5315 ( .B1(n16880), .B2(vis_r0_o[31]), .C1(n16879), .C2(
        vis_r3_o[31]), .A(n4619), .ZN(n4611) );
  OAI22_X1 U5316 ( .A1(n4962), .A2(n16876), .B1(n5305), .B2(n16873), .ZN(n4619) );
  OAI22_X1 U5319 ( .A1(n2461), .A2(n4620), .B1(n2462), .B2(n2083), .ZN(
        U180_Z_0) );
  INV_X1 U5320 ( .A(n2083), .ZN(n4620) );
  NAND4_X1 U5321 ( .A1(n4621), .A2(n4622), .A3(n4623), .A4(n4624), .ZN(n2083)
         );
  AOI221_X1 U5322 ( .B1(n16915), .B2(vis_r4_o[30]), .C1(n16912), .C2(
        vis_r5_o[30]), .A(n4625), .ZN(n4624) );
  OAI222_X1 U5323 ( .A1(n4955), .A2(n16910), .B1(n5174), .B2(n16908), .C1(
        n5455), .C2(n16905), .ZN(n4625) );
  AOI221_X1 U5326 ( .B1(n16901), .B2(vis_psp_o[28]), .C1(n16899), .C2(
        vis_r10_o[30]), .A(n4626), .ZN(n4623) );
  OAI22_X1 U5327 ( .A1(n5641), .A2(n16894), .B1(n5642), .B2(n16892), .ZN(n4626) );
  AOI221_X1 U5330 ( .B1(n16891), .B2(vis_r9_o[30]), .C1(n16888), .C2(
        vis_r12_o[30]), .A(n4627), .ZN(n4622) );
  OAI22_X1 U5331 ( .A1(n5080), .A2(n16885), .B1(n5397), .B2(n16881), .ZN(n4627) );
  AOI221_X1 U5334 ( .B1(n4224), .B2(vis_r0_o[30]), .C1(n16879), .C2(
        vis_r3_o[30]), .A(n4629), .ZN(n4621) );
  OAI22_X1 U5335 ( .A1(n5082), .A2(n16876), .B1(n5310), .B2(n16873), .ZN(n4629) );
  OAI22_X1 U5338 ( .A1(n2461), .A2(n4630), .B1(n2462), .B2(n2427), .ZN(
        U175_Z_0) );
  INV_X1 U5339 ( .A(n2427), .ZN(n4630) );
  NAND4_X1 U5340 ( .A1(n4631), .A2(n4632), .A3(n4633), .A4(n4634), .ZN(n2427)
         );
  AOI221_X1 U5341 ( .B1(n16915), .B2(vis_r4_o[27]), .C1(n16912), .C2(
        vis_r5_o[27]), .A(n4635), .ZN(n4634) );
  OAI222_X1 U5342 ( .A1(n4761), .A2(n16909), .B1(n5176), .B2(n16908), .C1(
        n5457), .C2(n16905), .ZN(n4635) );
  AOI221_X1 U5345 ( .B1(n16902), .B2(vis_psp_o[25]), .C1(n16899), .C2(
        vis_r10_o[27]), .A(n4636), .ZN(n4633) );
  OAI22_X1 U5346 ( .A1(n5628), .A2(n16894), .B1(n5629), .B2(n16892), .ZN(n4636) );
  AOI221_X1 U5349 ( .B1(n16891), .B2(vis_r9_o[27]), .C1(n16888), .C2(
        vis_r12_o[27]), .A(n4637), .ZN(n4632) );
  OAI22_X1 U5350 ( .A1(n5111), .A2(n16885), .B1(n5399), .B2(n16881), .ZN(n4637) );
  AOI221_X1 U5353 ( .B1(n4224), .B2(vis_r0_o[27]), .C1(n16879), .C2(
        vis_r3_o[27]), .A(n4639), .ZN(n4631) );
  OAI22_X1 U5354 ( .A1(n5113), .A2(n16876), .B1(n5312), .B2(n16873), .ZN(n4639) );
  OAI22_X1 U5357 ( .A1(n2461), .A2(n4640), .B1(n2462), .B2(n2496), .ZN(
        U163_Z_0) );
  INV_X1 U5358 ( .A(n2496), .ZN(n4640) );
  NAND4_X1 U5359 ( .A1(n4641), .A2(n4642), .A3(n4643), .A4(n4644), .ZN(n2496)
         );
  AOI221_X1 U5360 ( .B1(n16915), .B2(vis_r4_o[24]), .C1(n16912), .C2(
        vis_r5_o[24]), .A(n4645), .ZN(n4644) );
  OAI222_X1 U5361 ( .A1(n4971), .A2(n16909), .B1(n5179), .B2(n16907), .C1(
        n5460), .C2(n16904), .ZN(n4645) );
  AOI221_X1 U5364 ( .B1(n16901), .B2(vis_psp_o[22]), .C1(n16899), .C2(
        vis_r10_o[24]), .A(n4646), .ZN(n4643) );
  OAI22_X1 U5365 ( .A1(n5645), .A2(n16894), .B1(n5646), .B2(n16892), .ZN(n4646) );
  AOI221_X1 U5368 ( .B1(n16890), .B2(vis_r9_o[24]), .C1(n16888), .C2(
        vis_r12_o[24]), .A(n4647), .ZN(n4642) );
  OAI22_X1 U5369 ( .A1(n4982), .A2(n16884), .B1(n5402), .B2(n16881), .ZN(n4647) );
  AOI221_X1 U5372 ( .B1(n4224), .B2(vis_r0_o[24]), .C1(n16879), .C2(
        vis_r3_o[24]), .A(n4649), .ZN(n4641) );
  OAI22_X1 U5373 ( .A1(n4972), .A2(n16876), .B1(n5315), .B2(n16873), .ZN(n4649) );
  OAI22_X1 U5376 ( .A1(n2462), .A2(n1755), .B1(n2461), .B2(n4650), .ZN(
        U158_Z_0) );
  INV_X1 U5377 ( .A(n1755), .ZN(n4650) );
  INV_X1 U5378 ( .A(n2492), .ZN(n2461) );
  OAI21_X1 U5379 ( .B1(n16991), .B2(n3180), .A(n4651), .ZN(n2492) );
  NAND4_X1 U5381 ( .A1(n4652), .A2(n4653), .A3(n4654), .A4(n4655), .ZN(n1755)
         );
  AOI221_X1 U5382 ( .B1(n16915), .B2(vis_r4_o[29]), .C1(n16912), .C2(
        vis_r5_o[29]), .A(n4656), .ZN(n4655) );
  OAI222_X1 U5383 ( .A1(n4773), .A2(n16909), .B1(n5175), .B2(n16906), .C1(
        n5456), .C2(n16903), .ZN(n4656) );
  NAND2_X1 U5386 ( .A1(n4660), .A2(n4661), .ZN(n4211) );
  AOI221_X1 U5391 ( .B1(n16900), .B2(vis_psp_o[27]), .C1(n16897), .C2(
        vis_r10_o[29]), .A(n4664), .ZN(n4654) );
  OAI22_X1 U5392 ( .A1(n5289), .A2(n16894), .B1(n5078), .B2(n16892), .ZN(n4664) );
  NOR2_X1 U5397 ( .A1(n3489), .A2(n5545), .ZN(n4658) );
  AOI221_X1 U5401 ( .B1(n16889), .B2(vis_r9_o[29]), .C1(n16886), .C2(
        vis_r12_o[29]), .A(n4666), .ZN(n4653) );
  OAI22_X1 U5402 ( .A1(n5075), .A2(n16883), .B1(n5398), .B2(n16881), .ZN(n4666) );
  NOR2_X1 U5407 ( .A1(n5544), .A2(n5259), .ZN(n4660) );
  NOR2_X1 U5410 ( .A1(n1353), .A2(n5004), .ZN(n4662) );
  AOI221_X1 U5411 ( .B1(n4224), .B2(vis_r0_o[29]), .C1(n16877), .C2(
        vis_r3_o[29]), .A(n4668), .ZN(n4652) );
  OAI22_X1 U5412 ( .A1(n5077), .A2(n16876), .B1(n5311), .B2(n16873), .ZN(n4668) );
  NOR2_X1 U5414 ( .A1(n3493), .A2(n5544), .ZN(n4665) );
  NOR2_X1 U5416 ( .A1(n3496), .A2(n5259), .ZN(n4659) );
  NOR2_X1 U5419 ( .A1(n5004), .A2(n5545), .ZN(n4661) );
  INV_X1 U5421 ( .A(n4427), .ZN(n4224) );
  NOR2_X1 U5423 ( .A1(n3493), .A2(n3496), .ZN(n4657) );
  NOR2_X1 U5426 ( .A1(n1353), .A2(n3489), .ZN(n4663) );
  INV_X1 U5429 ( .A(n2493), .ZN(n2462) );
  OAI21_X1 U5430 ( .B1(n4669), .B2(n16990), .A(n4651), .ZN(n2493) );
  AOI21_X1 U5431 ( .B1(n16990), .B2(n4669), .A(n4670), .ZN(n4651) );
  NOR3_X1 U5432 ( .A1(n4669), .A2(n16988), .A3(n16990), .ZN(n4670) );
  OAI21_X1 U5434 ( .B1(n4671), .B2(n4672), .A(n1697), .ZN(n3180) );
  OAI222_X1 U5435 ( .A1(n1784), .A2(n673), .B1(n16851), .B2(n4673), .C1(n16833), .C2(n758), .ZN(n4672) );
  INV_X1 U5436 ( .A(n515), .ZN(n758) );
  NOR2_X1 U5437 ( .A1(n16805), .A2(n16825), .ZN(n515) );
  NOR4_X1 U5438 ( .A1(n3506), .A2(n2042), .A3(n529), .A4(n4674), .ZN(n4673) );
  NOR3_X1 U5439 ( .A1(n617), .A2(n16828), .A3(n16839), .ZN(n4674) );
  INV_X1 U5441 ( .A(n666), .ZN(n2042) );
  NAND2_X1 U5442 ( .A1(n16855), .A2(n16831), .ZN(n666) );
  INV_X1 U5443 ( .A(n1103), .ZN(n3506) );
  NAND2_X1 U5444 ( .A1(n16826), .A2(n16831), .ZN(n1103) );
  OAI221_X1 U5446 ( .B1(n617), .B2(n1278), .C1(n16824), .C2(n16867), .A(n4675), 
        .ZN(n4671) );
  NAND3_X1 U5447 ( .A1(n1805), .A2(n991), .A3(n1042), .ZN(n4675) );
  INV_X1 U5448 ( .A(n641), .ZN(n1042) );
  NAND2_X1 U5449 ( .A1(n16856), .A2(n16849), .ZN(n641) );
  INV_X1 U5452 ( .A(n1579), .ZN(n1805) );
  NAND2_X1 U5453 ( .A1(n16837), .A2(n16860), .ZN(n1579) );
  NAND2_X1 U5454 ( .A1(n565), .A2(n16831), .ZN(n1278) );
  OAI211_X1 U5456 ( .C1(n16859), .C2(n890), .A(n4677), .B(n4678), .ZN(n4676)
         );
  AOI21_X1 U5457 ( .B1(n667), .B2(n1564), .A(n4679), .ZN(n4678) );
  OAI33_X1 U5458 ( .A1(n1518), .A2(n16868), .A3(n16866), .B1(n16867), .B2(
        n16823), .B3(n4680), .ZN(n4679) );
  AOI21_X1 U5459 ( .B1(n16862), .B2(n16842), .A(n501), .ZN(n4680) );
  INV_X1 U5460 ( .A(n617), .ZN(n501) );
  NAND2_X1 U5462 ( .A1(n2646), .A2(n16860), .ZN(n1518) );
  INV_X1 U5463 ( .A(n1233), .ZN(n2646) );
  NAND2_X1 U5464 ( .A1(n16842), .A2(n16839), .ZN(n1233) );
  INV_X1 U5465 ( .A(n1580), .ZN(n1564) );
  NAND2_X1 U5466 ( .A1(n16851), .A2(n16843), .ZN(n1580) );
  INV_X1 U5467 ( .A(n1706), .ZN(n667) );
  NAND2_X1 U5468 ( .A1(n16830), .A2(n16839), .ZN(n1706) );
  INV_X1 U5469 ( .A(n1705), .ZN(n4677) );
  OAI222_X1 U5470 ( .A1(n1104), .A2(n849), .B1(n745), .B2(n568), .C1(n16868), 
        .C2(n1517), .ZN(n1705) );
  NAND2_X1 U5471 ( .A1(n16837), .A2(n16690), .ZN(n568) );
  NAND2_X1 U5472 ( .A1(n16866), .A2(n16839), .ZN(n849) );
  NAND2_X1 U5473 ( .A1(n565), .A2(n17096), .ZN(n890) );
  OR2_X1 U5475 ( .A1(n2732), .A2(n2716), .ZN(n4669) );
  NOR2_X1 U5476 ( .A1(n2543), .A2(n5254), .ZN(n2716) );
  NAND4_X1 U5477 ( .A1(n3430), .A2(n16833), .A3(n16826), .A4(n1697), .ZN(n2543) );
  INV_X1 U5478 ( .A(n1104), .ZN(n3430) );
  NAND2_X1 U5481 ( .A1(n3164), .A2(n1723), .ZN(n2719) );
  INV_X1 U5482 ( .A(n3186), .ZN(n3164) );
  NAND3_X1 U5483 ( .A1(n1095), .A2(n1697), .A3(n483), .ZN(n3186) );
  INV_X1 U5485 ( .A(n1784), .ZN(n1095) );
  NAND2_X1 U5486 ( .A1(n16854), .A2(n16843), .ZN(n1784) );
  OAI22_X1 U5487 ( .A1(n4959), .A2(n4681), .B1(n4682), .B2(n4683), .ZN(
        U144_Z_0) );
  AOI21_X1 U5488 ( .B1(n4684), .B2(n16798), .A(n4685), .ZN(n4682) );
  OAI21_X1 U5489 ( .B1(n16816), .B2(n4686), .A(n782), .ZN(n4684) );
  OAI22_X1 U5490 ( .A1(n4978), .A2(n4681), .B1(n4687), .B2(n4683), .ZN(
        U134_Z_0) );
  AOI211_X1 U5491 ( .C1(n4688), .C2(n451), .A(n4689), .B(n4685), .ZN(n4687) );
  OAI22_X1 U5492 ( .A1(n16794), .A2(n4690), .B1(n17099), .B2(n4691), .ZN(n4689) );
  OAI22_X1 U5493 ( .A1(n5004), .A2(n1713), .B1(n4692), .B2(n1715), .ZN(
        U122_Z_0) );
  AOI211_X1 U5494 ( .C1(n597), .C2(n486), .A(n4693), .B(n4694), .ZN(n4692) );
  OAI22_X1 U5495 ( .A1(n4695), .A2(n1307), .B1(n4967), .B2(n1719), .ZN(n4694)
         );
  NAND2_X1 U5496 ( .A1(n473), .A2(n16815), .ZN(n1719) );
  AOI221_X1 U5497 ( .B1(n4696), .B2(n1286), .C1(n4697), .C2(n664), .A(n4698), 
        .ZN(n4695) );
  OAI22_X1 U5498 ( .A1(n5003), .A2(n486), .B1(n4699), .B2(n437), .ZN(n4698) );
  NAND2_X1 U5499 ( .A1(n5258), .A2(n4697), .ZN(n664) );
  INV_X1 U5500 ( .A(n1294), .ZN(n4697) );
  OAI221_X1 U5501 ( .B1(n16794), .B2(n1721), .C1(n16801), .C2(n819), .A(n1720), 
        .ZN(n4693) );
  NOR3_X1 U5502 ( .A1(n483), .A2(n1478), .A3(n896), .ZN(n1720) );
  INV_X1 U5503 ( .A(n1170), .ZN(n896) );
  NOR2_X1 U5504 ( .A1(n784), .A2(n493), .ZN(n1170) );
  NOR2_X1 U5505 ( .A1(n640), .A2(n16845), .ZN(n493) );
  INV_X1 U5506 ( .A(n4318), .ZN(n784) );
  NAND2_X1 U5507 ( .A1(n608), .A2(n16843), .ZN(n4318) );
  INV_X1 U5508 ( .A(n745), .ZN(n608) );
  OAI21_X1 U5510 ( .B1(n822), .B2(n16817), .A(n1728), .ZN(n1721) );
  NAND2_X1 U5511 ( .A1(n1594), .A2(n1198), .ZN(n1728) );
  INV_X1 U5514 ( .A(n1715), .ZN(n1713) );
  NAND2_X1 U5515 ( .A1(n17124), .A2(n4700), .ZN(n1715) );
  NAND4_X1 U5516 ( .A1(n4701), .A2(n4702), .A3(n4703), .A4(n4704), .ZN(n4700)
         );
  NOR4_X1 U5517 ( .A1(n741), .A2(n495), .A3(n1302), .A4(n4705), .ZN(n4704) );
  NOR4_X1 U5518 ( .A1(n16828), .A2(n16821), .A3(n918), .A4(n1307), .ZN(n4705)
         );
  INV_X1 U5519 ( .A(n614), .ZN(n1307) );
  NOR2_X1 U5520 ( .A1(n4590), .A2(n16826), .ZN(n614) );
  NAND2_X1 U5521 ( .A1(n16870), .A2(n16851), .ZN(n4590) );
  NOR2_X1 U5523 ( .A1(n3528), .A2(n1467), .ZN(n1302) );
  INV_X1 U5524 ( .A(n911), .ZN(n1467) );
  NAND3_X1 U5525 ( .A1(n3313), .A2(vis_pc_o[2]), .A3(n5230), .ZN(n911) );
  NOR4_X1 U5528 ( .A1(n610), .A2(n640), .A3(n16826), .A4(n16853), .ZN(n495) );
  AOI222_X1 U5530 ( .A1(n486), .A2(n2774), .B1(n776), .B2(n16671), .C1(n437), 
        .C2(n1723), .ZN(n4708) );
  AOI22_X1 U5535 ( .A1(n455), .A2(n2731), .B1(n768), .B2(n2865), .ZN(n4707) );
  AOI22_X1 U5538 ( .A1(n1294), .A2(n2819), .B1(n1286), .B2(n2827), .ZN(n4706)
         );
  NAND2_X1 U5541 ( .A1(n5257), .A2(n1976), .ZN(n1294) );
  INV_X1 U5542 ( .A(n1286), .ZN(n1976) );
  NAND2_X1 U5543 ( .A1(n5256), .A2(n4696), .ZN(n1286) );
  INV_X1 U5544 ( .A(n768), .ZN(n4696) );
  NAND2_X1 U5545 ( .A1(n4699), .A2(n16810), .ZN(n768) );
  INV_X1 U5546 ( .A(n776), .ZN(n4699) );
  NAND2_X1 U5547 ( .A1(n5254), .A2(n1974), .ZN(n776) );
  INV_X1 U5548 ( .A(n437), .ZN(n1974) );
  NAND2_X1 U5549 ( .A1(n5253), .A2(n1975), .ZN(n437) );
  INV_X1 U5550 ( .A(n455), .ZN(n1975) );
  NAND2_X1 U5551 ( .A1(n5003), .A2(n5162), .ZN(n455) );
  INV_X1 U5552 ( .A(n619), .ZN(n741) );
  NAND2_X1 U5553 ( .A1(n1478), .A2(n16849), .ZN(n619) );
  INV_X1 U5554 ( .A(n694), .ZN(n1478) );
  NAND2_X1 U5555 ( .A1(n527), .A2(n16860), .ZN(n694) );
  AOI222_X1 U5556 ( .A1(n4709), .A2(n4710), .B1(n4711), .B2(n1265), .C1(n4712), 
        .C2(n589), .ZN(n4703) );
  NOR2_X1 U5557 ( .A1(n16837), .A2(n16848), .ZN(n4712) );
  INV_X1 U5558 ( .A(n1908), .ZN(n1265) );
  NAND3_X1 U5559 ( .A1(n16811), .A2(n16819), .A3(n732), .ZN(n1908) );
  INV_X1 U5560 ( .A(n819), .ZN(n732) );
  AOI21_X1 U5562 ( .B1(n16803), .B2(n1562), .A(n503), .ZN(n4711) );
  NAND2_X1 U5563 ( .A1(n16816), .A2(n16733), .ZN(n1562) );
  NAND2_X1 U5564 ( .A1(n1517), .A2(n1303), .ZN(n4710) );
  NAND2_X1 U5565 ( .A1(n526), .A2(n16867), .ZN(n1303) );
  NAND2_X1 U5566 ( .A1(n16866), .A2(n16838), .ZN(n1517) );
  INV_X1 U5567 ( .A(n514), .ZN(n4709) );
  NAND2_X1 U5568 ( .A1(n592), .A2(n16870), .ZN(n514) );
  AOI222_X1 U5569 ( .A1(n333), .A2(n4713), .B1(n16814), .B2(n4714), .C1(n4715), 
        .C2(n16821), .ZN(n4702) );
  INV_X1 U5570 ( .A(n3528), .ZN(n4715) );
  NAND2_X1 U5571 ( .A1(n195), .A2(n527), .ZN(n3528) );
  OAI33_X1 U5576 ( .A1(n4716), .A2(n1920), .A3(n583), .B1(n4717), .B2(n659), 
        .B3(n1928), .ZN(n4714) );
  NAND2_X1 U5577 ( .A1(n16725), .A2(n16686), .ZN(n1928) );
  NAND3_X1 U5579 ( .A1(n440), .A2(n505), .A3(n721), .ZN(n4717) );
  INV_X1 U5580 ( .A(n469), .ZN(n505) );
  INV_X1 U5581 ( .A(n892), .ZN(n440) );
  NAND3_X1 U5582 ( .A1(n708), .A2(n16819), .A3(n821), .ZN(n892) );
  INV_X1 U5583 ( .A(n1552), .ZN(n821) );
  NAND2_X1 U5584 ( .A1(n504), .A2(n17099), .ZN(n583) );
  NOR2_X1 U5585 ( .A1(n669), .A2(n5244), .ZN(n504) );
  NAND2_X1 U5586 ( .A1(n16800), .A2(n16674), .ZN(n669) );
  NAND2_X1 U5588 ( .A1(n476), .A2(n731), .ZN(n4716) );
  INV_X1 U5589 ( .A(n443), .ZN(n476) );
  NAND2_X1 U5592 ( .A1(n16804), .A2(n16820), .ZN(n579) );
  NAND2_X1 U5594 ( .A1(n16871), .A2(n16683), .ZN(n1198) );
  INV_X1 U5595 ( .A(n479), .ZN(n4713) );
  NAND2_X1 U5596 ( .A1(n1492), .A2(n16819), .ZN(n479) );
  INV_X1 U5597 ( .A(n725), .ZN(n1492) );
  NAND2_X1 U5598 ( .A1(n475), .A2(n16802), .ZN(n725) );
  INV_X1 U5599 ( .A(n932), .ZN(n333) );
  NAND2_X1 U5600 ( .A1(n16812), .A2(n791), .ZN(n932) );
  INV_X1 U5601 ( .A(n1261), .ZN(n791) );
  AOI221_X1 U5602 ( .B1(n1263), .B2(n16734), .C1(n506), .C2(n526), .A(n1883), 
        .ZN(n4701) );
  OAI21_X1 U5603 ( .B1(n650), .B2(n4718), .A(n1957), .ZN(n1883) );
  NAND2_X1 U5604 ( .A1(n17096), .A2(n16843), .ZN(n1957) );
  NAND2_X1 U5605 ( .A1(n997), .A2(n16831), .ZN(n4718) );
  INV_X1 U5606 ( .A(n653), .ZN(n997) );
  NAND2_X1 U5611 ( .A1(n16820), .A2(n16843), .ZN(n1882) );
  INV_X1 U5616 ( .A(n1465), .ZN(n506) );
  NAND2_X1 U5617 ( .A1(n589), .A2(n16831), .ZN(n1465) );
  INV_X1 U5618 ( .A(n696), .ZN(n589) );
  NOR3_X1 U5619 ( .A1(n851), .A2(n16839), .A3(n594), .ZN(n1263) );
  NAND4_X1 U5620 ( .A1(n483), .A2(n1468), .A3(n16803), .A4(n16851), .ZN(n594)
         );
  NAND2_X1 U5622 ( .A1(n16870), .A2(n16826), .ZN(n945) );
  OAI22_X1 U5625 ( .A1(n5036), .A2(n4681), .B1(n4719), .B2(n4683), .ZN(
        U121_Z_0) );
  AOI211_X1 U5626 ( .C1(n4688), .C2(n461), .A(n4720), .B(n4721), .ZN(n4719) );
  OAI221_X1 U5627 ( .B1(n16796), .B2(n4691), .C1(n5243), .C2(n4690), .A(n4722), 
        .ZN(n4720) );
  NAND4_X1 U5628 ( .A1(n16814), .A2(n1468), .A3(n592), .A4(n16683), .ZN(n4722)
         );
  OAI22_X1 U5629 ( .A1(n5252), .A2(n4681), .B1(n4723), .B2(n4683), .ZN(
        U105_Z_0) );
  AOI211_X1 U5630 ( .C1(n4688), .C2(n454), .A(n4724), .B(n4685), .ZN(n4723) );
  NAND4_X1 U5631 ( .A1(n4725), .A2(n755), .A3(n4726), .A4(n4727), .ZN(n4685)
         );
  AOI21_X1 U5632 ( .B1(n1468), .B2(n16683), .A(n4721), .ZN(n4727) );
  OAI221_X1 U5633 ( .B1(n4728), .B2(n4686), .C1(n4729), .C2(n1920), .A(n4730), 
        .ZN(n4721) );
  OR4_X1 U5634 ( .A1(n451), .A2(n461), .A3(n782), .A4(n16794), .ZN(n4730) );
  AOI21_X1 U5637 ( .B1(n731), .B2(n16686), .A(n16813), .ZN(n4728) );
  NOR2_X1 U5638 ( .A1(n16725), .A2(n16811), .ZN(n1468) );
  OAI21_X1 U5639 ( .B1(n16851), .B2(n16734), .A(n16805), .ZN(n4726) );
  OAI21_X1 U5640 ( .B1(n16796), .B2(n16807), .A(n630), .ZN(n4725) );
  OAI22_X1 U5641 ( .A1(n5244), .A2(n4690), .B1(n16816), .B2(n4691), .ZN(n4724)
         );
  OAI221_X1 U5642 ( .B1(n1547), .B2(n16659), .C1(n16811), .C2(n16802), .A(n592), .ZN(n4691) );
  NOR2_X1 U5643 ( .A1(n16802), .A2(n16807), .ZN(n1547) );
  OAI21_X1 U5644 ( .B1(n4731), .B2(n4732), .A(n592), .ZN(n4690) );
  OAI33_X1 U5645 ( .A1(n16683), .A2(n16802), .A3(n16725), .B1(n16683), .B2(
        n16795), .B3(n16659), .ZN(n4732) );
  NAND2_X1 U5646 ( .A1(n4733), .A2(n1552), .ZN(n4731) );
  NAND2_X1 U5647 ( .A1(n16802), .A2(n16683), .ZN(n1552) );
  NAND3_X1 U5648 ( .A1(n16657), .A2(n16683), .A3(n630), .ZN(n4733) );
  INV_X1 U5649 ( .A(n1920), .ZN(n630) );
  NAND2_X1 U5650 ( .A1(n16659), .A2(n16725), .ZN(n1920) );
  OAI21_X1 U5653 ( .B1(n782), .B2(n16734), .A(n4686), .ZN(n4688) );
  NAND4_X1 U5654 ( .A1(n16807), .A2(n16811), .A3(n2672), .A4(n16795), .ZN(
        n4686) );
  INV_X1 U5655 ( .A(n4729), .ZN(n2672) );
  NAND2_X1 U5656 ( .A1(n592), .A2(n16802), .ZN(n4729) );
  NAND2_X1 U5661 ( .A1(n16849), .A2(n16805), .ZN(n782) );
  INV_X1 U5663 ( .A(n4683), .ZN(n4681) );
  OAI21_X1 U5664 ( .B1(n4734), .B2(n4735), .A(n17124), .ZN(n4683) );
  OAI221_X1 U5665 ( .B1(n16867), .B2(n692), .C1(n1519), .C2(n696), .A(n488), 
        .ZN(n4735) );
  INV_X1 U5666 ( .A(n4736), .ZN(n488) );
  OAI211_X1 U5667 ( .C1(n1261), .C2(n1267), .A(n1953), .B(n4737), .ZN(n4736)
         );
  NOR2_X1 U5668 ( .A1(n1220), .A2(n4738), .ZN(n4737) );
  NOR4_X1 U5669 ( .A1(n721), .A2(n17098), .A3(n1297), .A4(n469), .ZN(n4738) );
  NAND2_X1 U5670 ( .A1(n16816), .A2(n16657), .ZN(n469) );
  INV_X1 U5671 ( .A(n1021), .ZN(n721) );
  NAND2_X1 U5672 ( .A1(n16801), .A2(n16798), .ZN(n1021) );
  NOR2_X1 U5674 ( .A1(n478), .A2(n16811), .ZN(n1220) );
  AOI21_X1 U5676 ( .B1(n550), .B2(n730), .A(n1471), .ZN(n1953) );
  INV_X1 U5677 ( .A(n738), .ZN(n1471) );
  NAND2_X1 U5678 ( .A1(n799), .A2(n753), .ZN(n738) );
  NAND4_X1 U5679 ( .A1(vis_pc_o[28]), .A2(vis_pc_o[30]), .A3(n2599), .A4(n4739), .ZN(n753) );
  NOR3_X1 U5680 ( .A1(n4843), .A2(n4817), .A3(n4822), .ZN(n4739) );
  NAND4_X1 U5681 ( .A1(n4382), .A2(n191), .A3(n4348), .A4(n170), .ZN(n2599) );
  NOR2_X1 U5683 ( .A1(vis_ipsr_o[5]), .A2(vis_ipsr_o[4]), .ZN(n4348) );
  NOR2_X1 U5685 ( .A1(vis_ipsr_o[2]), .A2(vis_ipsr_o[0]), .ZN(n4382) );
  INV_X1 U5688 ( .A(n755), .ZN(n799) );
  NAND2_X1 U5689 ( .A1(n17097), .A2(n16821), .ZN(n755) );
  INV_X1 U5691 ( .A(n1297), .ZN(n730) );
  NAND2_X1 U5692 ( .A1(n708), .A2(n16804), .ZN(n1297) );
  INV_X1 U5693 ( .A(n582), .ZN(n550) );
  NAND2_X1 U5694 ( .A1(n16796), .A2(n16817), .ZN(n582) );
  NAND2_X1 U5695 ( .A1(n4974), .A2(n16804), .ZN(n1267) );
  NAND2_X1 U5698 ( .A1(n16830), .A2(n16805), .ZN(n692) );
  INV_X1 U5699 ( .A(n16806), .ZN(n797) );
  OAI221_X1 U5702 ( .B1(n4740), .B2(n503), .C1(n16811), .C2(n941), .A(n4741), 
        .ZN(n4734) );
  AOI22_X1 U5703 ( .A1(n4742), .A2(n475), .B1(n4743), .B2(n16816), .ZN(n4741)
         );
  INV_X1 U5704 ( .A(n497), .ZN(n4743) );
  NAND2_X1 U5705 ( .A1(n16797), .A2(n1540), .ZN(n497) );
  INV_X1 U5706 ( .A(n580), .ZN(n1540) );
  NAND2_X1 U5707 ( .A1(n708), .A2(n16812), .ZN(n580) );
  NAND2_X1 U5709 ( .A1(n16871), .A2(n16659), .ZN(n1228) );
  AOI21_X1 U5712 ( .B1(n729), .B2(n16799), .A(n16870), .ZN(n4742) );
  INV_X1 U5713 ( .A(n625), .ZN(n729) );
  NAND2_X1 U5714 ( .A1(n16812), .A2(n16807), .ZN(n625) );
  NOR3_X1 U5716 ( .A1(n4744), .A2(n629), .A3(n4745), .ZN(n4740) );
  NOR3_X1 U5717 ( .A1(n329), .A2(n16803), .A3(n16813), .ZN(n4745) );
  NAND2_X1 U5719 ( .A1(n16871), .A2(n16725), .ZN(n329) );
  INV_X1 U5721 ( .A(n1486), .ZN(n629) );
  NAND2_X1 U5722 ( .A1(n822), .A2(n16803), .ZN(n1486) );
  OAI22_X1 U5723 ( .A1(n731), .A2(n1261), .B1(n941), .B2(n17098), .ZN(n4744)
         );
  NAND2_X1 U5725 ( .A1(n16812), .A2(n822), .ZN(n941) );
  INV_X1 U5726 ( .A(n1594), .ZN(n822) );
  NAND2_X1 U5727 ( .A1(n16795), .A2(n16871), .ZN(n1594) );
  NAND2_X1 U5728 ( .A1(n16807), .A2(n16871), .ZN(n1261) );
  NAND2_X1 U5731 ( .A1(n16657), .A2(n16817), .ZN(n1963) );
  DFFR_X1 Nbm2z4_reg ( .D(n16735), .CK(hclk), .RN(n17189), .Q(n194), .QN(n5034) );
  DFFR_X2 Ypi3z4_reg ( .D(n5654), .CK(hclk), .RN(n17195), .Q(sys_reset_req_o), 
        .QN(n4746) );
  DFFS_X1 F2o2z4_reg ( .D(n5736), .CK(hclk), .SN(n17191), .Q(sub_2068_A_0_), 
        .QN(n260) );
  DFFS_X1 Z8b3z4_reg ( .D(n5730), .CK(hclk), .SN(n17165), .Q(sub_2068_A_6_), 
        .QN(n300) );
  DFFS_X1 W0b3z4_reg ( .D(n5733), .CK(hclk), .SN(n17173), .Q(sub_2068_A_3_), 
        .QN(n306) );
  DFFS_X1 Qxa3z4_reg ( .D(n5731), .CK(hclk), .SN(n17143), .Q(sub_2068_A_5_), 
        .QN(n302) );
  DFFS_X1 M2b3z4_reg ( .D(n5734), .CK(hclk), .SN(n17173), .Q(sub_2068_A_2_), 
        .QN(n308) );
  DFFS_X1 Gza3z4_reg ( .D(n5732), .CK(hclk), .SN(n17173), .Q(sub_2068_A_4_), 
        .QN(n304) );
  DFFS_X1 C4b3z4_reg ( .D(n5735), .CK(hclk), .SN(n17173), .Q(sub_2068_A_1_), 
        .QN(n310) );
  DFFS_X1 Dhb3z4_reg ( .D(n5729), .CK(hclk), .SN(n17139), .Q(sub_2068_A_7_), 
        .QN(n298) );
  DFFS_X1 M5f3z4_reg ( .D(n5728), .CK(hclk), .SN(n17157), .Q(sub_2068_A_8_), 
        .QN(n296) );
  DFFS_X1 Aze3z4_reg ( .D(n5727), .CK(hclk), .SN(n17192), .Q(sub_2068_A_9_), 
        .QN(n294) );
  DFFS_X1 Zva3z4_reg ( .D(n5726), .CK(hclk), .SN(n17173), .Q(sub_2068_A_10_), 
        .QN(n292) );
  DFFS_X1 Jca3z4_reg ( .D(n5653), .CK(hclk), .SN(n17165), .QN(n262) );
  DFFS_X1 She3z4_reg ( .D(n5725), .CK(hclk), .SN(n17173), .Q(sub_2068_A_11_), 
        .QN(n290) );
  DFFS_X1 Iua3z4_reg ( .D(n5724), .CK(hclk), .SN(n17173), .Q(sub_2068_A_12_), 
        .QN(n288) );
  DFFS_X1 K7g3z4_reg ( .D(n5723), .CK(hclk), .SN(n17173), .Q(sub_2068_A_13_), 
        .QN(n286) );
  DFFS_X1 Rsa3z4_reg ( .D(n5722), .CK(hclk), .SN(n17157), .Q(sub_2068_A_14_), 
        .QN(n284) );
  DFFS_X1 Ara3z4_reg ( .D(n5721), .CK(hclk), .SN(n17186), .Q(sub_2068_A_15_), 
        .QN(n282) );
  DFFS_X1 Xeo2z4_reg ( .D(n5720), .CK(hclk), .SN(n17191), .Q(sub_2068_A_16_), 
        .QN(n280) );
  DFFS_X1 S3i3z4_reg ( .D(n5719), .CK(hclk), .SN(n17195), .Q(sub_2068_A_17_), 
        .QN(n278) );
  DFFS_X1 O0o2z4_reg ( .D(n5718), .CK(hclk), .SN(n17158), .Q(sub_2068_A_18_), 
        .QN(n276) );
  DFFS_X1 Jpa3z4_reg ( .D(n5717), .CK(hclk), .SN(n17195), .Q(sub_2068_A_19_), 
        .QN(n274) );
  DFFS_X1 Z2h3z4_reg ( .D(n5716), .CK(hclk), .SN(n17173), .Q(sub_2068_A_20_), 
        .QN(n272) );
  DFFS_X1 Ogo2z4_reg ( .D(n5715), .CK(hclk), .SN(n17172), .Q(sub_2068_A_21_), 
        .QN(n270) );
  DFFS_X1 Ddi3z4_reg ( .D(n5714), .CK(hclk), .SN(n17155), .Q(sub_2068_A_22_), 
        .QN(n268) );
  DFFS_X1 Uei3z4_reg ( .D(n5713), .CK(hclk), .SN(n17189), .Q(sub_2068_A_23_), 
        .QN(n264) );
  DFFS_X1 Ufy2z4_reg ( .D(n14432), .CK(hclk), .SN(n17151), .QN(n370) );
  DFFS_X1 T1y2z4_reg ( .D(n14934), .CK(hclk), .SN(n17155), .QN(n1319) );
  DFFS_X1 Fey2z4_reg ( .D(n5755), .CK(hclk), .SN(n17155), .QN(n335) );
  DFFS_X1 Y7y2z4_reg ( .D(n5760), .CK(hclk), .SN(n17139), .QN(n6) );
  DFFS_X1 I3y2z4_reg ( .D(n5763), .CK(hclk), .SN(n17139), .QN(n9) );
  DFFS_X1 Bdm2z4_reg ( .D(n5756), .CK(hclk), .SN(n17140), .QN(n2) );
  DFFS_X1 K6y2z4_reg ( .D(n5761), .CK(hclk), .SN(n17141), .QN(n7) );
  DFFS_X1 W4y2z4_reg ( .D(n5762), .CK(hclk), .SN(n17140), .QN(n8) );
  DFFS_X1 M9y2z4_reg ( .D(n5759), .CK(hclk), .SN(n17140), .QN(n5) );
  DFFS_X1 Bby2z4_reg ( .D(n5758), .CK(hclk), .SN(n17140), .QN(n4) );
  DFFS_X1 Qcy2z4_reg ( .D(n5757), .CK(hclk), .SN(n17139), .QN(n3) );
  DFFS_X1 Owq2z4_reg ( .D(n5765), .CK(hclk), .SN(n17154), .Q(n4806), .QN(n164)
         );
  DFFS_X1 Lbn2z4_reg ( .D(n5767), .CK(hclk), .SN(n17155), .Q(n4804), .QN(n175)
         );
  DFFS_X1 G0w2z4_reg ( .D(n5691), .CK(hclk), .SN(n17156), .Q(vis_ipsr_o[1]), 
        .QN(n191) );
  DFFS_X1 R1w2z4_reg ( .D(n5692), .CK(hclk), .SN(n17193), .Q(vis_ipsr_o[0]), 
        .QN(n186) );
  DFFR_X1 I6w2z4_reg ( .D(n5827), .CK(hclk), .RN(n17189), .QN(n184) );
  DFFR_X1 Uic3z4_reg ( .D(n5699), .CK(hclk), .RN(n17133), .Q(n4799), .QN(n3010) );
  DFFR_X1 Pab3z4_reg ( .D(U791_Z_0), .CK(hclk), .RN(n17135), .Q(n4753), .QN(
        n1885) );
  DFFR_X1 Fed3z4_reg ( .D(U763_Z_0), .CK(hclk), .RN(n17137), .Q(n4752), .QN(
        n1896) );
  DFFR_X1 W5c3z4_reg ( .D(n13907), .CK(hclk), .RN(n17132), .QN(n1411) );
  DFFR_X1 E9c3z4_reg ( .D(n13758), .CK(hclk), .RN(n17135), .QN(n1447) );
  DFFR_X1 Zqb3z4_reg ( .D(n14956), .CK(hclk), .RN(n17138), .QN(n1310) );
  DFFR_X1 D4g3z4_reg ( .D(n5707), .CK(hclk), .RN(n17133), .QN(n244) );
  DFFR_X1 Thm2z4_reg ( .D(n5824), .CK(hclk), .RN(n17135), .Q(vis_primask_o), 
        .QN(n1045) );
  DFFR_X1 Jje3z4_reg ( .D(n13846), .CK(hclk), .RN(n17132), .Q(n4755), .QN(
        n4338) );
  DFFR_X1 Wuq2z4_reg ( .D(n4897), .CK(hclk), .RN(n17132), .Q(n4751), .QN(n3775) );
  DFFR_X1 Uaj2z4_reg ( .D(n5689), .CK(hclk), .RN(n17131), .Q(vis_ipsr_o[2]), 
        .QN(n176) );
  DFFR_X1 Cam2z4_reg ( .D(n5687), .CK(hclk), .RN(n17130), .Q(vis_ipsr_o[3]), 
        .QN(n170) );
  DFFR_X1 Tdp2z4_reg ( .D(n5683), .CK(hclk), .RN(n17131), .Q(vis_ipsr_o[5]), 
        .QN(n159) );
  DFFR_X1 Trq2z4_reg ( .D(n5685), .CK(hclk), .RN(n17131), .Q(vis_ipsr_o[4]), 
        .QN(n165) );
  DFFR_X1 Idk2z4_reg ( .D(n5668), .CK(hclk), .RN(n17129), .Q(vis_apsr_o[0]), 
        .QN(n83) );
  DFFS_X1 Jcw2z4_reg ( .D(n4881), .CK(hclk), .SN(n17190), .QN(n4847) );
  DFFS_X1 Ydw2z4_reg ( .D(n4906), .CK(hclk), .SN(n17159), .Q(n367), .QN(n4777)
         );
  DFFS_X1 Xuw2z4_reg ( .D(n4917), .CK(hclk), .SN(n17194), .Q(n345), .QN(n4788)
         );
  DFFS_X1 Urw2z4_reg ( .D(n4915), .CK(hclk), .SN(n17192), .Q(n349), .QN(n4786)
         );
  DFFS_X1 Sow2z4_reg ( .D(n4913), .CK(hclk), .SN(n17159), .Q(n353), .QN(n4784)
         );
  DFFS_X1 Qzw2z4_reg ( .D(n4920), .CK(hclk), .SN(n17193), .Q(n339), .QN(n4791)
         );
  DFFS_X1 Qlw2z4_reg ( .D(n4911), .CK(hclk), .SN(n17159), .Q(n357), .QN(n4782)
         );
  DFFS_X1 Oiw2z4_reg ( .D(n4909), .CK(hclk), .SN(n17159), .Q(n361), .QN(n4780)
         );
  DFFS_X1 Mww2z4_reg ( .D(n4918), .CK(hclk), .SN(n17187), .Q(n343), .QN(n4789)
         );
  DFFS_X1 Mfw2z4_reg ( .D(n4907), .CK(hclk), .SN(n17159), .Q(n365), .QN(n4778)
         );
  DFFS_X1 Itw2z4_reg ( .D(n4916), .CK(hclk), .SN(n17188), .Q(n347), .QN(n4787)
         );
  DFFS_X1 Gqw2z4_reg ( .D(n4914), .CK(hclk), .SN(n17190), .Q(n351), .QN(n4785)
         );
  DFFS_X1 F1x2z4_reg ( .D(n4921), .CK(hclk), .SN(n17189), .Q(n372), .QN(n4792)
         );
  DFFS_X1 Enw2z4_reg ( .D(n4912), .CK(hclk), .SN(n17159), .Q(n355), .QN(n4783)
         );
  DFFS_X1 Ckw2z4_reg ( .D(n4910), .CK(hclk), .SN(n17159), .Q(n359), .QN(n4781)
         );
  DFFS_X1 Byw2z4_reg ( .D(n4919), .CK(hclk), .SN(n17191), .Q(n369), .QN(n4790)
         );
  DFFS_X1 Ahw2z4_reg ( .D(n4908), .CK(hclk), .SN(n17159), .Q(n363), .QN(n4779)
         );
  DFFS_X1 M1j2z4_reg ( .D(U691_Z_0), .CK(hclk), .SN(n17152), .Q(n3436), .QN(
        n4968) );
  DFFS_X1 B2i3z4_reg ( .D(n4885), .CK(hclk), .SN(n17156), .QN(n5639) );
  DFFS_X1 Ieh3z4_reg ( .D(n4890), .CK(hclk), .SN(n17153), .QN(n5625) );
  DFFS_X1 Xyn2z4_reg ( .D(n4888), .CK(hclk), .SN(n17187), .Q(n3250), .QN(n5067) );
  DFFS_X1 I1h3z4_reg ( .D(n4891), .CK(hclk), .SN(n17152), .QN(n5618) );
  DFFS_X1 Mka3z4_reg ( .D(n4871), .CK(hclk), .SN(n17164), .Q(n3012), .QN(n5514) );
  DFFS_X1 Gdo2z4_reg ( .D(n4892), .CK(hclk), .SN(n17152), .Q(n3381), .QN(n5074) );
  DFFS_X1 Gha3z4_reg ( .D(n4869), .CK(hclk), .SN(n17164), .Q(n3227), .QN(n5512) );
  DFFS_X1 Qfa3z4_reg ( .D(n4868), .CK(hclk), .SN(n17164), .Q(n3311), .QN(n5511) );
  DFFS_X1 Taa3z4_reg ( .D(n4867), .CK(hclk), .SN(n17164), .Q(n3056), .QN(n5509) );
  DFFS_X1 L8m2z4_reg ( .D(n4887), .CK(hclk), .SN(n17194), .Q(n3126), .QN(n5033) );
  DFFS_X1 Aea3z4_reg ( .D(n4861), .CK(hclk), .SN(n17172), .QN(n5510) );
  DFFS_X1 Wia3z4_reg ( .D(n4870), .CK(hclk), .SN(n17164), .Q(n3104), .QN(n5513) );
  DFFS_X1 Nfb3z4_reg ( .D(n4857), .CK(hclk), .SN(n17140), .QN(n5520) );
  DFFS_X1 J7b3z4_reg ( .D(n4859), .CK(hclk), .SN(n17166), .Q(n2946), .QN(n5517) );
  DFFS_X1 Cma3z4_reg ( .D(n4855), .CK(hclk), .SN(n17155), .Q(n2881), .QN(n5515) );
  DFFS_X1 Wzy2z4_reg ( .D(U105_Z_0), .CK(hclk), .SN(n17151), .Q(n3492), .QN(
        n5252) );
  DFFS_X1 Rni2z4_reg ( .D(U144_Z_0), .CK(hclk), .SN(n17141), .Q(n3495), .QN(
        n4959) );
  DFFS_X1 Kxe3z4_reg ( .D(n4889), .CK(hclk), .SN(n17188), .Q(n3326), .QN(n5579) );
  DFFS_X1 Bge3z4_reg ( .D(n4872), .CK(hclk), .SN(n17164), .Q(n3111), .QN(n5571) );
  DFFS_X1 C9a3z4_reg ( .D(n4866), .CK(hclk), .SN(n17164), .Q(n3268), .QN(n5508) );
  DFFS_X1 W3f3z4_reg ( .D(n4884), .CK(hclk), .SN(n17157), .QN(n5581) );
  DFFS_X1 T5g3z4_reg ( .D(n4873), .CK(hclk), .SN(n17164), .Q(n2986), .QN(n5600) );
  DFFS_X1 Hxx2z4_reg ( .D(n4879), .CK(hclk), .SN(n17143), .Q(n1008), .QN(n4845) );
  DFFS_X1 D4a3z4_reg ( .D(n4856), .CK(hclk), .SN(n17143), .QN(n5505) );
  DFFS_X1 U5a3z4_reg ( .D(n4858), .CK(hclk), .SN(n17165), .Q(n2917), .QN(n5506) );
  DFFS_X1 L7a3z4_reg ( .D(n4865), .CK(hclk), .SN(n17165), .QN(n5507) );
  DFFS_X1 Tyx2z4_reg ( .D(n5798), .CK(hclk), .SN(n17143), .Q(n1009) );
  DFFS_X1 Wai2z4_reg ( .D(n5800), .CK(hclk), .SN(n17165), .Q(n1759), .QN(n4947) );
  DFFS_X1 Yaz2z4_reg ( .D(U98_Z_0), .CK(hclk), .SN(n17141), .Q(n3493), .QN(
        n5259) );
  DFFS_X1 Svk2z4_reg ( .D(U122_Z_0), .CK(hclk), .SN(n17151), .Q(n3489), .QN(
        n5004) );
  DFFS_X1 T1d3z4_reg ( .D(U97_Z_0), .CK(hclk), .SN(n17141), .Q(n3496), .QN(
        n5544) );
  DFFS_X1 H3d3z4_reg ( .D(U754_Z_0), .CK(hclk), .SN(n17142), .Q(n1353), .QN(
        n5545) );
  DFFS_X1 W7z2z4_reg ( .D(n8706), .CK(hclk), .SN(n17141), .Q(n2827), .QN(n5257) );
  DFFS_X1 K9z2z4_reg ( .D(n8698), .CK(hclk), .SN(n17159), .Q(n2819), .QN(n5258) );
  DFFS_X1 I6z2z4_reg ( .D(n5779), .CK(hclk), .SN(n17141), .Q(n2865), .QN(n5256) );
  DFFS_X1 Qzq2z4_reg ( .D(U811_Z_0), .CK(hclk), .SN(n17154), .Q(n2172), .QN(
        n5120) );
  DFFS_X1 I2t2z4_reg ( .D(n5771), .CK(hclk), .SN(n17140), .Q(n486), .QN(n5162)
         );
  DFFS_X1 C3z2z4_reg ( .D(n5770), .CK(hclk), .SN(n17141), .Q(n1723), .QN(n5254) );
  DFFS_X1 K1z2z4_reg ( .D(n5772), .CK(hclk), .SN(n17140), .Q(n2731), .QN(n5253) );
  DFFS_X1 Auk2z4_reg ( .D(n5773), .CK(hclk), .SN(n17141), .Q(n2774), .QN(n5003) );
  DFFS_X1 Fzl2z4_reg ( .D(U795_Z_0), .CK(hclk), .SN(n17154), .Q(n2231), .QN(
        n5027) );
  DFFS_X1 Uup2z4_reg ( .D(U755_Z_0), .CK(hclk), .SN(n17153), .Q(n795), .QN(
        n5100) );
  DFFS_X1 Iwp2z4_reg ( .D(n5738), .CK(hclk), .SN(n17165), .Q(n2188), .QN(n5101) );
  DFFS_X1 Jw93z4_reg ( .D(n5786), .CK(hclk), .SN(n17163), .Q(n2620), .QN(n5500) );
  DFFS_X1 U4z2z4_reg ( .D(n5776), .CK(hclk), .SN(n17141), .Q(n2635), .QN(n5255) );
  DFFS_X1 Xx93z4_reg ( .D(n5784), .CK(hclk), .SN(n17163), .Q(n2593), .QN(n5501) );
  DFFS_X1 Ovc3z4_reg ( .D(n4944), .CK(hclk), .SN(n17164), .Q(n2570), .QN(n4853) );
  DFFS_X1 Qdj2z4_reg ( .D(n14928), .CK(hclk), .SN(n17155), .Q(n503), .QN(n4974) );
  DFFS_X1 Dvy2z4_reg ( .D(n5742), .CK(hclk), .SN(n17139), .Q(n16687), .QN(
        n16818) );
  DFFS_X1 Rxl2z4_reg ( .D(n5751), .CK(hclk), .SN(n17140), .Q(n461), .QN(n5026)
         );
  DFFS_X1 Viy2z4_reg ( .D(n5750), .CK(hclk), .SN(n17141), .Q(n454), .QN(n5241)
         );
  DFFS_X1 Efp2z4_reg ( .D(n4943), .CK(hclk), .SN(n17141), .Q(n2539), .QN(n4852) );
  DFFS_X1 U593z4_reg ( .D(n4927), .CK(hclk), .SN(n17165), .Q(n1152) );
  DFFS_X1 I793z4_reg ( .D(n4923), .CK(hclk), .SN(n17140), .Q(n2221), .QN(n4828) );
  DFFS_X1 Szr2z4_reg ( .D(n4940), .CK(hclk), .SN(n17157), .Q(n1161), .QN(n4851) );
  DFFS_X1 Rkd3z4_reg ( .D(n17212), .CK(hclk), .SN(n17144), .Q(n3142), .QN(
        n4771) );
  DFFS_X1 G1s2z4_reg ( .D(n5783), .CK(hclk), .SN(n17186), .Q(n869), .QN(n5140)
         );
  DFFS_X1 Dkr2z4_reg ( .D(n4937), .CK(hclk), .SN(n17161), .Q(n3028), .QN(n4830) );
  DFFS_X1 Wce3z4_reg ( .D(n4938), .CK(hclk), .SN(n17153), .Q(n3049), .QN(n4831) );
  DFFS_X1 G9w2z4_reg ( .D(n5828), .CK(hclk), .SN(n17156), .Q(n651), .QN(n5230)
         );
  DFFS_X1 Slr2z4_reg ( .D(n4936), .CK(hclk), .SN(n17153), .Q(n2970), .QN(n4832) );
  DFFS_X1 J7q2z4_reg ( .D(n4935), .CK(hclk), .SN(n17155), .Q(n2961), .QN(n4850) );
  DFFS_X1 Y8q2z4_reg ( .D(n4941), .CK(hclk), .SN(n17156), .Q(n1163), .QN(n4827) );
  DFFS_X1 H4p2z4_reg ( .D(n4933), .CK(hclk), .SN(n17192), .Q(n2817), .QN(n4769) );
  DFFS_X1 Ym93z4_reg ( .D(n4934), .CK(hclk), .SN(n17152), .Q(n2841), .QN(n4770) );
  DFFS_X1 F0y2z4_reg ( .D(n5764), .CK(hclk), .SN(n17155), .Q(n403), .QN(n5240)
         );
  DFFS_X1 Kyi2z4_reg ( .D(n5769), .CK(hclk), .SN(n17154), .Q(n413), .QN(n4966)
         );
  DFFS_X1 Gtp2z4_reg ( .D(n5766), .CK(hclk), .SN(n17153), .Q(n415), .QN(n5099)
         );
  DFFS_X1 Dwl2z4_reg ( .D(n5768), .CK(hclk), .SN(n17195), .QN(n5025) );
  DFFS_X1 W5p2z4_reg ( .D(n4932), .CK(hclk), .SN(n17190), .Q(n2795), .QN(n4768) );
  DFFS_X1 L7p2z4_reg ( .D(n4931), .CK(hclk), .SN(n17193), .Q(n2772), .QN(n4767) );
  DFFS_X1 Llq2z4_reg ( .D(n4929), .CK(hclk), .SN(n17153), .Q(n2714), .QN(n4765) );
  DFFS_X1 Tzg3z4_reg ( .D(n4930), .CK(hclk), .SN(n17152), .Q(n2746), .QN(n4766) );
  DFFS_X1 G6d3z4_reg ( .D(U317_Z_0), .CK(hclk), .SN(n17163), .QN(n5546) );
  DFFS_X1 Zfh3z4_reg ( .D(n4928), .CK(hclk), .SN(n17165), .Q(n2713), .QN(n4764) );
  DFFS_X1 B6j2z4_reg ( .D(n4942), .CK(hclk), .SN(n17152), .Q(n2515), .QN(n4772) );
  DFFS_X1 Q7j2z4_reg ( .D(n5737), .CK(hclk), .SN(n17152), .Q(n2481), .QN(n4971) );
  DFFS_X1 S8k2z4_reg ( .D(n4925), .CK(hclk), .SN(n17154), .Q(n2441), .QN(n4762) );
  DFFS_X1 Lgi3z4_reg ( .D(n4926), .CK(hclk), .SN(n17187), .Q(n2460), .QN(n4763) );
  DFFS_X1 Ohh3z4_reg ( .D(n5787), .CK(hclk), .SN(n17154), .Q(n2279), .QN(n5626) );
  DFFS_X1 Hak2z4_reg ( .D(n4924), .CK(hclk), .SN(n17153), .Q(n2280), .QN(n4761) );
  DFFS_X1 Cqo2z4_reg ( .D(n5788), .CK(hclk), .SN(n17154), .Q(n881), .QN(n4773)
         );
  DFFS_X1 Rhi2z4_reg ( .D(n5785), .CK(hclk), .SN(n17151), .Q(n874), .QN(n4955)
         );
  DFFS_X1 Rbi3z4_reg ( .D(n4945), .CK(hclk), .SN(n17151), .QN(n4846) );
  DFFS_X1 V1l2z4_reg ( .D(n5782), .CK(hclk), .SN(n17154), .Q(n867), .QN(n4774)
         );
  DFFR_X1 Nen2z4_reg ( .D(U692_Z_0), .CK(hclk), .RN(n17195), .Q(vis_control_o), 
        .QN(n5055) );
  DFFR_X1 Zei2z4_reg ( .D(U809_Z_0), .CK(hclk), .RN(n17128), .Q(vis_apsr_o[1]), 
        .QN(n4953) );
  DFFR_X1 S4w2z4_reg ( .D(n4880), .CK(hclk), .RN(hreset_n), .Q(n596), .QN(
        n5228) );
  DFFR_X1 J6i2z4_reg ( .D(n5711), .CK(hclk), .RN(n17129), .Q(n251), .QN(n4905)
         );
  DFFR_X1 Ffs2z4_reg ( .D(n5791), .CK(hclk), .RN(n17130), .Q(n1110), .QN(n5149) );
  DFFR_X1 Lz93z4_reg ( .D(n5790), .CK(hclk), .RN(n17132), .Q(n4073), .QN(n5502) );
  DFFS_X1 Zjq2z4_reg ( .D(n5665), .CK(hclk), .SN(n17191), .Q(vis_pc_o[18]), 
        .QN(n5114) );
  DFFS_X1 Plx2z4_reg ( .D(n5663), .CK(hclk), .SN(n17188), .Q(vis_pc_o[16]), 
        .QN(n5236) );
  DFFS_X1 Foe3z4_reg ( .D(n5660), .CK(hclk), .SN(n17153), .Q(vis_pc_o[20]), 
        .QN(n5573) );
  DFFS_X1 Dkx2z4_reg ( .D(n5664), .CK(hclk), .SN(n17152), .Q(vis_pc_o[15]), 
        .QN(n5235) );
  DFFS_X1 Bnx2z4_reg ( .D(n5662), .CK(hclk), .SN(n17186), .Q(vis_pc_o[17]), 
        .QN(n5237) );
  DFFS_X1 B9g3z4_reg ( .D(n5659), .CK(hclk), .SN(n17152), .Q(vis_pc_o[19]), 
        .QN(n5601) );
  DFFS_X1 Rix2z4_reg ( .D(n5677), .CK(hclk), .SN(n17155), .Q(vis_pc_o[13]), 
        .QN(n4813) );
  DFFS_X1 Gmd3z4_reg ( .D(n5675), .CK(hclk), .SN(n17143), .Q(vis_pc_o[10]), 
        .QN(n4815) );
  DFFS_X1 Fhx2z4_reg ( .D(n5678), .CK(hclk), .SN(n17143), .Q(vis_pc_o[11]), 
        .QN(n4812) );
  DFFS_X1 V4d3z4_reg ( .D(n5676), .CK(hclk), .SN(n17144), .Q(vis_pc_o[8]), 
        .QN(n4814) );
  DFFS_X1 Ycx2z4_reg ( .D(n5656), .CK(hclk), .SN(n17160), .Q(vis_pc_o[6]), 
        .QN(n4825) );
  DFFS_X1 Nbx2z4_reg ( .D(n5681), .CK(hclk), .SN(n17160), .Q(vis_pc_o[5]) );
  DFFS_X1 J4x2z4_reg ( .D(n5688), .CK(hclk), .SN(n17160), .Q(vis_pc_o[1]), 
        .QN(n5233) );
  DFFS_X1 G7x2z4_reg ( .D(n5686), .CK(hclk), .SN(n17160), .Q(vis_pc_o[2]) );
  DFFS_X1 Cax2z4_reg ( .D(n5682), .CK(hclk), .SN(n17160), .Q(vis_pc_o[4]) );
  DFFS_X1 R8x2z4_reg ( .D(n5684), .CK(hclk), .SN(n17160), .Q(vis_pc_o[3]) );
  DFFS_X1 Zjg3z4_reg ( .D(U474_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r10_o[20]), 
        .QN(n5608) );
  DFFS_X1 Z523z4_reg ( .D(U407_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r11_o[16]), 
        .QN(n5325) );
  DFFS_X1 Y6o2z4_reg ( .D(U409_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r5_o[16]), 
        .QN(n5070) );
  DFFS_X1 Wu53z4_reg ( .D(U438_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r8_o[18]), 
        .QN(n5410) );
  DFFS_X1 Wrg3z4_reg ( .D(U479_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r7_o[20]), 
        .QN(n5613) );
  DFFS_X1 Vgg3z4_reg ( .D(U472_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r8_o[20]), 
        .QN(n5606) );
  DFFS_X1 V223z4_reg ( .D(U441_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r11_o[18]), 
        .QN(n5323) );
  DFFS_X1 Tvn2z4_reg ( .D(U448_Z_0), .CK(hclk), .SN(n17170), .Q(vis_msp_o[16]), 
        .QN(n5065) );
  DFFS_X1 Sog3z4_reg ( .D(U477_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r5_o[20]), 
        .QN(n5611) );
  DFFS_X1 Skv2z4_reg ( .D(U408_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r4_o[16]), 
        .QN(n5218) );
  DFFS_X1 Sg83z4_reg ( .D(U402_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r2_o[16]), 
        .QN(n5470) );
  DFFS_X1 Ro43z4_reg ( .D(U405_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r9_o[16]), 
        .QN(n5383) );
  DFFS_X1 Rdg3z4_reg ( .D(U470_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r2_o[20]), 
        .QN(n5604) );
  DFFS_X1 Rbo2z4_reg ( .D(U415_Z_0), .CK(hclk), .SN(n17171), .Q(vis_psp_o[14]), 
        .QN(n5073) );
  DFFS_X1 Pwg3z4_reg ( .D(U482_Z_0), .CK(hclk), .SN(n17168), .Q(vis_msp_o[18]), 
        .QN(n5616) );
  DFFS_X1 Psn2z4_reg ( .D(U443_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r5_o[18]), 
        .QN(n5063) );
  DFFS_X1 Olg3z4_reg ( .D(U475_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r11_o[20]), 
        .QN(n5609) );
  DFFS_X1 Ohv2z4_reg ( .D(U442_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r4_o[18]), 
        .QN(n5216) );
  DFFS_X1 Od83z4_reg ( .D(U436_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r2_o[18]), 
        .QN(n5468) );
  DFFS_X1 O403z4_reg ( .D(U412_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r12_o[16]), 
        .QN(n5278) );
  DFFS_X1 Nl43z4_reg ( .D(U439_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r9_o[18]), 
        .QN(n5381) );
  DFFS_X1 Nag3z4_reg ( .D(U468_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r0_o[20]), 
        .QN(n5602) );
  DFFS_X1 N8o2z4_reg ( .D(U411_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r7_o[16]), 
        .QN(n5071) );
  DFFS_X1 Ltg3z4_reg ( .D(U480_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r12_o[20]), 
        .QN(n5614) );
  DFFS_X1 Kig3z4_reg ( .D(U473_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r9_o[20]), 
        .QN(n5607) );
  DFFS_X1 K103z4_reg ( .D(U446_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r12_o[18]), 
        .QN(n5276) );
  DFFS_X1 Jl93z4_reg ( .D(U400_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r0_o[16]), 
        .QN(n5494) );
  DFFS_X1 Jbu2z4_reg ( .D(U410_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r6_o[16]), 
        .QN(n5189) );
  DFFS_X1 J773z4_reg ( .D(U403_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r3_o[16]), 
        .QN(n5441) );
  DFFS_X1 J5o2z4_reg ( .D(U401_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r1_o[16]), 
        .QN(n5069) );
  DFFS_X1 Ixn2z4_reg ( .D(U449_Z_0), .CK(hclk), .SN(n17170), .Q(vis_psp_o[16]), 
        .QN(n5066) );
  DFFS_X1 If33z4_reg ( .D(U406_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r10_o[16]), 
        .QN(n5354) );
  DFFS_X1 I113z4_reg ( .D(U413_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r14_o[16]), 
        .QN(n5299) );
  DFFS_X1 Hqg3z4_reg ( .D(U478_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r6_o[20]), 
        .QN(n5612) );
  DFFS_X1 Gfg3z4_reg ( .D(U471_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r3_o[20]), 
        .QN(n5605) );
  DFFS_X1 Fi93z4_reg ( .D(U434_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r0_o[18]), 
        .QN(n5492) );
  DFFS_X1 F473z4_reg ( .D(U437_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r3_o[18]), 
        .QN(n5439) );
  DFFS_X1 F8u2z4_reg ( .D(U444_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r6_o[18]), 
        .QN(n5187) );
  DFFS_X1 Eyg3z4_reg ( .D(U483_Z_0), .CK(hclk), .SN(n17168), .Q(vis_psp_o[18]), 
        .QN(n5617) );
  DFFS_X1 Ey03z4_reg ( .D(U447_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r14_o[18]), 
        .QN(n5297) );
  DFFS_X1 Eun2z4_reg ( .D(U445_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r7_o[18]), 
        .QN(n5064) );
  DFFS_X1 Ec33z4_reg ( .D(U440_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r10_o[18]), 
        .QN(n5352) );
  DFFS_X1 Dng3z4_reg ( .D(U476_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r4_o[20]), 
        .QN(n5610) );
  DFFS_X1 Ccg3z4_reg ( .D(U469_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r1_o[20]), 
        .QN(n5603) );
  DFFS_X1 Cao2z4_reg ( .D(U414_Z_0), .CK(hclk), .SN(n17171), .Q(vis_msp_o[14]), 
        .QN(n5072) );
  DFFS_X1 Ay53z4_reg ( .D(U404_Z_0), .CK(hclk), .SN(n17172), .Q(vis_r8_o[16]), 
        .QN(n5412) );
  DFFS_X1 Avg3z4_reg ( .D(U481_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r14_o[20]), 
        .QN(n5615) );
  DFFS_X1 Arn2z4_reg ( .D(U435_Z_0), .CK(hclk), .SN(n17171), .Q(vis_r1_o[18]), 
        .QN(n5062) );
  DFFS_X1 Zxo2z4_reg ( .D(U427_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[17]), 
        .QN(n5084) );
  DFFS_X1 Zfv2z4_reg ( .D(U460_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r4_o[19]), 
        .QN(n5215) );
  DFFS_X1 Zb83z4_reg ( .D(U454_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r2_o[19]), 
        .QN(n5467) );
  DFFS_X1 Z203z4_reg ( .D(U430_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[17]), 
        .QN(n5277) );
  DFFS_X1 Yj43z4_reg ( .D(U457_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r9_o[19]), 
        .QN(n5380) );
  DFFS_X1 Xyh3z4_reg ( .D(U466_Z_0), .CK(hclk), .SN(n17169), .Q(vis_msp_o[17]), 
        .QN(n5637) );
  DFFS_X1 Uj93z4_reg ( .D(U418_Z_0), .CK(hclk), .SN(n17191), .Q(vis_r0_o[17]), 
        .QN(n5493) );
  DFFS_X1 U573z4_reg ( .D(U421_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[17]), 
        .QN(n5440) );
  DFFS_X1 U9u2z4_reg ( .D(U428_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[17]), 
        .QN(n5188) );
  DFFS_X1 Tz03z4_reg ( .D(U431_Z_0), .CK(hclk), .SN(n17143), .Q(vis_r14_o[17]), 
        .QN(n5298) );
  DFFS_X1 Tvh3z4_reg ( .D(U464_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r12_o[19]), 
        .QN(n5635) );
  DFFS_X1 Td33z4_reg ( .D(U424_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[17]), 
        .QN(n5353) );
  DFFS_X1 S2p2z4_reg ( .D(U433_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[15]), 
        .QN(n5087) );
  DFFS_X1 Qg93z4_reg ( .D(U452_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r0_o[19]), 
        .QN(n5491) );
  DFFS_X1 Q273z4_reg ( .D(U455_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r3_o[19]), 
        .QN(n5438) );
  DFFS_X1 Q6u2z4_reg ( .D(U462_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r6_o[19]), 
        .QN(n5186) );
  DFFS_X1 Pap2z4_reg ( .D(U461_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r5_o[19]), 
        .QN(n5089) );
  DFFS_X1 Pa33z4_reg ( .D(U458_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r10_o[19]), 
        .QN(n5351) );
  DFFS_X1 Ozo2z4_reg ( .D(U429_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[17]), 
        .QN(n5085) );
  DFFS_X1 M0i3z4_reg ( .D(U467_Z_0), .CK(hclk), .SN(n17169), .Q(vis_psp_o[17]), 
        .QN(n5638) );
  DFFS_X1 Lw53z4_reg ( .D(U422_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[17]), 
        .QN(n5411) );
  DFFS_X1 Kwo2z4_reg ( .D(U419_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[17]), 
        .QN(n5083) );
  DFFS_X1 K423z4_reg ( .D(U425_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[17]), 
        .QN(n5324) );
  DFFS_X1 Ixh3z4_reg ( .D(U465_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r14_o[19]), 
        .QN(n5636) );
  DFFS_X1 Ht53z4_reg ( .D(U456_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r8_o[19]), 
        .QN(n5409) );
  DFFS_X1 G123z4_reg ( .D(U459_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r11_o[19]), 
        .QN(n5322) );
  DFFS_X1 Ecp2z4_reg ( .D(U463_Z_0), .CK(hclk), .SN(n17169), .Q(vis_r7_o[19]), 
        .QN(n5090) );
  DFFS_X1 Djv2z4_reg ( .D(U426_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[17]), 
        .QN(n5217) );
  DFFS_X1 Df83z4_reg ( .D(U420_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[17]), 
        .QN(n5469) );
  DFFS_X1 D1p2z4_reg ( .D(U432_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[15]), 
        .QN(n5086) );
  DFFS_X1 Cn43z4_reg ( .D(U423_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[17]), 
        .QN(n5382) );
  DFFS_X1 A9p2z4_reg ( .D(U453_Z_0), .CK(hclk), .SN(n17170), .Q(vis_r1_o[19]), 
        .QN(n5088) );
  DFFS_X1 Nox2z4_reg ( .D(n5661), .CK(hclk), .SN(n17165), .Q(vis_pc_o[21]), 
        .QN(n5238) );
  DFFS_X1 Tch3z4_reg ( .D(U501_Z_0), .CK(hclk), .SN(n17167), .Q(vis_psp_o[19]), 
        .QN(n5624) );
  DFFS_X1 Sr53z4_reg ( .D(U490_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r8_o[21]), 
        .QN(n5408) );
  DFFS_X1 Rz13z4_reg ( .D(U493_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r11_o[21]), 
        .QN(n5321) );
  DFFS_X1 Poq2z4_reg ( .D(U495_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r5_o[21]), 
        .QN(n5116) );
  DFFS_X1 P9h3z4_reg ( .D(U499_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r14_o[21]), 
        .QN(n5622) );
  DFFS_X1 Kev2z4_reg ( .D(U494_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r4_o[21]), 
        .QN(n5214) );
  DFFS_X1 Ka83z4_reg ( .D(U488_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r2_o[21]), 
        .QN(n5466) );
  DFFS_X1 Ji43z4_reg ( .D(U491_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r9_o[21]), 
        .QN(n5379) );
  DFFS_X1 Eqq2z4_reg ( .D(U497_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r7_o[21]), 
        .QN(n5117) );
  DFFS_X1 Ebh3z4_reg ( .D(U500_Z_0), .CK(hclk), .SN(n17167), .Q(vis_msp_o[19]), 
        .QN(n5623) );
  DFFS_X1 Bf93z4_reg ( .D(U486_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r0_o[21]), 
        .QN(n5490) );
  DFFS_X1 B173z4_reg ( .D(U489_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r3_o[21]), 
        .QN(n5437) );
  DFFS_X1 B5u2z4_reg ( .D(U496_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r6_o[21]), 
        .QN(n5185) );
  DFFS_X1 Anq2z4_reg ( .D(U487_Z_0), .CK(hclk), .SN(n17168), .Q(vis_r1_o[21]), 
        .QN(n5115) );
  DFFS_X1 A933z4_reg ( .D(U492_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r10_o[21]), 
        .QN(n5350) );
  DFFS_X1 A8h3z4_reg ( .D(U498_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r12_o[21]), 
        .QN(n5621) );
  DFFS_X1 Kaf3z4_reg ( .D(n5657), .CK(hclk), .SN(n17190), .Q(vis_pc_o[22]), 
        .QN(n4824) );
  DFFS_X1 Tme3z4_reg ( .D(n5674), .CK(hclk), .SN(n17153), .Q(vis_pc_o[12]), 
        .QN(n4816) );
  DFFS_X1 Ufx2z4_reg ( .D(n5679), .CK(hclk), .SN(n17143), .Q(vis_pc_o[9]), 
        .QN(n4811) );
  DFFS_X1 Jwf3z4_reg ( .D(n5658), .CK(hclk), .SN(n17143), .Q(vis_pc_o[14]) );
  DFFS_X1 Jex2z4_reg ( .D(n5680), .CK(hclk), .SN(n17160), .Q(vis_pc_o[7]) );
  DFFS_X1 W5s2z4_reg ( .D(U295_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r7_o[9]), 
        .QN(n5143) );
  DFFS_X1 Uku2z4_reg ( .D(U294_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r6_o[9]), 
        .QN(n5195) );
  DFFS_X1 Ug73z4_reg ( .D(U287_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[9]), 
        .QN(n5447) );
  DFFS_X1 U2s2z4_reg ( .D(U285_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[9]), 
        .QN(n5141) );
  DFFS_X1 Tse3z4_reg ( .D(U298_Z_0), .CK(hclk), .SN(n17175), .Q(vis_msp_o[7]), 
        .QN(n5576) );
  DFFS_X1 To33z4_reg ( .D(U290_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[9]), 
        .QN(n5360) );
  DFFS_X1 Rpe3z4_reg ( .D(U296_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[9]), 
        .QN(n5574) );
  DFFS_X1 L763z4_reg ( .D(U288_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[9]), 
        .QN(n5418) );
  DFFS_X1 Kf23z4_reg ( .D(U291_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r11_o[9]), 
        .QN(n5331) );
  DFFS_X1 I4s2z4_reg ( .D(U293_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[9]), 
        .QN(n5142) );
  DFFS_X1 Hue3z4_reg ( .D(U299_Z_0), .CK(hclk), .SN(n17180), .Q(vis_psp_o[7]), 
        .QN(n5577) );
  DFFS_X1 Fre3z4_reg ( .D(U297_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r14_o[9]), 
        .QN(n5575) );
  DFFS_X1 Duv2z4_reg ( .D(U292_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[9]), 
        .QN(n5224) );
  DFFS_X1 Dq83z4_reg ( .D(U286_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[9]), 
        .QN(n5476) );
  DFFS_X1 Cy43z4_reg ( .D(U289_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[9]), 
        .QN(n5389) );
  DFFS_X1 Cxc3z4_reg ( .D(U284_Z_0), .CK(hclk), .SN(n17152), .Q(vis_r0_o[9]), 
        .QN(n5541) );
  DFFS_X1 Zgr2z4_reg ( .D(U366_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[10]), 
        .QN(n5130) );
  DFFS_X1 Vdr2z4_reg ( .D(U361_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[12]), 
        .QN(n5128) );
  DFFS_X1 T263z4_reg ( .D(U356_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[12]), 
        .QN(n5415) );
  DFFS_X1 Sa23z4_reg ( .D(U359_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[12]), 
        .QN(n5328) );
  DFFS_X1 S703z4_reg ( .D(U364_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[12]), 
        .QN(n5280) );
  DFFS_X1 Rr93z4_reg ( .D(U352_Z_0), .CK(hclk), .SN(n17153), .Q(vis_r0_o[12]), 
        .QN(n5497) );
  DFFS_X1 Oir2z4_reg ( .D(U367_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[10]), 
        .QN(n5131) );
  DFFS_X1 M413z4_reg ( .D(U365_Z_0), .CK(hclk), .SN(n17143), .Q(vis_r14_o[12]), 
        .QN(n5301) );
  DFFS_X1 Lpv2z4_reg ( .D(U360_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[12]), 
        .QN(n5221) );
  DFFS_X1 Ll83z4_reg ( .D(U354_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[12]), 
        .QN(n5473) );
  DFFS_X1 Kt43z4_reg ( .D(U357_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[12]), 
        .QN(n5386) );
  DFFS_X1 Kfr2z4_reg ( .D(U363_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r7_o[12]), 
        .QN(n5129) );
  DFFS_X1 Gcr2z4_reg ( .D(U353_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[12]), 
        .QN(n5127) );
  DFFS_X1 Cgu2z4_reg ( .D(U362_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[12]), 
        .QN(n5192) );
  DFFS_X1 Cc73z4_reg ( .D(U355_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[12]), 
        .QN(n5444) );
  DFFS_X1 Bk33z4_reg ( .D(U358_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[12]), 
        .QN(n5357) );
  DFFS_X1 Y1n2z4_reg ( .D(U511_Z_0), .CK(hclk), .SN(n17164), .Q(vis_r5_o[22]), 
        .QN(n5049) );
  DFFS_X1 Vzz2z4_reg ( .D(U514_Z_0), .CK(hclk), .SN(n17165), .Q(vis_r12_o[22]), 
        .QN(n5275) );
  DFFS_X1 Vcv2z4_reg ( .D(U510_Z_0), .CK(hclk), .SN(n17164), .Q(vis_r4_o[22]), 
        .QN(n5213) );
  DFFS_X1 V883z4_reg ( .D(U504_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r2_o[22]), 
        .QN(n5465) );
  DFFS_X1 Ug43z4_reg ( .D(U507_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r9_o[22]), 
        .QN(n5378) );
  DFFS_X1 R6n2z4_reg ( .D(U517_Z_0), .CK(hclk), .SN(n17165), .Q(vis_psp_o[20]), 
        .QN(n5052) );
  DFFS_X1 Pw03z4_reg ( .D(U515_Z_0), .CK(hclk), .SN(n17165), .Q(vis_r14_o[22]), 
        .QN(n5296) );
  DFFS_X1 N3n2z4_reg ( .D(U513_Z_0), .CK(hclk), .SN(n17165), .Q(vis_r7_o[22]), 
        .QN(n5050) );
  DFFS_X1 Mz63z4_reg ( .D(U505_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r3_o[22]), 
        .QN(n5436) );
  DFFS_X1 Md93z4_reg ( .D(U502_Z_0), .CK(hclk), .SN(n17141), .Q(vis_r0_o[22]), 
        .QN(n5489) );
  DFFS_X1 M3u2z4_reg ( .D(U512_Z_0), .CK(hclk), .SN(n17164), .Q(vis_r6_o[22]), 
        .QN(n5184) );
  DFFS_X1 L733z4_reg ( .D(U508_Z_0), .CK(hclk), .SN(n17164), .Q(vis_r10_o[22]), 
        .QN(n5349) );
  DFFS_X1 J0n2z4_reg ( .D(U503_Z_0), .CK(hclk), .SN(n17140), .Q(vis_r1_o[22]), 
        .QN(n5048) );
  DFFS_X1 Dq53z4_reg ( .D(U506_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r8_o[22]), 
        .QN(n5407) );
  DFFS_X1 Cy13z4_reg ( .D(U509_Z_0), .CK(hclk), .SN(n17164), .Q(vis_r11_o[22]), 
        .QN(n5320) );
  DFFS_X1 C5n2z4_reg ( .D(U516_Z_0), .CK(hclk), .SN(n17165), .Q(vis_msp_o[20]), 
        .QN(n5051) );
  DFFS_X1 Z853z4_reg ( .D(U738_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r8_o[0]), 
        .QN(n5396) );
  DFFS_X1 Yg13z4_reg ( .D(U723_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r11_o[0]), 
        .QN(n5309) );
  DFFS_X1 Unm2z4_reg ( .D(U803_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r0_o[0]), 
        .QN(n5040) );
  DFFS_X1 Skm2z4_reg ( .D(U708_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r7_o[0]), 
        .QN(n5038) );
  DFFS_X1 Rvu2z4_reg ( .D(U693_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r4_o[0]), 
        .QN(n5202) );
  DFFS_X1 Rr73z4_reg ( .D(U748_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r2_o[0]), 
        .QN(n5454) );
  DFFS_X1 Qz33z4_reg ( .D(U733_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r9_o[0]), 
        .QN(n5367) );
  DFFS_X1 Knz2z4_reg ( .D(U713_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r12_o[0]), 
        .QN(n5267) );
  DFFS_X1 Imt2z4_reg ( .D(U703_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r6_o[0]), 
        .QN(n5173) );
  DFFS_X1 Ii63z4_reg ( .D(U743_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r3_o[0]), 
        .QN(n5425) );
  DFFS_X1 Hq23z4_reg ( .D(U728_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r10_o[0]), 
        .QN(n5338) );
  DFFS_X1 Gmm2z4_reg ( .D(U797_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r1_o[0]), 
        .QN(n5039) );
  DFFS_X1 Ek03z4_reg ( .D(U718_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r14_o[0]), 
        .QN(n5288) );
  DFFS_X1 Ejm2z4_reg ( .D(U698_Z_0), .CK(hclk), .SN(n17166), .Q(vis_r5_o[0]), 
        .QN(n5037) );
  DFFS_X1 Yfn2z4_reg ( .D(U301_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[2]), 
        .QN(n5056) );
  DFFS_X1 X563z4_reg ( .D(U304_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[2]), 
        .QN(n5417) );
  DFFS_X1 Wd23z4_reg ( .D(U307_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r11_o[2]), 
        .QN(n5330) );
  DFFS_X1 Wa03z4_reg ( .D(U312_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[2]), 
        .QN(n5282) );
  DFFS_X1 Vu93z4_reg ( .D(U300_Z_0), .CK(hclk), .SN(n17154), .Q(vis_r0_o[2]), 
        .QN(n5499) );
  DFFS_X1 Q713z4_reg ( .D(U313_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r14_o[2]), 
        .QN(n5303) );
  DFFS_X1 Psv2z4_reg ( .D(U308_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[2]), 
        .QN(n5223) );
  DFFS_X1 Po83z4_reg ( .D(U302_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[2]), 
        .QN(n5475) );
  DFFS_X1 Ow43z4_reg ( .D(U305_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[2]), 
        .QN(n5388) );
  DFFS_X1 Okn2z4_reg ( .D(U314_Z_0), .CK(hclk), .SN(n17175), .Q(vis_msp_o[0]), 
        .QN(n5059) );
  DFFS_X1 Mhn2z4_reg ( .D(U309_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[2]), 
        .QN(n5057) );
  DFFS_X1 Gju2z4_reg ( .D(U310_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r6_o[2]), 
        .QN(n5194) );
  DFFS_X1 Gf73z4_reg ( .D(U303_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[2]), 
        .QN(n5446) );
  DFFS_X1 Fn33z4_reg ( .D(U306_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[2]), 
        .QN(n5359) );
  DFFS_X1 Cmn2z4_reg ( .D(U315_Z_0), .CK(hclk), .SN(n17151), .Q(vis_psp_o[0]), 
        .QN(n5060) );
  DFFS_X1 Ajn2z4_reg ( .D(U311_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r7_o[2]), 
        .QN(n5058) );
  DFFS_X1 Z7i2z4_reg ( .D(n14825), .CK(hclk), .SN(n17140), .Q(vis_tbit_o), 
        .QN(n4922) );
  DFFS_X1 Yx63z4_reg ( .D(U522_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[3]), 
        .QN(n5435) );
  DFFS_X1 Yb93z4_reg ( .D(U519_Z_0), .CK(hclk), .SN(n17151), .Q(vis_r0_o[3]), 
        .QN(n5488) );
  DFFS_X1 Y1u2z4_reg ( .D(U529_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[3]), 
        .QN(n5183) );
  DFFS_X1 X533z4_reg ( .D(U525_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[3]), 
        .QN(n5348) );
  DFFS_X1 X6m2z4_reg ( .D(U534_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[1]), 
        .QN(n5032) );
  DFFS_X1 V3m2z4_reg ( .D(U530_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[3]), 
        .QN(n5030) );
  DFFS_X1 T0m2z4_reg ( .D(U520_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[3]), 
        .QN(n5028) );
  DFFS_X1 Po53z4_reg ( .D(U523_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[3]), 
        .QN(n5406) );
  DFFS_X1 Ow13z4_reg ( .D(U526_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[3]), 
        .QN(n5319) );
  DFFS_X1 J5m2z4_reg ( .D(U533_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[1]), 
        .QN(n5031) );
  DFFS_X1 Hyz2z4_reg ( .D(U531_Z_0), .CK(hclk), .SN(n17160), .Q(vis_r12_o[3]), 
        .QN(n5274) );
  DFFS_X1 Hbv2z4_reg ( .D(U527_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[3]), 
        .QN(n5212) );
  DFFS_X1 H783z4_reg ( .D(U521_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[3]), 
        .QN(n5464) );
  DFFS_X1 H2m2z4_reg ( .D(U528_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[3]), 
        .QN(n5029) );
  DFFS_X1 Gf43z4_reg ( .D(U524_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[3]), 
        .QN(n5377) );
  DFFS_X1 Bv03z4_reg ( .D(U532_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[3]), 
        .QN(n5295) );
  DFFS_X1 Zr03z4_reg ( .D(U564_Z_0), .CK(hclk), .SN(n17143), .Q(vis_r14_o[5]), 
        .QN(n5293) );
  DFFS_X1 Wyt2z4_reg ( .D(U561_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[5]), 
        .QN(n5181) );
  DFFS_X1 Wu63z4_reg ( .D(U554_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[5]), 
        .QN(n5433) );
  DFFS_X1 Wmp2z4_reg ( .D(U566_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[3]), 
        .QN(n5095) );
  DFFS_X1 W893z4_reg ( .D(U551_Z_0), .CK(hclk), .SN(n17194), .Q(vis_r0_o[5]), 
        .QN(n5486) );
  DFFS_X1 V233z4_reg ( .D(U557_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[5]), 
        .QN(n5346) );
  DFFS_X1 Ujp2z4_reg ( .D(U562_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[5]), 
        .QN(n5093) );
  DFFS_X1 Sgp2z4_reg ( .D(U552_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[5]), 
        .QN(n5091) );
  DFFS_X1 Nl53z4_reg ( .D(U555_Z_0), .CK(hclk), .SN(n17156), .Q(vis_r8_o[5]), 
        .QN(n5404) );
  DFFS_X1 Mt13z4_reg ( .D(U558_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[5]), 
        .QN(n5317) );
  DFFS_X1 Ilp2z4_reg ( .D(U565_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[3]), 
        .QN(n5094) );
  DFFS_X1 Gip2z4_reg ( .D(U560_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[5]), 
        .QN(n5092) );
  DFFS_X1 Fvz2z4_reg ( .D(U563_Z_0), .CK(hclk), .SN(n17160), .Q(vis_r12_o[5]), 
        .QN(n5272) );
  DFFS_X1 F483z4_reg ( .D(U553_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[5]), 
        .QN(n5462) );
  DFFS_X1 F8v2z4_reg ( .D(U559_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[5]), 
        .QN(n5210) );
  DFFS_X1 Ec43z4_reg ( .D(U556_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[5]), 
        .QN(n5375) );
  DFFS_X1 U5r2z4_reg ( .D(U549_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[2]), 
        .QN(n5124) );
  DFFS_X1 Twz2z4_reg ( .D(U547_Z_0), .CK(hclk), .SN(n17160), .Q(vis_r12_o[4]), 
        .QN(n5273) );
  DFFS_X1 T583z4_reg ( .D(U537_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[4]), 
        .QN(n5463) );
  DFFS_X1 T9v2z4_reg ( .D(U543_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[4]), 
        .QN(n5211) );
  DFFS_X1 Sd43z4_reg ( .D(U540_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[4]), 
        .QN(n5376) );
  DFFS_X1 S2r2z4_reg ( .D(U544_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[4]), 
        .QN(n5122) );
  DFFS_X1 Nt03z4_reg ( .D(U548_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[4]), 
        .QN(n5294) );
  DFFS_X1 Kw63z4_reg ( .D(U538_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[4]), 
        .QN(n5434) );
  DFFS_X1 Ka93z4_reg ( .D(U535_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r0_o[4]), 
        .QN(n5487) );
  DFFS_X1 K0u2z4_reg ( .D(U545_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[4]), 
        .QN(n5182) );
  DFFS_X1 J433z4_reg ( .D(U541_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[4]), 
        .QN(n5347) );
  DFFS_X1 I7r2z4_reg ( .D(U550_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[2]), 
        .QN(n5125) );
  DFFS_X1 G4r2z4_reg ( .D(U546_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[4]), 
        .QN(n5123) );
  DFFS_X1 E1r2z4_reg ( .D(U536_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[4]), 
        .QN(n5121) );
  DFFS_X1 Bn53z4_reg ( .D(U539_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r8_o[4]), 
        .QN(n5405) );
  DFFS_X1 Av13z4_reg ( .D(U542_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[4]), 
        .QN(n5318) );
  DFFS_X1 Zu43z4_reg ( .D(U323_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[10]), 
        .QN(n5387) );
  DFFS_X1 Z8s2z4_reg ( .D(U327_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[10]), 
        .QN(n5145) );
  DFFS_X1 Rhu2z4_reg ( .D(U328_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[10]), 
        .QN(n5193) );
  DFFS_X1 Rds2z4_reg ( .D(U333_Z_0), .CK(hclk), .SN(n17151), .Q(vis_psp_o[8]), 
        .QN(n5148) );
  DFFS_X1 Rd73z4_reg ( .D(U321_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[10]), 
        .QN(n5445) );
  DFFS_X1 Ql33z4_reg ( .D(U324_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[10]), 
        .QN(n5358) );
  DFFS_X1 Oas2z4_reg ( .D(U329_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r7_o[10]), 
        .QN(n5146) );
  DFFS_X1 K7s2z4_reg ( .D(U319_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[10]), 
        .QN(n5144) );
  DFFS_X1 I463z4_reg ( .D(U322_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[10]), 
        .QN(n5416) );
  DFFS_X1 Hc23z4_reg ( .D(U325_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[10]), 
        .QN(n5329) );
  DFFS_X1 H903z4_reg ( .D(U330_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[10]), 
        .QN(n5281) );
  DFFS_X1 Gt93z4_reg ( .D(U318_Z_0), .CK(hclk), .SN(n17153), .Q(vis_r0_o[10]), 
        .QN(n5498) );
  DFFS_X1 Dcs2z4_reg ( .D(U332_Z_0), .CK(hclk), .SN(n17175), .Q(vis_msp_o[8]), 
        .QN(n5147) );
  DFFS_X1 B613z4_reg ( .D(U331_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r14_o[10]), 
        .QN(n5302) );
  DFFS_X1 Arv2z4_reg ( .D(U326_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[10]), 
        .QN(n5222) );
  DFFS_X1 An83z4_reg ( .D(U320_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[10]), 
        .QN(n5474) );
  DFFS_X1 Xyk2z4_reg ( .D(n5672), .CK(hclk), .SN(n17152), .Q(vis_pc_o[23]) );
  DFFS_X1 Wnu2z4_reg ( .D(U260_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r6_o[15]), 
        .QN(n5197) );
  DFFS_X1 Wj73z4_reg ( .D(U253_Z_0), .CK(hclk), .SN(n17195), .Q(vis_r3_o[15]), 
        .QN(n5449) );
  DFFS_X1 Vr33z4_reg ( .D(U256_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r10_o[15]), 
        .QN(n5362) );
  DFFS_X1 Rdq2z4_reg ( .D(U261_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r7_o[15]), 
        .QN(n5110) );
  DFFS_X1 Psh3z4_reg ( .D(U264_Z_0), .CK(hclk), .SN(n17175), .Q(vis_msp_o[13]), 
        .QN(n5633) );
  DFFS_X1 Naq2z4_reg ( .D(U251_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[15]), 
        .QN(n5108) );
  DFFS_X1 Na63z4_reg ( .D(U254_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r8_o[15]), 
        .QN(n5420) );
  DFFS_X1 Mi23z4_reg ( .D(U257_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r11_o[15]), 
        .QN(n5333) );
  DFFS_X1 Lph3z4_reg ( .D(U262_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[15]), 
        .QN(n5631) );
  DFFS_X1 Fxv2z4_reg ( .D(U258_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[15]), 
        .QN(n5226) );
  DFFS_X1 Ft83z4_reg ( .D(U252_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[15]), 
        .QN(n5478) );
  DFFS_X1 Euh3z4_reg ( .D(U265_Z_0), .CK(hclk), .SN(n17173), .Q(vis_psp_o[13]), 
        .QN(n5634) );
  DFFS_X1 E153z4_reg ( .D(U255_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[15]), 
        .QN(n5391) );
  DFFS_X1 E0d3z4_reg ( .D(U250_Z_0), .CK(hclk), .SN(n17186), .Q(vis_r0_o[15]), 
        .QN(n5543) );
  DFFS_X1 Ccq2z4_reg ( .D(U259_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r5_o[15]), 
        .QN(n5109) );
  DFFS_X1 Arh3z4_reg ( .D(U263_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r14_o[15]), 
        .QN(n5632) );
  DFFS_X1 Z863z4_reg ( .D(U272_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[8]), 
        .QN(n5419) );
  DFFS_X1 Yg23z4_reg ( .D(U275_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r11_o[8]), 
        .QN(n5332) );
  DFFS_X1 Rvv2z4_reg ( .D(U276_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[8]), 
        .QN(n5225) );
  DFFS_X1 Rr83z4_reg ( .D(U270_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[8]), 
        .QN(n5477) );
  DFFS_X1 Qz43z4_reg ( .D(U273_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[8]), 
        .QN(n5390) );
  DFFS_X1 Qyc3z4_reg ( .D(U268_Z_0), .CK(hclk), .SN(n17152), .Q(vis_r0_o[8]), 
        .QN(n5542) );
  DFFS_X1 Qwr2z4_reg ( .D(U282_Z_0), .CK(hclk), .SN(n17175), .Q(vis_msp_o[6]), 
        .QN(n5138) );
  DFFS_X1 Otr2z4_reg ( .D(U277_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r5_o[8]), 
        .QN(n5136) );
  DFFS_X1 Kc03z4_reg ( .D(U280_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[8]), 
        .QN(n5283) );
  DFFS_X1 Imu2z4_reg ( .D(U278_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r6_o[8]), 
        .QN(n5196) );
  DFFS_X1 Ii73z4_reg ( .D(U271_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[8]), 
        .QN(n5448) );
  DFFS_X1 Hq33z4_reg ( .D(U274_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[8]), 
        .QN(n5361) );
  DFFS_X1 Eyr2z4_reg ( .D(U283_Z_0), .CK(hclk), .SN(n17173), .Q(vis_psp_o[6]), 
        .QN(n5139) );
  DFFS_X1 E913z4_reg ( .D(U281_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r14_o[8]), 
        .QN(n5304) );
  DFFS_X1 Cvr2z4_reg ( .D(U279_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r7_o[8]), 
        .QN(n5137) );
  DFFS_X1 Asr2z4_reg ( .D(U269_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[8]), 
        .QN(n5135) );
  DFFS_X1 Fcj2z4_reg ( .D(n5690), .CK(hclk), .SN(n17158), .Q(vis_pc_o[0]), 
        .QN(n4973) );
  DFFS_X1 Zj53z4_reg ( .D(U571_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r8_o[6]), 
        .QN(n5403) );
  DFFS_X1 Ytm2z4_reg ( .D(U581_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[4]), 
        .QN(n5044) );
  DFFS_X1 Yr13z4_reg ( .D(U574_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[6]), 
        .QN(n5316) );
  DFFS_X1 Wqm2z4_reg ( .D(U576_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[6]), 
        .QN(n5042) );
  DFFS_X1 Rtz2z4_reg ( .D(U579_Z_0), .CK(hclk), .SN(n17160), .Q(vis_r12_o[6]), 
        .QN(n5271) );
  DFFS_X1 R283z4_reg ( .D(U569_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[6]), 
        .QN(n5461) );
  DFFS_X1 R6v2z4_reg ( .D(U575_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[6]), 
        .QN(n5209) );
  DFFS_X1 Qa43z4_reg ( .D(U572_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[6]), 
        .QN(n5374) );
  DFFS_X1 Mvm2z4_reg ( .D(U582_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[4]), 
        .QN(n5045) );
  DFFS_X1 Lq03z4_reg ( .D(U580_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[6]), 
        .QN(n5292) );
  DFFS_X1 Ksm2z4_reg ( .D(U578_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[6]), 
        .QN(n5043) );
  DFFS_X1 Ixt2z4_reg ( .D(U577_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[6]), 
        .QN(n5180) );
  DFFS_X1 It63z4_reg ( .D(U570_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[6]), 
        .QN(n5432) );
  DFFS_X1 Ipm2z4_reg ( .D(U568_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[6]), 
        .QN(n5041) );
  DFFS_X1 H133z4_reg ( .D(U573_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[6]), 
        .QN(n5345) );
  DFFS_X1 G493z4_reg ( .D(U567_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r0_o[6]), 
        .QN(n5485) );
  DFFS_X1 X553z4_reg ( .D(U740_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r8_o[7]), 
        .QN(n5394) );
  DFFS_X1 Wd13z4_reg ( .D(U725_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r11_o[7]), 
        .QN(n5307) );
  DFFS_X1 Spl2z4_reg ( .D(U799_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[7]), 
        .QN(n5021) );
  DFFS_X1 Qml2z4_reg ( .D(U700_Z_0), .CK(hclk), .SN(n17175), .Q(vis_r5_o[7]), 
        .QN(n5019) );
  DFFS_X1 Psu2z4_reg ( .D(U695_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r4_o[7]), 
        .QN(n5200) );
  DFFS_X1 Po73z4_reg ( .D(U750_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[7]), 
        .QN(n5452) );
  DFFS_X1 Ow33z4_reg ( .D(U735_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[7]), 
        .QN(n5365) );
  DFFS_X1 Mcz2z4_reg ( .D(U687_Z_0), .CK(hclk), .SN(n17149), .Q(vis_psp_o[5]), 
        .QN(n5260) );
  DFFS_X1 Ikz2z4_reg ( .D(U715_Z_0), .CK(hclk), .SN(n17186), .Q(vis_r12_o[7]), 
        .QN(n5265) );
  DFFS_X1 Grl2z4_reg ( .D(U804_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r0_o[7]), 
        .QN(n5022) );
  DFFS_X1 Gjt2z4_reg ( .D(U705_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r6_o[7]), 
        .QN(n5171) );
  DFFS_X1 Gf63z4_reg ( .D(U745_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r3_o[7]), 
        .QN(n5423) );
  DFFS_X1 Fn23z4_reg ( .D(U730_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r10_o[7]), 
        .QN(n5336) );
  DFFS_X1 Eol2z4_reg ( .D(U710_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r7_o[7]), 
        .QN(n5020) );
  DFFS_X1 Cll2z4_reg ( .D(U684_Z_0), .CK(hclk), .SN(n17158), .Q(vis_msp_o[5]), 
        .QN(n5018) );
  DFFS_X1 Ch03z4_reg ( .D(U720_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[7]), 
        .QN(n5286) );
  DFFS_X1 Ycu2z4_reg ( .D(U394_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[14]), 
        .QN(n5190) );
  DFFS_X1 Y873z4_reg ( .D(U387_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[14]), 
        .QN(n5442) );
  DFFS_X1 Xg33z4_reg ( .D(U390_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[14]), 
        .QN(n5355) );
  DFFS_X1 X213z4_reg ( .D(U397_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[14]), 
        .QN(n5300) );
  DFFS_X1 U5q2z4_reg ( .D(U399_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[12]), 
        .QN(n5107) );
  DFFS_X1 Q2q2z4_reg ( .D(U395_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[14]), 
        .QN(n5105) );
  DFFS_X1 Pz53z4_reg ( .D(U388_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[14]), 
        .QN(n5413) );
  DFFS_X1 O723z4_reg ( .D(U391_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[14]), 
        .QN(n5326) );
  DFFS_X1 No93z4_reg ( .D(U384_Z_0), .CK(hclk), .SN(n17153), .Q(vis_r0_o[14]), 
        .QN(n5495) );
  DFFS_X1 Mzp2z4_reg ( .D(U385_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[14]), 
        .QN(n5103) );
  DFFS_X1 Hmv2z4_reg ( .D(U392_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[14]), 
        .QN(n5219) );
  DFFS_X1 Hi83z4_reg ( .D(U386_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[14]), 
        .QN(n5471) );
  DFFS_X1 Gq43z4_reg ( .D(U389_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[14]), 
        .QN(n5384) );
  DFFS_X1 F4q2z4_reg ( .D(U398_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[12]), 
        .QN(n5106) );
  DFFS_X1 D603z4_reg ( .D(U396_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[14]), 
        .QN(n5279) );
  DFFS_X1 B1q2z4_reg ( .D(U393_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[14]), 
        .QN(n5104) );
  DFFS_X1 Wlz2z4_reg ( .D(U714_Z_0), .CK(hclk), .SN(n17194), .Q(vis_r12_o[1]), 
        .QN(n5266) );
  DFFS_X1 Ukt2z4_reg ( .D(U704_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r6_o[1]), 
        .QN(n5172) );
  DFFS_X1 Ug63z4_reg ( .D(U744_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r3_o[1]), 
        .QN(n5424) );
  DFFS_X1 Txj2z4_reg ( .D(U810_Z_0), .CK(hclk), .SN(n17192), .Q(vis_r0_o[1]), 
        .QN(n4987) );
  DFFS_X1 To23z4_reg ( .D(U729_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r10_o[1]), 
        .QN(n5337) );
  DFFS_X1 Ruj2z4_reg ( .D(U709_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[1]), 
        .QN(n4985) );
  DFFS_X1 Qi03z4_reg ( .D(U719_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[1]), 
        .QN(n5287) );
  DFFS_X1 L753z4_reg ( .D(U739_Z_0), .CK(hclk), .SN(n17156), .Q(vis_r8_o[1]), 
        .QN(n5395) );
  DFFS_X1 Kf13z4_reg ( .D(U724_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r11_o[1]), 
        .QN(n5308) );
  DFFS_X1 Fwj2z4_reg ( .D(U798_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[1]), 
        .QN(n4986) );
  DFFS_X1 Duu2z4_reg ( .D(U694_Z_0), .CK(hclk), .SN(n17193), .Q(vis_r4_o[1]), 
        .QN(n5201) );
  DFFS_X1 Dtj2z4_reg ( .D(U699_Z_0), .CK(hclk), .SN(n17175), .Q(vis_r5_o[1]), 
        .QN(n4984) );
  DFFS_X1 Dq73z4_reg ( .D(U749_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[1]), 
        .QN(n5453) );
  DFFS_X1 Cy33z4_reg ( .D(U734_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[1]), 
        .QN(n5366) );
  DFFS_X1 Xmf3z4_reg ( .D(U240_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[23]), 
        .QN(n5590) );
  DFFS_X1 Wbf3z4_reg ( .D(U232_Z_0), .CK(hclk), .SN(n17155), .Q(vis_r0_o[23]), 
        .QN(n5583) );
  DFFS_X1 Uuf3z4_reg ( .D(U247_Z_0), .CK(hclk), .SN(n17173), .Q(vis_psp_o[21]), 
        .QN(n5595) );
  DFFS_X1 Tjf3z4_reg ( .D(U238_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r10_o[23]), 
        .QN(n5588) );
  DFFS_X1 Qrf3z4_reg ( .D(U244_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[23]), 
        .QN(n5593) );
  DFFS_X1 Mof3z4_reg ( .D(U241_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r5_o[23]), 
        .QN(n5591) );
  DFFS_X1 Eif3z4_reg ( .D(U237_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[23]), 
        .QN(n5587) );
  DFFS_X1 Orj2z4_reg ( .D(U233_Z_0), .CK(hclk), .SN(n17155), .Q(vis_r1_o[23]), 
        .QN(n4983) );
  DFFS_X1 Ftf3z4_reg ( .D(U245_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r14_o[23]), 
        .QN(n5594) );
  DFFS_X1 Pgf3z4_reg ( .D(U236_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r8_o[23]), 
        .QN(n5586) );
  DFFS_X1 M4j2z4_reg ( .D(U246_Z_0), .CK(hclk), .SN(n17175), .Q(vis_msp_o[21]), 
        .QN(n4970) );
  DFFS_X1 Ilf3z4_reg ( .D(U239_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r11_o[23]), 
        .QN(n5589) );
  DFFS_X1 Aff3z4_reg ( .D(U235_Z_0), .CK(hclk), .SN(n17192), .Q(vis_r3_o[23]), 
        .QN(n5585) );
  DFFS_X1 Bqf3z4_reg ( .D(U242_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r6_o[23]), 
        .QN(n5592) );
  DFFS_X1 Ldf3z4_reg ( .D(U234_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[23]), 
        .QN(n5584) );
  DFFS_X1 Fpi2z4_reg ( .D(U243_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r7_o[23]), 
        .QN(n4960) );
  DFFS_X1 Zpx2z4_reg ( .D(n5671), .CK(hclk), .SN(n17156), .Q(vis_pc_o[24]), 
        .QN(n4819) );
  DFFS_X1 X1e3z4_reg ( .D(U343_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[11]), 
        .QN(n5563) );
  DFFS_X1 Wqd3z4_reg ( .D(U336_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[11]), 
        .QN(n5556) );
  DFFS_X1 U9e3z4_reg ( .D(U348_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[9]), 
        .QN(n5568) );
  DFFS_X1 Tyd3z4_reg ( .D(U341_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[11]), 
        .QN(n5561) );
  DFFS_X1 Snd3z4_reg ( .D(U334_Z_0), .CK(hclk), .SN(n17153), .Q(vis_r0_o[11]), 
        .QN(n5554) );
  DFFS_X1 Q6e3z4_reg ( .D(U346_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[11]), 
        .QN(n5566) );
  DFFS_X1 Pvd3z4_reg ( .D(U339_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[11]), 
        .QN(n5559) );
  DFFS_X1 M3e3z4_reg ( .D(U344_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[11]), 
        .QN(n5564) );
  DFFS_X1 Lsd3z4_reg ( .D(U337_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[11]), 
        .QN(n5557) );
  DFFS_X1 Ibe3z4_reg ( .D(U349_Z_0), .CK(hclk), .SN(n17151), .Q(vis_psp_o[9]), 
        .QN(n5569) );
  DFFS_X1 I0e3z4_reg ( .D(U342_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[11]), 
        .QN(n5562) );
  DFFS_X1 Hpd3z4_reg ( .D(U335_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[11]), 
        .QN(n5555) );
  DFFS_X1 F8e3z4_reg ( .D(U347_Z_0), .CK(hclk), .SN(n17143), .Q(vis_r14_o[11]), 
        .QN(n5567) );
  DFFS_X1 Exd3z4_reg ( .D(U340_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[11]), 
        .QN(n5560) );
  DFFS_X1 B5e3z4_reg ( .D(U345_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r7_o[11]), 
        .QN(n5565) );
  DFFS_X1 Aud3z4_reg ( .D(U338_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[11]), 
        .QN(n5558) );
  DFFS_X1 Z0g3z4_reg ( .D(U382_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[11]), 
        .QN(n5598) );
  DFFS_X1 Wor2z4_reg ( .D(U377_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[13]), 
        .QN(n5133) );
  DFFS_X1 Wnv2z4_reg ( .D(U376_Z_0), .CK(hclk), .SN(n17163), .Q(vis_r4_o[13]), 
        .QN(n5220) );
  DFFS_X1 Wj83z4_reg ( .D(U370_Z_0), .CK(hclk), .SN(n17149), .Q(vis_r2_o[13]), 
        .QN(n5472) );
  DFFS_X1 Vxf3z4_reg ( .D(U380_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r12_o[13]), 
        .QN(n5596) );
  DFFS_X1 Vr43z4_reg ( .D(U373_Z_0), .CK(hclk), .SN(n17178), .Q(vis_r9_o[13]), 
        .QN(n5385) );
  DFFS_X1 O2g3z4_reg ( .D(U383_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[11]), 
        .QN(n5599) );
  DFFS_X1 Neu2z4_reg ( .D(U378_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[13]), 
        .QN(n5191) );
  DFFS_X1 Na73z4_reg ( .D(U371_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[13]), 
        .QN(n5443) );
  DFFS_X1 Mi33z4_reg ( .D(U374_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[13]), 
        .QN(n5356) );
  DFFS_X1 Lqr2z4_reg ( .D(U379_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[13]), 
        .QN(n5134) );
  DFFS_X1 Kzf3z4_reg ( .D(U381_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[13]), 
        .QN(n5597) );
  DFFS_X1 Hnr2z4_reg ( .D(U369_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r1_o[13]), 
        .QN(n5132) );
  DFFS_X1 E163z4_reg ( .D(U372_Z_0), .CK(hclk), .SN(n17157), .Q(vis_r8_o[13]), 
        .QN(n5414) );
  DFFS_X1 D923z4_reg ( .D(U375_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[13]), 
        .QN(n5327) );
  DFFS_X1 Cq93z4_reg ( .D(U368_Z_0), .CK(hclk), .SN(n17152), .Q(vis_r0_o[13]), 
        .QN(n5496) );
  DFFS_X1 Zpj2z4_reg ( .D(U584_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[24]), 
        .QN(n4982) );
  DFFS_X1 Vmj2z4_reg ( .D(U592_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[24]), 
        .QN(n4980) );
  DFFS_X1 Umi3z4_reg ( .D(U597_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[22]), 
        .QN(n5646) );
  DFFS_X1 Tvt2z4_reg ( .D(U593_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[24]), 
        .QN(n5179) );
  DFFS_X1 Tr63z4_reg ( .D(U586_Z_0), .CK(hclk), .SN(n17185), .Q(vis_r3_o[24]), 
        .QN(n5431) );
  DFFS_X1 Sz23z4_reg ( .D(U589_Z_0), .CK(hclk), .SN(n17147), .Q(vis_r10_o[24]), 
        .QN(n5344) );
  DFFS_X1 R293z4_reg ( .D(U583_Z_0), .CK(hclk), .SN(n17189), .Q(vis_r0_o[24]), 
        .QN(n5484) );
  DFFS_X1 Qji3z4_reg ( .D(U595_Z_0), .CK(hclk), .SN(n17160), .Q(vis_r12_o[24]), 
        .QN(n5644) );
  DFFS_X1 Ki53z4_reg ( .D(U587_Z_0), .CK(hclk), .SN(n17156), .Q(vis_r8_o[24]), 
        .QN(n5402) );
  DFFS_X1 Jq13z4_reg ( .D(U590_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[24]), 
        .QN(n5315) );
  DFFS_X1 Joi3z4_reg ( .D(U598_Z_0), .CK(hclk), .SN(n17139), .Q(vis_psp_o[22]), 
        .QN(n5647) );
  DFFS_X1 Fli3z4_reg ( .D(U596_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[24]), 
        .QN(n5645) );
  DFFS_X1 F9j2z4_reg ( .D(U594_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[24]), 
        .QN(n4972) );
  DFFS_X1 C183z4_reg ( .D(U585_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[24]), 
        .QN(n5460) );
  DFFS_X1 C5v2z4_reg ( .D(U591_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[24]), 
        .QN(n5208) );
  DFFS_X1 B943z4_reg ( .D(U588_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[24]), 
        .QN(n5373) );
  DFFS_X1 Lrx2z4_reg ( .D(n5670), .CK(hclk), .SN(n17187), .Q(vis_pc_o[25]), 
        .QN(n4820) );
  DFFS_X1 Xhl2z4_reg ( .D(U614_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[23]), 
        .QN(n5016) );
  DFFS_X1 Wo03z4_reg ( .D(U612_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[25]), 
        .QN(n5291) );
  DFFS_X1 Vg53z4_reg ( .D(U603_Z_0), .CK(hclk), .SN(n17156), .Q(vis_r8_o[25]), 
        .QN(n5401) );
  DFFS_X1 Uo13z4_reg ( .D(U606_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[25]), 
        .QN(n5314) );
  DFFS_X1 Tel2z4_reg ( .D(U610_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[25]), 
        .QN(n5014) );
  DFFS_X1 Pbl2z4_reg ( .D(U600_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[25]), 
        .QN(n5012) );
  DFFS_X1 Nz73z4_reg ( .D(U601_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[25]), 
        .QN(n5459) );
  DFFS_X1 N3v2z4_reg ( .D(U607_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[25]), 
        .QN(n5207) );
  DFFS_X1 M743z4_reg ( .D(U604_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[25]), 
        .QN(n5372) );
  DFFS_X1 Igl2z4_reg ( .D(U613_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[23]), 
        .QN(n5015) );
  DFFS_X1 Eut2z4_reg ( .D(U609_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[25]), 
        .QN(n5178) );
  DFFS_X1 Eq63z4_reg ( .D(U602_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r3_o[25]), 
        .QN(n5430) );
  DFFS_X1 Edl2z4_reg ( .D(U608_Z_0), .CK(hclk), .SN(n17176), .Q(vis_r5_o[25]), 
        .QN(n5013) );
  DFFS_X1 Dy23z4_reg ( .D(U605_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r10_o[25]), 
        .QN(n5343) );
  DFFS_X1 Csz2z4_reg ( .D(U611_Z_0), .CK(hclk), .SN(n17160), .Q(vis_r12_o[25]), 
        .QN(n5270) );
  DFFS_X1 C193z4_reg ( .D(U599_Z_0), .CK(hclk), .SN(n17194), .Q(vis_r0_o[25]), 
        .QN(n5483) );
  DFFS_X1 Xsx2z4_reg ( .D(n5669), .CK(hclk), .SN(n17188), .Q(vis_pc_o[26]), 
        .QN(n4821) );
  DFFS_X1 Z3k2z4_reg ( .D(U628_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[26]), 
        .QN(n4991) );
  DFFS_X1 Yx73z4_reg ( .D(U619_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[26]), 
        .QN(n5458) );
  DFFS_X1 Y1v2z4_reg ( .D(U625_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[26]), 
        .QN(n5206) );
  DFFS_X1 X543z4_reg ( .D(U622_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[26]), 
        .QN(n5371) );
  DFFS_X1 V0k2z4_reg ( .D(U618_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[26]), 
        .QN(n4989) );
  DFFS_X1 Pst2z4_reg ( .D(U627_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[26]), 
        .QN(n5177) );
  DFFS_X1 Po63z4_reg ( .D(U620_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r3_o[26]), 
        .QN(n5429) );
  DFFS_X1 Ow23z4_reg ( .D(U623_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r10_o[26]), 
        .QN(n5342) );
  DFFS_X1 O5k2z4_reg ( .D(U631_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[24]), 
        .QN(n4992) );
  DFFS_X1 Nz83z4_reg ( .D(U617_Z_0), .CK(hclk), .SN(n17191), .Q(vis_r0_o[26]), 
        .QN(n5482) );
  DFFS_X1 Nqz2z4_reg ( .D(U629_Z_0), .CK(hclk), .SN(n17167), .Q(vis_r12_o[26]), 
        .QN(n5269) );
  DFFS_X1 K2k2z4_reg ( .D(U626_Z_0), .CK(hclk), .SN(n17175), .Q(vis_r5_o[26]), 
        .QN(n4990) );
  DFFS_X1 Hn03z4_reg ( .D(U630_Z_0), .CK(hclk), .SN(n17143), .Q(vis_r14_o[26]), 
        .QN(n5290) );
  DFFS_X1 Gf53z4_reg ( .D(U621_Z_0), .CK(hclk), .SN(n17156), .Q(vis_r8_o[26]), 
        .QN(n5400) );
  DFFS_X1 Fn13z4_reg ( .D(U624_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[26]), 
        .QN(n5313) );
  DFFS_X1 D7k2z4_reg ( .D(U632_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[24]), 
        .QN(n4993) );
  DFFS_X1 Jux2z4_reg ( .D(n5667), .CK(hclk), .SN(n17191), .Q(vis_pc_o[27]), 
        .QN(n4822) );
  DFFS_X1 Aez2z4_reg ( .D(U686_Z_0), .CK(hclk), .SN(n17151), .Q(vis_psp_o[26]), 
        .QN(n5261) );
  DFFS_X1 Zu33z4_reg ( .D(U736_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[28]), 
        .QN(n5364) );
  DFFS_X1 Zkk2z4_reg ( .D(U806_Z_0), .CK(hclk), .SN(n17155), .Q(vis_r0_o[28]), 
        .QN(n4998) );
  DFFS_X1 Tiz2z4_reg ( .D(U716_Z_0), .CK(hclk), .SN(n17193), .Q(vis_r12_o[28]), 
        .QN(n5264) );
  DFFS_X1 Ql23z4_reg ( .D(U731_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r10_o[28]), 
        .QN(n5335) );
  DFFS_X1 Ggk2z4_reg ( .D(U701_Z_0), .CK(hclk), .SN(n17175), .Q(vis_r5_o[28]), 
        .QN(n4995) );
  DFFS_X1 Aru2z4_reg ( .D(U696_Z_0), .CK(hclk), .SN(n17154), .Q(vis_r4_o[28]), 
        .QN(n5199) );
  DFFS_X1 Nf03z4_reg ( .D(U721_Z_0), .CK(hclk), .SN(n17141), .Q(vis_r14_o[28]), 
        .QN(n5285) );
  DFFS_X1 Kjk2z4_reg ( .D(U800_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[28]), 
        .QN(n4997) );
  DFFS_X1 Rek2z4_reg ( .D(U683_Z_0), .CK(hclk), .SN(n17160), .Q(vis_msp_o[26]), 
        .QN(n4994) );
  DFFS_X1 Rd63z4_reg ( .D(U746_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r3_o[28]), 
        .QN(n5422) );
  DFFS_X1 I453z4_reg ( .D(U741_Z_0), .CK(hclk), .SN(n17156), .Q(vis_r8_o[28]), 
        .QN(n5393) );
  DFFS_X1 Hc13z4_reg ( .D(U726_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r11_o[28]), 
        .QN(n5306) );
  DFFS_X1 Rht2z4_reg ( .D(U706_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r6_o[28]), 
        .QN(n5170) );
  DFFS_X1 An73z4_reg ( .D(U751_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[28]), 
        .QN(n5451) );
  DFFS_X1 Vhk2z4_reg ( .D(U711_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r7_o[28]), 
        .QN(n4996) );
  DFFS_X1 Zu23z4_reg ( .D(U639_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r10_o[27]), 
        .QN(n5341) );
  DFFS_X1 Yx83z4_reg ( .D(U633_Z_0), .CK(hclk), .SN(n17154), .Q(vis_r0_o[27]), 
        .QN(n5481) );
  DFFS_X1 Wnh3z4_reg ( .D(U648_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[25]), 
        .QN(n5630) );
  DFFS_X1 Vgq2z4_reg ( .D(U642_Z_0), .CK(hclk), .SN(n17175), .Q(vis_r5_o[27]), 
        .QN(n5112) );
  DFFS_X1 Skh3z4_reg ( .D(U646_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[27]), 
        .QN(n5628) );
  DFFS_X1 Rd53z4_reg ( .D(U637_Z_0), .CK(hclk), .SN(n17156), .Q(vis_r8_o[27]), 
        .QN(n5399) );
  DFFS_X1 Ql13z4_reg ( .D(U640_Z_0), .CK(hclk), .SN(n17183), .Q(vis_r11_o[27]), 
        .QN(n5312) );
  DFFS_X1 Kiq2z4_reg ( .D(U644_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[27]), 
        .QN(n5113) );
  DFFS_X1 Jw73z4_reg ( .D(U635_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[27]), 
        .QN(n5457) );
  DFFS_X1 J0v2z4_reg ( .D(U641_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[27]), 
        .QN(n5205) );
  DFFS_X1 I443z4_reg ( .D(U638_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[27]), 
        .QN(n5370) );
  DFFS_X1 Hmh3z4_reg ( .D(U647_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[25]), 
        .QN(n5629) );
  DFFS_X1 Gfq2z4_reg ( .D(U634_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[27]), 
        .QN(n5111) );
  DFFS_X1 Djh3z4_reg ( .D(U645_Z_0), .CK(hclk), .SN(n17187), .Q(vis_r12_o[27]), 
        .QN(n5627) );
  DFFS_X1 Art2z4_reg ( .D(U643_Z_0), .CK(hclk), .SN(n17145), .Q(vis_r6_o[27]), 
        .QN(n5176) );
  DFFS_X1 An63z4_reg ( .D(U636_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r3_o[27]), 
        .QN(n5428) );
  DFFS_X1 Vvx2z4_reg ( .D(n5666), .CK(hclk), .SN(n17153), .Q(vis_pc_o[28]), 
        .QN(n5239) );
  DFFS_X1 Omk2z4_reg ( .D(n5673), .CK(hclk), .SN(n17155), .Q(vis_pc_o[29]), 
        .QN(n4817) );
  DFFS_X1 J0l2z4_reg ( .D(n5655), .CK(hclk), .SN(n17152), .Q(vis_pc_o[30]), 
        .QN(n5006) );
  DFFS_X1 Y6i3z4_reg ( .D(U679_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[30]), 
        .QN(n5641) );
  DFFS_X1 Wnt2z4_reg ( .D(U676_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r6_o[30]), 
        .QN(n5174) );
  DFFS_X1 Wj63z4_reg ( .D(U669_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r3_o[30]), 
        .QN(n5426) );
  DFFS_X1 Vuo2z4_reg ( .D(U677_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[30]), 
        .QN(n5082) );
  DFFS_X1 Vr23z4_reg ( .D(U672_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r10_o[30]), 
        .QN(n5339) );
  DFFS_X1 Uu83z4_reg ( .D(U666_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r0_o[30]), 
        .QN(n5479) );
  DFFS_X1 Rro2z4_reg ( .D(U667_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[30]), 
        .QN(n5080) );
  DFFS_X1 Na53z4_reg ( .D(U670_Z_0), .CK(hclk), .SN(n17158), .Q(vis_r8_o[30]), 
        .QN(n5397) );
  DFFS_X1 N8i3z4_reg ( .D(U680_Z_0), .CK(hclk), .SN(n17173), .Q(vis_msp_o[28]), 
        .QN(n5642) );
  DFFS_X1 Mi13z4_reg ( .D(U673_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r11_o[30]), 
        .QN(n5310) );
  DFFS_X1 J5i3z4_reg ( .D(U678_Z_0), .CK(hclk), .SN(n17188), .Q(vis_r12_o[30]), 
        .QN(n5640) );
  DFFS_X1 Gto2z4_reg ( .D(U675_Z_0), .CK(hclk), .SN(n17175), .Q(vis_r5_o[30]), 
        .QN(n5081) );
  DFFS_X1 Fxu2z4_reg ( .D(U674_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[30]), 
        .QN(n5203) );
  DFFS_X1 Ft73z4_reg ( .D(U668_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[30]), 
        .QN(n5455) );
  DFFS_X1 E143z4_reg ( .D(U671_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[30]), 
        .QN(n5368) );
  DFFS_X1 Cai3z4_reg ( .D(U681_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[28]), 
        .QN(n5643) );
  DFFS_X1 Yoz2z4_reg ( .D(U661_Z_0), .CK(hclk), .SN(n17195), .Q(vis_r12_o[29]), 
        .QN(n5268) );
  DFFS_X1 Ymo2z4_reg ( .D(U663_Z_0), .CK(hclk), .SN(n17174), .Q(vis_msp_o[27]), 
        .QN(n5078) );
  DFFS_X1 Uyu2z4_reg ( .D(U657_Z_0), .CK(hclk), .SN(n17162), .Q(vis_r4_o[29]), 
        .QN(n5204) );
  DFFS_X1 Uu73z4_reg ( .D(U651_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[29]), 
        .QN(n5456) );
  DFFS_X1 Ujo2z4_reg ( .D(U658_Z_0), .CK(hclk), .SN(n17175), .Q(vis_r5_o[29]), 
        .QN(n5076) );
  DFFS_X1 T243z4_reg ( .D(U654_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[29]), 
        .QN(n5369) );
  DFFS_X1 Sl03z4_reg ( .D(U662_Z_0), .CK(hclk), .SN(n17142), .Q(vis_r14_o[29]), 
        .QN(n5289) );
  DFFS_X1 Noo2z4_reg ( .D(U664_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[27]), 
        .QN(n5079) );
  DFFS_X1 Lpt2z4_reg ( .D(U659_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r6_o[29]), 
        .QN(n5175) );
  DFFS_X1 Ll63z4_reg ( .D(U652_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r3_o[29]), 
        .QN(n5427) );
  DFFS_X1 Kt23z4_reg ( .D(U655_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r10_o[29]), 
        .QN(n5340) );
  DFFS_X1 Jw83z4_reg ( .D(U649_Z_0), .CK(hclk), .SN(n17151), .Q(vis_r0_o[29]), 
        .QN(n5480) );
  DFFS_X1 Jlo2z4_reg ( .D(U660_Z_0), .CK(hclk), .SN(n17181), .Q(vis_r7_o[29]), 
        .QN(n5077) );
  DFFS_X1 Fio2z4_reg ( .D(U650_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[29]), 
        .QN(n5075) );
  DFFS_X1 Cc53z4_reg ( .D(U653_Z_0), .CK(hclk), .SN(n17156), .Q(vis_r8_o[29]), 
        .QN(n5398) );
  DFFS_X1 Bk13z4_reg ( .D(U656_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r11_o[29]), 
        .QN(n5311) );
  DFFS_X1 Yd03z4_reg ( .D(U722_Z_0), .CK(hclk), .SN(n17143), .Q(vis_r14_o[31]), 
        .QN(n5284) );
  DFFS_X1 Xti2z4_reg ( .D(U805_Z_0), .CK(hclk), .SN(n17155), .Q(vis_r0_o[31]), 
        .QN(n4963) );
  DFFS_X1 X2j2z4_reg ( .D(U682_Z_0), .CK(hclk), .SN(n17173), .Q(vis_msp_o[29]), 
        .QN(n4969) );
  DFFS_X1 T253z4_reg ( .D(U742_Z_0), .CK(hclk), .SN(n17156), .Q(vis_r8_o[31]), 
        .QN(n5392) );
  DFFS_X1 Sa13z4_reg ( .D(U727_Z_0), .CK(hclk), .SN(n17182), .Q(vis_r11_o[31]), 
        .QN(n5305) );
  DFFS_X1 Pfz2z4_reg ( .D(U685_Z_0), .CK(hclk), .SN(n17150), .Q(vis_psp_o[29]), 
        .QN(n5262) );
  DFFS_X1 Lpu2z4_reg ( .D(U697_Z_0), .CK(hclk), .SN(n17161), .Q(vis_r4_o[31]), 
        .QN(n5198) );
  DFFS_X1 Ll73z4_reg ( .D(U752_Z_0), .CK(hclk), .SN(n17148), .Q(vis_r2_o[31]), 
        .QN(n5450) );
  DFFS_X1 Kt33z4_reg ( .D(U737_Z_0), .CK(hclk), .SN(n17177), .Q(vis_r9_o[31]), 
        .QN(n5363) );
  DFFS_X1 Koj2z4_reg ( .D(U801_Z_0), .CK(hclk), .SN(n17179), .Q(vis_r1_o[31]), 
        .QN(n4981) );
  DFFS_X1 Isi2z4_reg ( .D(U712_Z_0), .CK(hclk), .SN(n17180), .Q(vis_r7_o[31]), 
        .QN(n4962) );
  DFFS_X1 Glj2z4_reg ( .D(U702_Z_0), .CK(hclk), .SN(n17175), .Q(vis_r5_o[31]), 
        .QN(n4979) );
  DFFS_X1 Ehz2z4_reg ( .D(U717_Z_0), .CK(hclk), .SN(n17186), .Q(vis_r12_o[31]), 
        .QN(n5263) );
  DFFS_X1 Cgt2z4_reg ( .D(U707_Z_0), .CK(hclk), .SN(n17144), .Q(vis_r6_o[31]), 
        .QN(n5169) );
  DFFS_X1 Cc63z4_reg ( .D(U747_Z_0), .CK(hclk), .SN(n17184), .Q(vis_r3_o[31]), 
        .QN(n5421) );
  DFFS_X1 Bk23z4_reg ( .D(U732_Z_0), .CK(hclk), .SN(n17146), .Q(vis_r10_o[31]), 
        .QN(n5334) );
  DFFS_X1 Gci2z4_reg ( .D(U229_Z_0), .CK(hclk), .SN(n17154), .Q(vis_apsr_o[3]), 
        .QN(n4948) );
  DFFS_X1 Igi2z4_reg ( .D(U665_Z_0), .CK(hclk), .SN(n17151), .Q(vis_apsr_o[2]), 
        .QN(n4954) );
  DFFR_X1 Pet2z4_reg ( .D(n4878), .CK(hclk), .RN(hreset_n), .Q(n2029), .QN(
        n4843) );
  DFFR_X1 Y6t2z4_reg ( .D(n4876), .CK(hclk), .RN(n17132), .Q(n808), .QN(n5165)
         );
  DFFR_X1 V3o2z4_reg ( .D(n5712), .CK(hclk), .RN(n17135), .QN(n5068) );
  DFFR_X1 Y9t2z4_reg ( .D(n4886), .CK(hclk), .RN(n17129), .Q(n1063), .QN(n5167) );
  DFFR_X1 Mbt2z4_reg ( .D(n4864), .CK(hclk), .RN(n17133), .Q(n3229), .QN(n4829) );
  DFFR_X1 S5b3z4_reg ( .D(n4874), .CK(hclk), .RN(n17133), .QN(n4833) );
  DFFR_X1 R0t2z4_reg ( .D(n4882), .CK(hclk), .RN(n17130), .Q(n3313), .QN(n4848) );
  DFFR_X1 Adt2z4_reg ( .D(n4863), .CK(hclk), .RN(n17133), .Q(n3059), .QN(n5168) );
  DFFR_X1 Tna3z4_reg ( .D(n4860), .CK(hclk), .RN(n17135), .QN(n5516) );
  DFFR_X1 Bec3z4_reg ( .D(n5696), .CK(hclk), .RN(n17133), .Q(n217), .QN(n4801)
         );
  DFFR_X1 Zad3z4_reg ( .D(U766_Z_0), .CK(hclk), .RN(n17138), .Q(n3847), .QN(
        n5549) );
  DFFR_X1 Bmb3z4_reg ( .D(U774_Z_0), .CK(hclk), .RN(n17138), .QN(n5523) );
  DFFR_X1 Kkb3z4_reg ( .D(U782_Z_0), .CK(hclk), .RN(n17138), .Q(n3812), .QN(
        n5522) );
  DFFR_X1 Tib3z4_reg ( .D(U790_Z_0), .CK(hclk), .RN(n17137), .Q(n3784), .QN(
        n5521) );
  DFFR_X1 Mcc3z4_reg ( .D(n5695), .CK(hclk), .RN(n17133), .Q(n214), .QN(n5535)
         );
  DFFR_X1 Fhc3z4_reg ( .D(n5698), .CK(hclk), .RN(n17133), .Q(n223), .QN(n4800)
         );
  DFFR_X1 Ztc3z4_reg ( .D(n5710), .CK(hclk), .RN(n17135), .QN(n5540) );
  DFFR_X1 U5x2z4_reg ( .D(n5826), .CK(hclk), .RN(n17131), .QN(n5234) );
  DFFR_X1 Qfc3z4_reg ( .D(n5697), .CK(hclk), .RN(n17133), .Q(n220), .QN(n5536)
         );
  DFFR_X1 X9n2z4_reg ( .D(n4854), .CK(hclk), .RN(n17136), .Q(n2889), .QN(n4826) );
  DFFR_X1 Ylc3z4_reg ( .D(n5701), .CK(hclk), .RN(n17137), .Q(n231), .QN(n4797)
         );
  DFFR_X1 J9d3z4_reg ( .D(U767_Z_0), .CK(hclk), .RN(n17136), .Q(n2951), .QN(
        n5548) );
  DFFR_X1 Xdb3z4_reg ( .D(U775_Z_0), .CK(hclk), .RN(n17136), .Q(n2952), .QN(
        n5519) );
  DFFR_X1 Gcb3z4_reg ( .D(U783_Z_0), .CK(hclk), .RN(n17135), .QN(n5518) );
  DFFR_X1 G8n2z4_reg ( .D(U771_Z_0), .CK(hclk), .RN(n17137), .Q(n4367), .QN(
        n5053) );
  DFFR_X1 Bus2z4_reg ( .D(U779_Z_0), .CK(hclk), .RN(n17137), .Q(n2888), .QN(
        n5158) );
  DFFR_X1 Dks2z4_reg ( .D(U787_Z_0), .CK(hclk), .RN(n17137), .Q(n2890), .QN(
        n5152) );
  DFFR_X1 Jkc3z4_reg ( .D(n5700), .CK(hclk), .RN(n17135), .Q(n228), .QN(n4798)
         );
  DFFR_X1 Uqi2z4_reg ( .D(n5652), .CK(hclk), .RN(n17130), .Q(n3731), .QN(n4961) );
  DFFR_X1 Aqp2z4_reg ( .D(n4883), .CK(hclk), .RN(n17130), .Q(n2929), .QN(n5097) );
  DFFR_X1 B1a3z4_reg ( .D(n4862), .CK(hclk), .RN(n17134), .QN(n5503) );
  DFFR_X1 Vfd3z4_reg ( .D(U762_Z_0), .CK(hclk), .RN(n17129), .Q(n3834), .QN(
        n5551) );
  DFFR_X1 Z4l2z4_reg ( .D(U770_Z_0), .CK(hclk), .RN(n17134), .Q(n3863), .QN(
        n5008) );
  DFFR_X1 Svs2z4_reg ( .D(U778_Z_0), .CK(hclk), .RN(n17134), .Q(n3793), .QN(
        n5159) );
  DFFR_X1 Uls2z4_reg ( .D(U786_Z_0), .CK(hclk), .RN(n17134), .Q(n3790), .QN(
        n5153) );
  DFFR_X1 Lns2z4_reg ( .D(U785_Z_0), .CK(hclk), .RN(n17134), .Q(n2927), .QN(
        n5154) );
  DFFR_X1 Lhd3z4_reg ( .D(U761_Z_0), .CK(hclk), .RN(n17129), .Q(n2933), .QN(
        n5552) );
  DFFR_X1 Q6l2z4_reg ( .D(U769_Z_0), .CK(hclk), .RN(n17134), .Q(n2931), .QN(
        n5009) );
  DFFR_X1 Jxs2z4_reg ( .D(U777_Z_0), .CK(hclk), .RN(n17134), .Q(n2932), .QN(
        n5160) );
  DFFR_X1 Wbk2z4_reg ( .D(n5694), .CK(hclk), .RN(n17128), .Q(n209), .QN(n4802)
         );
  DFFR_X1 Yvb3z4_reg ( .D(n13951), .CK(hclk), .RN(n17131), .QN(n5527) );
  DFFR_X1 Qsb3z4_reg ( .D(n13963), .CK(hclk), .RN(n17135), .QN(n5525) );
  DFFR_X1 Vve3z4_reg ( .D(n5703), .CK(hclk), .RN(n17138), .QN(n5578) );
  DFFR_X1 Rnb3z4_reg ( .D(n13894), .CK(hclk), .RN(n17132), .QN(n5524) );
  DFFR_X1 T7d3z4_reg ( .D(U764_Z_0), .CK(hclk), .RN(n17138), .Q(n3719), .QN(
        n5547) );
  DFFR_X1 Usl2z4_reg ( .D(U772_Z_0), .CK(hclk), .RN(n17138), .Q(n3720), .QN(
        n5023) );
  DFFR_X1 Tqs2z4_reg ( .D(U780_Z_0), .CK(hclk), .RN(n17138), .Q(n3813), .QN(
        n5156) );
  DFFR_X1 Vgs2z4_reg ( .D(U788_Z_0), .CK(hclk), .RN(n17138), .Q(n4356), .QN(
        n5150) );
  DFFR_X1 Pcd3z4_reg ( .D(U765_Z_0), .CK(hclk), .RN(n17136), .Q(n2901), .QN(
        n5550) );
  DFFR_X1 Axm2z4_reg ( .D(U773_Z_0), .CK(hclk), .RN(n17136), .Q(n2902), .QN(
        n5046) );
  DFFR_X1 Kss2z4_reg ( .D(U781_Z_0), .CK(hclk), .RN(n17137), .QN(n5157) );
  DFFR_X1 Mis2z4_reg ( .D(U789_Z_0), .CK(hclk), .RN(n17136), .QN(n5151) );
  DFFR_X1 Lee3z4_reg ( .D(n5705), .CK(hclk), .RN(n17133), .QN(n5570) );
  DFFR_X1 Gzb3z4_reg ( .D(n13932), .CK(hclk), .RN(n17137), .QN(n5529) );
  DFFR_X1 Hzj2z4_reg ( .D(n5693), .CK(hclk), .RN(n17129), .Q(n203), .QN(n4988)
         );
  DFFR_X1 Aok2z4_reg ( .D(n10055), .CK(hclk), .RN(n17129), .Q(n16846), .QN(
        n16844) );
  DFFR_X1 Nnc3z4_reg ( .D(n5704), .CK(hclk), .RN(n17133), .QN(n5537) );
  DFFR_X1 H2f3z4_reg ( .D(n5702), .CK(hclk), .RN(n17137), .QN(n4796) );
  DFFR_X1 N7c3z4_reg ( .D(n11945), .CK(hclk), .RN(n17132), .Q(n3861), .QN(
        n5533) );
  DFFR_X1 Pxb3z4_reg ( .D(n4894), .CK(hclk), .RN(n17131), .Q(n3238), .QN(n5528) );
  DFFR_X1 Jsc3z4_reg ( .D(n5709), .CK(hclk), .RN(n17139), .Q(n3785), .QN(n5539) );
  DFFR_X1 Vac3z4_reg ( .D(n11939), .CK(hclk), .RN(n17136), .QN(n5534) );
  DFFR_X1 Tqc3z4_reg ( .D(n5708), .CK(hclk), .RN(n17136), .Q(n2916), .QN(n5538) );
  DFFR_X1 Dpc3z4_reg ( .D(n5706), .CK(hclk), .RN(n17133), .QN(n4795) );
  DFFR_X1 Gxk2z4_reg ( .D(n11929), .CK(hclk), .RN(n17139), .QN(n5005) );
  DFFR_X1 Hub3z4_reg ( .D(n4893), .CK(hclk), .RN(n17131), .Q(n3107), .QN(n5526) );
  DFFR_X1 O2c3z4_reg ( .D(n13919), .CK(hclk), .RN(n17135), .QN(n5531) );
  DFFR_X1 Ipb3z4_reg ( .D(n4901), .CK(hclk), .RN(n17132), .Q(n3060), .QN(n4750) );
  DFFR_X1 X0c3z4_reg ( .D(n4899), .CK(hclk), .RN(n17137), .QN(n5530) );
  DFFR_X1 Q0f3z4_reg ( .D(n4904), .CK(hclk), .RN(n17139), .Q(n1129), .QN(n5580) );
  DFFR_X1 Qnn2z4_reg ( .D(n13835), .CK(hclk), .RN(n17128), .QN(n5061) );
  DFFR_X1 Etq2z4_reg ( .D(n13989), .CK(hclk), .RN(n17132), .QN(n5118) );
  DFFR_X1 C7f3z4_reg ( .D(n13813), .CK(hclk), .RN(n17137), .QN(n5582) );
  DFFR_X1 Fij2z4_reg ( .D(n5781), .CK(hclk), .RN(n17131), .Q(n16852), .QN(
        n16850) );
  DFFR_X1 W8r2z4_reg ( .D(n13795), .CK(hclk), .RN(n17132), .Q(n4333), .QN(
        n5126) );
  DFFR_X1 Uyv2z4_reg ( .D(n5825), .CK(hclk), .RN(n17136), .Q(n1053) );
  DFFR_X1 F4c3z4_reg ( .D(n4898), .CK(hclk), .RN(n17135), .Q(n2953), .QN(n5532) );
  DFFR_X1 Qrp2z4_reg ( .D(n5651), .CK(hclk), .RN(n17130), .Q(n3740), .QN(n5098) );
  DFFR_X1 Cps2z4_reg ( .D(U784_Z_0), .CK(hclk), .RN(n17134), .Q(n3791), .QN(
        n5155) );
  DFFR_X1 Bjd3z4_reg ( .D(U760_Z_0), .CK(hclk), .RN(n17134), .Q(n3833), .QN(
        n5553) );
  DFFR_X1 H8l2z4_reg ( .D(U768_Z_0), .CK(hclk), .RN(n17134), .Q(n3862), .QN(
        n5010) );
  DFFR_X1 Azs2z4_reg ( .D(U776_Z_0), .CK(hclk), .RN(n17134), .Q(n3792), .QN(
        n5161) );
  DFFR_X1 P2a3z4_reg ( .D(n5650), .CK(hclk), .RN(n17134), .Q(n3732), .QN(n5504) );
  DFFR_X1 Nsk2z4_reg ( .D(n9796), .CK(hclk), .RN(n17130), .Q(n16690), .QN(
        n16827) );
  DFFR_X1 Npk2z4_reg ( .D(n9972), .CK(hclk), .RN(n17131), .Q(n16728), .QN(
        n16840) );
  DFFR_X1 Oar2z4_reg ( .D(n4900), .CK(hclk), .RN(n17128), .Q(n3089), .QN(n4749) );
  DFFR_X1 Y9l2z4_reg ( .D(n11957), .CK(hclk), .RN(n17137), .QN(n5011) );
  DFFR_X1 Ble3z4_reg ( .D(n11971), .CK(hclk), .RN(n17128), .QN(n5572) );
  DFFR_X1 I6h3z4_reg ( .D(n14001), .CK(hclk), .RN(n17138), .Q(n1379), .QN(
        n5620) );
  DFFR_X1 Mvi2z4_reg ( .D(n13870), .CK(hclk), .RN(n17138), .QN(n4964) );
  DFFR_X1 Ipn2z4_reg ( .D(n4903), .CK(hclk), .RN(n17128), .QN(n4748) );
  DFFR_X1 T8f3z4_reg ( .D(n4902), .CK(hclk), .RN(n17136), .QN(n4747) );
  DFFR_X1 Lul2z4_reg ( .D(n4895), .CK(hclk), .RN(n17138), .Q(n3786), .QN(n5024) );
  DFFR_X1 Rym2z4_reg ( .D(n4896), .CK(hclk), .RN(n17136), .Q(n2914), .QN(n5047) );
  DFFR_X1 Ywi2z4_reg ( .D(n11928), .CK(hclk), .RN(n17129), .Q(n1066), .QN(
        n4965) );
  DFFR_X1 Q4h3z4_reg ( .D(n13747), .CK(hclk), .RN(n17136), .QN(n5619) );
  DFFR_X1 Ark2z4_reg ( .D(n5777), .CK(hclk), .RN(n17130), .Q(n16835), .QN(
        n16834) );
  DFFR_X1 U7w2z4_reg ( .D(n5799), .CK(hclk), .RN(n17139), .Q(n3066), .QN(n5229) );
  DFFR_X1 Ffj2z4_reg ( .D(n5789), .CK(hclk), .RN(n17129), .Q(n16863), .QN(
        n16861) );
  DFFR_X1 Sgj2z4_reg ( .D(n5774), .CK(hclk), .RN(n17130), .Q(n16694), .QN(
        n16857) );
  DFFR_X1 C3w2z4_reg ( .D(U802_Z_0), .CK(hclk), .RN(n17135), .Q(n3222), .QN(
        n5227) );
  DFFR_X1 Vaw2z4_reg ( .D(n5795), .CK(hclk), .RN(n17130), .Q(n375), .QN(n5231)
         );
  DFFR_X1 Wxp2z4_reg ( .D(U518_Z_0), .CK(hclk), .RN(n17128), .Q(n3223), .QN(
        n5102) );
  DFFR_X1 Gji2z4_reg ( .D(U227_Z_0), .CK(hclk), .RN(n17128), .Q(n1096), .QN(
        n4956) );
  DFFR_X1 L8t2z4_reg ( .D(n5823), .CK(hclk), .RN(n17131), .Q(n16681), .QN(
        n16822) );
  DFFR_X1 Aii3z4_reg ( .D(n4875), .CK(hclk), .RN(n17132), .QN(n4834) );
  DFFR_X1 Jhy2z4_reg ( .D(n5796), .CK(hclk), .RN(n17131), .Q(n1002) );
  DFFR_X1 Kop2z4_reg ( .D(n5792), .CK(hclk), .RN(n17129), .Q(n3874), .QN(n5096) );
  DFFR_X1 Mjl2z4_reg ( .D(n5793), .CK(hclk), .RN(n17128), .Q(n3875), .QN(n5017) );
  DFFR_X1 Tki2z4_reg ( .D(n5775), .CK(hclk), .RN(n17128), .Q(n16689), .QN(
        n16872) );
  DFFS_X1 O5t2z4_reg ( .D(n5778), .CK(hclk), .SN(n17190), .Q(n16805), .QN(
        n16806) );
  DFFS_X1 Sjj2z4_reg ( .D(U134_Z_0), .CK(hclk), .SN(n17142), .Q(n3488), .QN(
        n4978) );
  DFFS_X1 Fgm2z4_reg ( .D(U121_Z_0), .CK(hclk), .SN(n17190), .Q(n3480), .QN(
        n5036) );
  DFFS_X1 Cyq2z4_reg ( .D(n5780), .CK(hclk), .SN(n17154), .Q(n16671), .QN(
        n16810) );
  DFFS_X1 Zcn2z4_reg ( .D(U756_Z_0), .CK(hclk), .SN(n17154), .Q(n16656), .QN(
        n16809) );
  DFFS_X1 Yzi2z4_reg ( .D(n5752), .CK(hclk), .SN(n17159), .Q(n451), .QN(n4967)
         );
  DFFS_X1 Xly2z4_reg ( .D(n5748), .CK(hclk), .SN(n17159), .Q(n781), .QN(n5243)
         );
  DFFS_X1 Lny2z4_reg ( .D(n5747), .CK(hclk), .SN(n17159), .Q(n659), .QN(n5244)
         );
  DFFS_X1 Bsy2z4_reg ( .D(n5744), .CK(hclk), .SN(n17140), .Q(n16686), .QN(
        n16797) );
  DFFS_X1 Pdi2z4_reg ( .D(n11746), .CK(hclk), .SN(n17151), .Q(n1697), .QN(
        n4950) );
  DFFS_X2 Pty2z4_reg ( .D(n5743), .CK(hclk), .SN(n17139), .Q(n16657), .QN(
        n16796) );
  DFFS_X2 Qem2z4_reg ( .D(n5753), .CK(hclk), .SN(n17158), .Q(n16683), .QN(
        n16807) );
  DFFS_X2 U2x2z4_reg ( .D(n5754), .CK(hclk), .SN(n17151), .Q(n16659), .QN(
        n16811) );
  DFFS_X2 Zoy2z4_reg ( .D(n5746), .CK(hclk), .SN(n17139), .Q(n16674), .QN(
        n16801) );
  DFFR_X2 K3l2z4_reg ( .D(U792_Z_0), .CK(hclk), .RN(n17128), .Q(n253), .QN(
        n5007) );
  DFFS_X2 Jky2z4_reg ( .D(n5749), .CK(hclk), .SN(n17141), .Q(n16734), .QN(
        n16794) );
  DFFS_X2 Hyy2z4_reg ( .D(n5740), .CK(hclk), .SN(n17139), .Q(n16725), .QN(
        n16795) );
  DFFS_X2 Swy2z4_reg ( .D(n5741), .CK(hclk), .SN(n17140), .Q(n16733), .QN(
        n16814) );
  DFFR_X2 A4t2z4_reg ( .D(n5794), .CK(hclk), .RN(n17130), .Q(n16808), .QN(
        n16680) );
  DFFS_X2 Nqy2z4_reg ( .D(n5745), .CK(hclk), .SN(n17140), .Q(n16798), .QN(
        n16800) );
  DFFR_X2 Emi2z4_reg ( .D(n10553), .CK(hclk), .RN(n17129), .Q(n16867), .QN(
        n16865) );
  DFFS_X2 H9i2z4_reg ( .D(n5739), .CK(hclk), .SN(n17159), .Q(n16802), .QN(
        n16803) );
  OR2_X4 U108 ( .A1(n42), .A2(n187), .ZN(n16644) );
  NOR2_X4 U112 ( .A1(n2998), .A2(n16789), .ZN(n16645) );
  NOR3_X4 U124 ( .A1(n376), .A2(n374), .A3(n377), .ZN(n16646) );
  OR3_X4 U135 ( .A1(n17108), .A2(n258), .A3(n314), .ZN(n16647) );
  AND2_X4 U137 ( .A1(n4665), .A2(n4663), .ZN(n16648) );
  AND2_X4 U141 ( .A1(n4661), .A2(n4659), .ZN(n16649) );
  AND2_X4 U144 ( .A1(n4665), .A2(n4661), .ZN(n16650) );
  AND3_X4 U145 ( .A1(n4660), .A2(n4662), .A3(n4968), .ZN(n16651) );
  AND2_X4 U159 ( .A1(n4660), .A2(n4658), .ZN(n16652) );
  XOR2_X2 U190 ( .A(add_2073_A_13_), .B(n16714), .Z(n16653) );
  AND2_X4 U191 ( .A1(add_2073_A_30_), .A2(n16661), .ZN(n16654) );
  NAND2_X2 U197 ( .A1(n1697), .A2(n4676), .ZN(n2169) );
  XOR2_X2 U200 ( .A(add_2073_A_26_), .B(n16665), .Z(n16655) );
  XOR2_X2 U213 ( .A(add_2073_A_15_), .B(n16707), .Z(n16658) );
  OAI22_X2 U224 ( .A1(n4401), .A2(n2196), .B1(n16786), .B2(n2254), .ZN(n247)
         );
  AND2_X4 U227 ( .A1(add_2073_A_31_), .A2(n16654), .ZN(n16660) );
  AND2_X4 U236 ( .A1(add_2073_A_29_), .A2(n16692), .ZN(n16661) );
  AND2_X4 U239 ( .A1(add_2073_A_27_), .A2(n16697), .ZN(n16662) );
  XOR2_X2 U242 ( .A(add_2073_A_27_), .B(n16697), .Z(n16663) );
  AND2_X4 U250 ( .A1(add_2073_A_23_), .A2(n16700), .ZN(n16664) );
  AND2_X4 U251 ( .A1(add_2073_A_25_), .A2(n16696), .ZN(n16665) );
  AND2_X4 U253 ( .A1(add_2073_A_17_), .A2(n16708), .ZN(n16666) );
  AND2_X4 U254 ( .A1(add_2073_A_20_), .A2(n16704), .ZN(n16667) );
  XOR2_X2 U260 ( .A(add_2073_A_22_), .B(n16699), .Z(n16668) );
  AND2_X4 U267 ( .A1(add_2073_A_15_), .A2(n16707), .ZN(n16669) );
  AND2_X4 U270 ( .A1(add_2073_A_13_), .A2(n16714), .ZN(n16670) );
  XOR2_X2 U273 ( .A(add_2073_A_19_), .B(n16703), .Z(n16672) );
  AND2_X4 U276 ( .A1(add_2073_A_9_), .A2(n16718), .ZN(n16673) );
  XOR2_X2 U279 ( .A(add_2082_B_1_), .B(add_2082_A_1_), .Z(n16675) );
  AND2_X4 U282 ( .A1(add_2073_A_5_), .A2(n16717), .ZN(n16676) );
  AND2_X4 U285 ( .A1(add_2073_A_6_), .A2(n16676), .ZN(n16677) );
  AND2_X4 U288 ( .A1(add_2073_A_3_), .A2(n16721), .ZN(n16678) );
  XOR2_X2 U291 ( .A(add_2073_A_14_), .B(n16670), .Z(n16679) );
  XOR2_X2 U294 ( .A(add_2073_A_4_), .B(n16678), .Z(n16682) );
  XOR2_X2 U297 ( .A(n4068), .B(n4168), .Z(n16684) );
  OR3_X4 U300 ( .A1(n2926), .A2(n4905), .A3(n261), .ZN(n16685) );
  XOR2_X2 U303 ( .A(add_2073_A_32_), .B(n16660), .Z(n16688) );
  AND2_X4 U306 ( .A1(add_2082_B_1_), .A2(add_2082_A_1_), .ZN(n16691) );
  AND2_X4 U309 ( .A1(add_2073_A_28_), .A2(n16662), .ZN(n16692) );
  XOR2_X2 U312 ( .A(add_2073_A_30_), .B(n16661), .Z(n16693) );
  XOR2_X2 U313 ( .A(add_2073_A_29_), .B(n16692), .Z(n16695) );
  AND2_X4 U315 ( .A1(add_2073_A_24_), .A2(n16664), .ZN(n16696) );
  AND2_X4 U316 ( .A1(add_2073_A_26_), .A2(n16665), .ZN(n16697) );
  XOR2_X2 U319 ( .A(add_2073_A_28_), .B(n16662), .Z(n16698) );
  AND2_X4 U353 ( .A1(add_2073_A_21_), .A2(n16667), .ZN(n16699) );
  AND2_X4 U359 ( .A1(add_2073_A_22_), .A2(n16699), .ZN(n16700) );
  XOR2_X2 U468 ( .A(add_2073_A_25_), .B(n16696), .Z(n16701) );
  XOR2_X2 U512 ( .A(add_2073_A_23_), .B(n16700), .Z(n16702) );
  AND2_X4 U582 ( .A1(add_2073_A_18_), .A2(n16666), .ZN(n16703) );
  AND2_X4 U648 ( .A1(add_2073_A_19_), .A2(n16703), .ZN(n16704) );
  XOR2_X2 U711 ( .A(add_2073_A_24_), .B(n16664), .Z(n16705) );
  XOR2_X2 U742 ( .A(add_2073_A_21_), .B(n16667), .Z(n16706) );
  AND2_X4 U751 ( .A1(add_2073_A_14_), .A2(n16670), .ZN(n16707) );
  AND2_X4 U752 ( .A1(add_2073_A_16_), .A2(n16669), .ZN(n16708) );
  XOR2_X2 U753 ( .A(add_2073_A_20_), .B(n16704), .Z(n16709) );
  XOR2_X2 U754 ( .A(add_2073_A_18_), .B(n16666), .Z(n16710) );
  XOR2_X2 U756 ( .A(add_2073_A_17_), .B(n16708), .Z(n16711) );
  AND2_X4 U757 ( .A1(add_2073_A_10_), .A2(n16673), .ZN(n16712) );
  AND2_X4 U758 ( .A1(add_2073_A_11_), .A2(n16712), .ZN(n16713) );
  AND2_X4 U759 ( .A1(add_2073_A_12_), .A2(n16713), .ZN(n16714) );
  XOR2_X2 U785 ( .A(add_2073_A_16_), .B(n16669), .Z(n16715) );
  AND2_X4 U812 ( .A1(add_2073_A_7_), .A2(n16677), .ZN(n16716) );
  AND2_X4 U820 ( .A1(add_2073_A_4_), .A2(n16678), .ZN(n16717) );
  AND2_X4 U837 ( .A1(add_2073_A_8_), .A2(n16716), .ZN(n16718) );
  XOR2_X2 U840 ( .A(add_2073_A_12_), .B(n16713), .Z(n16719) );
  AND2_X4 U841 ( .A1(add_2073_B_1_), .A2(n16675), .ZN(n16720) );
  AND2_X4 U845 ( .A1(add_2073_A_2_), .A2(n16720), .ZN(n16721) );
  XOR2_X2 U850 ( .A(add_2073_A_9_), .B(n16718), .Z(n16722) );
  XOR2_X2 U851 ( .A(add_2073_A_11_), .B(n16712), .Z(n16723) );
  OR2_X4 U852 ( .A1(n16736), .A2(n16737), .ZN(haddr_o[15]) );
  NAND3_X2 U856 ( .A1(n373), .A2(n379), .A3(n400), .ZN(n381) );
  XOR2_X2 U857 ( .A(add_2073_A_8_), .B(n16716), .Z(n16726) );
  XOR2_X2 U858 ( .A(add_2073_A_10_), .B(n16673), .Z(n16727) );
  NOR2_X2 U879 ( .A1(n4131), .A2(n4130), .ZN(n3118) );
  XOR2_X2 U880 ( .A(add_2073_A_3_), .B(n16721), .Z(n16729) );
  XOR2_X2 U996 ( .A(add_2073_A_5_), .B(n16717), .Z(n16730) );
  XOR2_X2 U997 ( .A(add_2073_A_6_), .B(n16676), .Z(n16731) );
  NOR2_X2 U1000 ( .A1(n4142), .A2(n4131), .ZN(n3275) );
  XOR2_X2 U1006 ( .A(add_2073_A_2_), .B(n16720), .Z(n16732) );
  NAND4_X2 U1013 ( .A1(n2674), .A2(n2675), .A3(n2676), .A4(n2677), .ZN(n979)
         );
  OAI22_X2 U1022 ( .A1(n4401), .A2(n2250), .B1(n16786), .B2(n2253), .ZN(n245)
         );
  NAND2_X1 U1024 ( .A1(n5649), .A2(n422), .ZN(n16735) );
  OAI21_X2 U1027 ( .B1(n2643), .B2(n2644), .A(n979), .ZN(n1632) );
  OAI221_X2 U1031 ( .B1(n16845), .B2(n1086), .C1(n16862), .C2(n715), .A(n2645), 
        .ZN(n2644) );
  NOR2_X1 U1051 ( .A1(n1661), .A2(n1622), .ZN(n16736) );
  INV_X1 U1054 ( .A(n1662), .ZN(n16737) );
  OAI21_X4 U1112 ( .B1(n2626), .B2(n2627), .A(n979), .ZN(n1622) );
  INV_X4 U1259 ( .A(n876), .ZN(haddr_o[2]) );
  AOI221_X2 U1260 ( .B1(n16729), .B2(n17086), .C1(n1640), .C2(n1628), .A(n1641), .ZN(n876) );
  OAI221_X4 U1264 ( .B1(n1654), .B2(n1622), .C1(n1655), .C2(n1632), .A(n1656), 
        .ZN(haddr_o[19]) );
  NAND4_X2 U1265 ( .A1(n1603), .A2(n4588), .A3(n4589), .A4(n4590), .ZN(n1612)
         );
  XOR2_X2 U1266 ( .A(n16990), .B(n3407), .Z(n5818) );
  NOR2_X2 U1267 ( .A1(n1614), .A2(n5167), .ZN(n4240) );
  INV_X4 U1270 ( .A(n968), .ZN(haddr_o[5]) );
  AOI221_X2 U1271 ( .B1(n1634), .B2(n1628), .C1(n16731), .C2(n17087), .A(n1635), .ZN(n968) );
  OAI21_X4 U1273 ( .B1(n1695), .B2(n1622), .A(n1731), .ZN(haddr_o[11]) );
  XOR2_X2 U1275 ( .A(n16990), .B(n2730), .Z(n5815) );
  INV_X4 U1278 ( .A(n4260), .ZN(hwdata_o[31]) );
  INV_X4 U1280 ( .A(n24), .ZN(hwdata_o[26]) );
  INV_X4 U1281 ( .A(n967), .ZN(haddr_o[4]) );
  AOI221_X2 U1283 ( .B1(n1636), .B2(n1628), .C1(n16730), .C2(n17087), .A(n1637), .ZN(n967) );
  OAI22_X4 U1284 ( .A1(n1607), .A2(n1608), .B1(n1609), .B2(n999), .ZN(
        htrans_o[1]) );
  NOR3_X4 U1286 ( .A1(n1614), .A2(n17090), .A3(n1613), .ZN(hsize_o[0]) );
  OAI221_X4 U1288 ( .B1(n1630), .B2(n1622), .C1(n16782), .C2(n1632), .A(n1633), 
        .ZN(haddr_o[6]) );
  XOR2_X2 U1289 ( .A(n2169), .B(n3035), .Z(n5807) );
  INV_X4 U1294 ( .A(n1149), .ZN(haddr_o[26]) );
  AOI221_X2 U1296 ( .B1(n1645), .B2(n1628), .C1(n16663), .C2(n17087), .A(n1646), .ZN(n1149) );
  INV_X4 U1297 ( .A(n1158), .ZN(haddr_o[17]) );
  AOI221_X2 U1299 ( .B1(n1658), .B2(n1628), .C1(n16710), .C2(n17087), .A(n1659), .ZN(n1158) );
  INV_X4 U1301 ( .A(n208), .ZN(hwdata_o[27]) );
  INV_X4 U1303 ( .A(n1155), .ZN(haddr_o[20]) );
  OAI21_X2 U1305 ( .B1(n3218), .B2(n3213), .A(n2756), .ZN(n2004) );
  INV_X4 U1307 ( .A(n4272), .ZN(hwdata_o[29]) );
  INV_X4 U1308 ( .A(n948), .ZN(haddr_o[10]) );
  AOI221_X2 U1310 ( .B1(n1667), .B2(n1628), .C1(n16723), .C2(n17087), .A(n1668), .ZN(n948) );
  NAND2_X2 U1312 ( .A1(n1620), .A2(n1869), .ZN(haddr_o[29]) );
  OAI21_X4 U1313 ( .B1(n1621), .B2(n1622), .A(n1623), .ZN(haddr_o[9]) );
  OAI22_X2 U1315 ( .A1(n2461), .A2(n4610), .B1(n2462), .B2(n3534), .ZN(
        U186_Z_0) );
  XOR2_X2 U1317 ( .A(n16990), .B(n3356), .Z(n5819) );
  INV_X4 U1318 ( .A(n1116), .ZN(hwdata_o[21]) );
  AOI22_X2 U1320 ( .A1(n4202), .A2(n2556), .B1(n21), .B2(n4203), .ZN(n1116) );
  INV_X4 U1322 ( .A(n1148), .ZN(haddr_o[27]) );
  INV_X4 U1324 ( .A(n1157), .ZN(haddr_o[18]) );
  INV_X4 U1326 ( .A(n205), .ZN(hwdata_o[28]) );
  INV_X4 U1328 ( .A(n1112), .ZN(hwdata_o[17]) );
  AOI22_X2 U1329 ( .A1(n4202), .A2(n2028), .B1(n2258), .B2(n4203), .ZN(n1112)
         );
  INV_X4 U1331 ( .A(n25), .ZN(hwdata_o[24]) );
  INV_X4 U1332 ( .A(n1154), .ZN(haddr_o[21]) );
  AOI221_X2 U1334 ( .B1(n1651), .B2(n1628), .C1(n16668), .C2(n17087), .A(n1652), .ZN(n1154) );
  OAI21_X2 U1367 ( .B1(n1168), .B2(n1169), .A(n17125), .ZN(n866) );
  OAI211_X2 U1396 ( .C1(n650), .C2(n912), .A(n1170), .B(n1171), .ZN(n1169) );
  NAND4_X2 U1402 ( .A1(n1875), .A2(n1876), .A3(n1877), .A4(n1878), .ZN(
        hwrite_o) );
  OAI21_X2 U1465 ( .B1(n3427), .B2(n3213), .A(n2756), .ZN(n2871) );
  NOR3_X4 U1466 ( .A1(n1612), .A2(n683), .A3(n1613), .ZN(haddr_o[1]) );
  AOI222_X2 U1500 ( .A1(n17090), .A2(n2625), .B1(n16732), .B2(n17087), .C1(
        n2232), .C2(n1628), .ZN(n683) );
  OAI211_X2 U1501 ( .C1(n3242), .C2(n3243), .A(n3244), .B(n3245), .ZN(n2011)
         );
  INV_X4 U1509 ( .A(n1077), .ZN(hwdata_o[30]) );
  AOI222_X2 U1512 ( .A1(n2250), .A2(n16786), .B1(n2253), .B2(n4240), .C1(n2083), .C2(n4203), .ZN(n1077) );
  OAI21_X4 U1519 ( .B1(n1616), .B2(n1617), .A(hprot_o[2]), .ZN(hprot_o[3]) );
  OAI21_X4 U1521 ( .B1(n1638), .B2(n1622), .A(n1639), .ZN(haddr_o[3]) );
  NOR2_X2 U1524 ( .A1(n3962), .A2(n2926), .ZN(n2895) );
  NAND2_X2 U1529 ( .A1(n1759), .A2(n4172), .ZN(n2926) );
  INV_X4 U1531 ( .A(n4261), .ZN(hwdata_o[23]) );
  AOI22_X2 U1533 ( .A1(n3450), .A2(n4203), .B1(n4202), .B2(n2196), .ZN(n4261)
         );
  INV_X4 U1546 ( .A(n1115), .ZN(hwdata_o[18]) );
  AOI22_X2 U1551 ( .A1(n4202), .A2(n3177), .B1(n2249), .B2(n4203), .ZN(n1115)
         );
  INV_X4 U1561 ( .A(n955), .ZN(hsize_o[1]) );
  AOI21_X2 U1571 ( .B1(n1612), .B2(n979), .A(n1613), .ZN(n955) );
  INV_X4 U1581 ( .A(n1117), .ZN(hwdata_o[20]) );
  AOI22_X2 U1598 ( .A1(n4202), .A2(n2578), .B1(n20), .B2(n4203), .ZN(n1117) );
  INV_X4 U1604 ( .A(n1118), .ZN(hwdata_o[16]) );
  AOI22_X2 U1607 ( .A1(n4202), .A2(n1354), .B1(n17), .B2(n4203), .ZN(n1118) );
  INV_X4 U1761 ( .A(n973), .ZN(haddr_o[23]) );
  INV_X4 U1767 ( .A(n952), .ZN(haddr_o[12]) );
  AOI221_X2 U1775 ( .B1(n1665), .B2(n1628), .C1(n16653), .C2(n17087), .A(n1666), .ZN(n952) );
  INV_X4 U1776 ( .A(n317), .ZN(haddr_o[24]) );
  INV_X4 U1807 ( .A(n956), .ZN(haddr_o[14]) );
  INV_X4 U1813 ( .A(n957), .ZN(haddr_o[13]) );
  INV_X4 U1818 ( .A(n240), .ZN(hwdata_o[12]) );
  AOI22_X2 U1835 ( .A1(n2578), .A2(n16786), .B1(n4401), .B2(n2247), .ZN(n240)
         );
  INV_X4 U1900 ( .A(n185), .ZN(lockup_o) );
  NOR2_X2 U1948 ( .A1(n1861), .A2(n1862), .ZN(n185) );
  INV_X4 U1950 ( .A(n1114), .ZN(hwdata_o[19]) );
  AOI22_X2 U1951 ( .A1(n4202), .A2(n2257), .B1(n22), .B2(n4203), .ZN(n1114) );
  INV_X4 U1953 ( .A(n1150), .ZN(haddr_o[25]) );
  INV_X4 U1962 ( .A(n1159), .ZN(haddr_o[16]) );
  INV_X4 U1964 ( .A(n201), .ZN(hwdata_o[25]) );
  INV_X4 U1965 ( .A(n1153), .ZN(haddr_o[22]) );
  OR2_X4 U1967 ( .A1(haddr_o[29]), .A2(haddr_o[30]), .ZN(hprot_o[2]) );
  OAI221_X4 U2016 ( .B1(n1677), .B2(n1622), .C1(n16783), .C2(n1632), .A(n1874), 
        .ZN(haddr_o[30]) );
  AOI22_X2 U2019 ( .A1(n2260), .A2(n2461), .B1(n2462), .B2(n2463), .ZN(n4952)
         );
  NOR2_X2 U2026 ( .A1(n4834), .A2(n16821), .ZN(sleeping_o) );
  INV_X4 U2028 ( .A(n221), .ZN(hwdata_o[4]) );
  NAND2_X2 U2029 ( .A1(n2578), .A2(n1063), .ZN(n221) );
  OAI221_X2 U2031 ( .B1(n3754), .B2(n3760), .C1(n3761), .C2(n3762), .A(n3763), 
        .ZN(n2909) );
  INV_X4 U2033 ( .A(n229), .ZN(hwdata_o[7]) );
  INV_X4 U2034 ( .A(n224), .ZN(hwdata_o[5]) );
  NAND2_X2 U2056 ( .A1(n2556), .A2(n1063), .ZN(n224) );
  INV_X4 U2066 ( .A(n218), .ZN(hwdata_o[3]) );
  NAND2_X2 U2068 ( .A1(n2257), .A2(n1063), .ZN(n218) );
  INV_X4 U2069 ( .A(n226), .ZN(hwdata_o[6]) );
  INV_X4 U2071 ( .A(n210), .ZN(hwdata_o[1]) );
  NAND2_X2 U2073 ( .A1(n2028), .A2(n1063), .ZN(n210) );
  INV_X4 U2091 ( .A(n249), .ZN(hwdata_o[0]) );
  NAND2_X2 U2099 ( .A1(n1354), .A2(n1063), .ZN(n249) );
  INV_X4 U2101 ( .A(n878), .ZN(haddr_o[28]) );
  AOI221_X2 U2102 ( .B1(n1832), .B2(n1628), .C1(n16695), .C2(n17087), .A(n1833), .ZN(n878) );
  INV_X4 U2104 ( .A(n236), .ZN(hwdata_o[10]) );
  AOI22_X2 U2106 ( .A1(n3177), .A2(n16786), .B1(n4401), .B2(n3145), .ZN(n236)
         );
  INV_X4 U2107 ( .A(n242), .ZN(hwdata_o[13]) );
  AOI22_X2 U2128 ( .A1(n2556), .A2(n16786), .B1(n4401), .B2(n2259), .ZN(n242)
         );
  INV_X4 U2137 ( .A(n232), .ZN(hwdata_o[8]) );
  AOI22_X2 U2139 ( .A1(n1354), .A2(n16786), .B1(n4401), .B2(n2261), .ZN(n232)
         );
  OAI211_X2 U2140 ( .C1(n3215), .C2(n3217), .A(n3284), .B(n3285), .ZN(n2008)
         );
  NAND2_X2 U2142 ( .A1(n1777), .A2(n3867), .ZN(n3217) );
  NOR4_X4 U2144 ( .A1(n1669), .A2(n1670), .A3(n1613), .A4(n1612), .ZN(
        haddr_o[0]) );
  NAND4_X2 U2165 ( .A1(n1876), .A2(n2674), .A3(n2685), .A4(n2686), .ZN(
        hprot_o[0]) );
  INV_X4 U2174 ( .A(n215), .ZN(hwdata_o[2]) );
  NAND2_X2 U2176 ( .A1(n3177), .A2(n1063), .ZN(n215) );
  INV_X4 U2177 ( .A(n247), .ZN(hwdata_o[15]) );
  INV_X4 U2179 ( .A(n245), .ZN(hwdata_o[14]) );
  OR4_X4 U2181 ( .A1(n948), .A2(n963), .A3(haddr_o[7]), .A4(haddr_o[9]), .ZN(
        n969) );
  INV_X4 U2203 ( .A(n1147), .ZN(haddr_o[7]) );
  INV_X4 U2219 ( .A(n238), .ZN(hwdata_o[11]) );
  AOI22_X2 U2240 ( .A1(n2257), .A2(n16786), .B1(n4401), .B2(n2246), .ZN(n238)
         );
  INV_X4 U2274 ( .A(n234), .ZN(hwdata_o[9]) );
  AOI22_X2 U2309 ( .A1(n4401), .A2(n3287), .B1(n2028), .B2(n16786), .ZN(n234)
         );
  INV_X4 U2331 ( .A(n19), .ZN(hwdata_o[22]) );
  OAI22_X2 U2332 ( .A1(n4203), .A2(n2250), .B1(n4202), .B2(n2251), .ZN(n19) );
  NOR3_X4 U2333 ( .A1(n1088), .A2(n16823), .A3(n1784), .ZN(txev_o) );
  AOI211_X2 U2341 ( .C1(n2376), .C2(n3213), .A(n3609), .B(n3425), .ZN(n2076)
         );
  INV_X4 U2344 ( .A(n3209), .ZN(n3425) );
  OAI21_X4 U2345 ( .B1(n1618), .B2(n979), .A(n1871), .ZN(haddr_o[31]) );
  OAI21_X4 U2346 ( .B1(n1625), .B2(n1622), .A(n1626), .ZN(haddr_o[8]) );
  INV_X4 U2347 ( .A(n16738), .ZN(n16792) );
  INV_X4 U2355 ( .A(n16738), .ZN(n16793) );
  INV_X4 U2379 ( .A(n17104), .ZN(n17103) );
  INV_X4 U2385 ( .A(n17076), .ZN(n17074) );
  INV_X4 U2386 ( .A(n17076), .ZN(n17073) );
  INV_X4 U2402 ( .A(n17056), .ZN(n17053) );
  INV_X4 U2414 ( .A(n17056), .ZN(n17054) );
  INV_X4 U2443 ( .A(n17021), .ZN(n17018) );
  INV_X4 U2452 ( .A(n17021), .ZN(n17019) );
  INV_X4 U2454 ( .A(n17051), .ZN(n17048) );
  INV_X4 U2455 ( .A(n17051), .ZN(n17049) );
  INV_X4 U2457 ( .A(n17071), .ZN(n17068) );
  INV_X4 U2481 ( .A(n17071), .ZN(n17069) );
  INV_X4 U2486 ( .A(n17041), .ZN(n17038) );
  INV_X4 U2491 ( .A(n17041), .ZN(n17039) );
  INV_X4 U2493 ( .A(n17026), .ZN(n17023) );
  INV_X4 U2494 ( .A(n17026), .ZN(n17024) );
  INV_X4 U2496 ( .A(n17076), .ZN(n17075) );
  INV_X4 U2498 ( .A(n17056), .ZN(n17055) );
  INV_X4 U2518 ( .A(n17021), .ZN(n17020) );
  INV_X4 U2530 ( .A(n17051), .ZN(n17050) );
  INV_X4 U2532 ( .A(n17071), .ZN(n17070) );
  INV_X4 U2533 ( .A(n17041), .ZN(n17040) );
  INV_X4 U2535 ( .A(n17026), .ZN(n17025) );
  INV_X4 U2537 ( .A(n16644), .ZN(n17116) );
  INV_X4 U2556 ( .A(n36), .ZN(n17117) );
  INV_X4 U2566 ( .A(n36), .ZN(n17118) );
  INV_X4 U2568 ( .A(n36), .ZN(n17119) );
  INV_X4 U2569 ( .A(n532), .ZN(n597) );
  INV_X4 U2571 ( .A(n16957), .ZN(n16956) );
  INV_X4 U2573 ( .A(n4427), .ZN(n16880) );
  INV_X4 U2593 ( .A(n16788), .ZN(n2337) );
  INV_X4 U2605 ( .A(n1632), .ZN(n17088) );
  INV_X4 U2607 ( .A(n979), .ZN(n17090) );
  INV_X4 U2608 ( .A(n1632), .ZN(n17086) );
  INV_X4 U2610 ( .A(n1632), .ZN(n17087) );
  INV_X4 U2612 ( .A(n979), .ZN(n17091) );
  INV_X4 U2631 ( .A(n979), .ZN(n17089) );
  AND2_X2 U2641 ( .A1(n17102), .A2(n527), .ZN(n16738) );
  INV_X4 U2643 ( .A(n866), .ZN(n17102) );
  INV_X4 U2644 ( .A(n318), .ZN(n17104) );
  NAND2_X2 U2646 ( .A1(n195), .A2(n17096), .ZN(n699) );
  INV_X4 U2648 ( .A(n16742), .ZN(n17077) );
  INV_X4 U2668 ( .A(n16740), .ZN(n17057) );
  INV_X4 U2682 ( .A(n16741), .ZN(n17022) );
  INV_X4 U2684 ( .A(n16743), .ZN(n17052) );
  INV_X4 U2685 ( .A(n16744), .ZN(n17027) );
  INV_X4 U2687 ( .A(n16745), .ZN(n17042) );
  INV_X4 U2689 ( .A(n16740), .ZN(n17056) );
  INV_X4 U2709 ( .A(n16741), .ZN(n17021) );
  INV_X4 U2715 ( .A(n16739), .ZN(n17071) );
  INV_X4 U2719 ( .A(n16742), .ZN(n17076) );
  INV_X4 U2731 ( .A(n16743), .ZN(n17051) );
  INV_X4 U2751 ( .A(n16744), .ZN(n17026) );
  INV_X4 U2755 ( .A(n16745), .ZN(n17041) );
  INV_X4 U2763 ( .A(n200), .ZN(n17092) );
  INV_X4 U2765 ( .A(n200), .ZN(n17093) );
  INV_X4 U2766 ( .A(n866), .ZN(n17100) );
  INV_X4 U2768 ( .A(n866), .ZN(n17101) );
  INV_X4 U2790 ( .A(n16644), .ZN(n17115) );
  INV_X4 U2798 ( .A(n17046), .ZN(n17043) );
  INV_X4 U2803 ( .A(n17046), .ZN(n17044) );
  INV_X4 U2821 ( .A(n17031), .ZN(n17028) );
  INV_X4 U2827 ( .A(n17031), .ZN(n17029) );
  INV_X4 U2828 ( .A(n16644), .ZN(n17114) );
  INV_X4 U2830 ( .A(n17046), .ZN(n17045) );
  INV_X4 U2832 ( .A(n17031), .ZN(n17030) );
  INV_X4 U2833 ( .A(n54), .ZN(n29) );
  INV_X4 U2855 ( .A(n16739), .ZN(n17072) );
  INV_X4 U2859 ( .A(n17113), .ZN(n17112) );
  INV_X4 U2865 ( .A(n17113), .ZN(n17111) );
  INV_X4 U2867 ( .A(n17061), .ZN(n17058) );
  INV_X4 U2868 ( .A(n17061), .ZN(n17059) );
  INV_X4 U2870 ( .A(n17081), .ZN(n17078) );
  INV_X4 U2872 ( .A(n17081), .ZN(n17079) );
  INV_X4 U2880 ( .A(n17066), .ZN(n17063) );
  INV_X4 U2882 ( .A(n17066), .ZN(n17064) );
  INV_X4 U2910 ( .A(n17016), .ZN(n17013) );
  INV_X4 U2927 ( .A(n17016), .ZN(n17014) );
  INV_X4 U2936 ( .A(n17036), .ZN(n17033) );
  INV_X4 U2941 ( .A(n17036), .ZN(n17034) );
  INV_X4 U2956 ( .A(n17061), .ZN(n17060) );
  INV_X4 U2964 ( .A(n17081), .ZN(n17080) );
  INV_X4 U2966 ( .A(n17066), .ZN(n17065) );
  INV_X4 U2967 ( .A(n17036), .ZN(n17035) );
  INV_X4 U2969 ( .A(n17016), .ZN(n17015) );
  NAND2_X2 U2971 ( .A1(n473), .A2(n466), .ZN(n443) );
  NAND2_X2 U2991 ( .A1(n16870), .A2(n16849), .ZN(n532) );
  NAND2_X2 U3000 ( .A1(n16825), .A2(n16860), .ZN(n653) );
  INV_X4 U3002 ( .A(n585), .ZN(n991) );
  INV_X4 U3003 ( .A(n2222), .ZN(n16957) );
  INV_X4 U3005 ( .A(n2637), .ZN(n16979) );
  INV_X4 U3007 ( .A(n2184), .ZN(n16971) );
  INV_X4 U3034 ( .A(n640), .ZN(n527) );
  INV_X4 U3037 ( .A(n17097), .ZN(n17096) );
  INV_X4 U3071 ( .A(n3180), .ZN(n16988) );
  INV_X4 U3078 ( .A(n2184), .ZN(n16970) );
  INV_X4 U3086 ( .A(n2637), .ZN(n16981) );
  NAND2_X2 U3088 ( .A1(n16825), .A2(n16805), .ZN(n696) );
  NAND2_X2 U3094 ( .A1(n16859), .A2(n17096), .ZN(n745) );
  INV_X4 U3098 ( .A(n715), .ZN(n526) );
  INV_X4 U3112 ( .A(n1086), .ZN(n1574) );
  INV_X4 U3127 ( .A(n673), .ZN(n827) );
  INV_X4 U3130 ( .A(n1519), .ZN(n529) );
  INV_X4 U3141 ( .A(n918), .ZN(n565) );
  INV_X4 U3148 ( .A(n1514), .ZN(n17083) );
  INV_X4 U3157 ( .A(n1514), .ZN(n17084) );
  INV_X4 U3159 ( .A(n2184), .ZN(n16972) );
  INV_X4 U3160 ( .A(n16957), .ZN(n16955) );
  INV_X4 U3162 ( .A(n16991), .ZN(n16990) );
  INV_X4 U3164 ( .A(n16652), .ZN(n16895) );
  NOR2_X2 U3175 ( .A1(n1754), .A2(n2233), .ZN(n2391) );
  INV_X4 U3188 ( .A(n16957), .ZN(n16954) );
  INV_X4 U3220 ( .A(n2637), .ZN(n16980) );
  INV_X4 U3224 ( .A(n16648), .ZN(n16882) );
  INV_X4 U3225 ( .A(n1514), .ZN(n17085) );
  INV_X4 U3241 ( .A(n16911), .ZN(n16910) );
  INV_X4 U3244 ( .A(n16652), .ZN(n16894) );
  INV_X4 U3248 ( .A(n16649), .ZN(n16875) );
  INV_X4 U3262 ( .A(n16648), .ZN(n16881) );
  INV_X4 U3264 ( .A(n16650), .ZN(n16873) );
  INV_X4 U3265 ( .A(n16650), .ZN(n16874) );
  INV_X4 U3267 ( .A(n17099), .ZN(n17098) );
  INV_X4 U3269 ( .A(n16911), .ZN(n16909) );
  INV_X4 U3275 ( .A(n851), .ZN(n592) );
  INV_X4 U3296 ( .A(n16652), .ZN(n16896) );
  INV_X4 U3327 ( .A(n16649), .ZN(n16876) );
  INV_X4 U3338 ( .A(n16684), .ZN(n16788) );
  INV_X4 U3342 ( .A(n2127), .ZN(n16992) );
  INV_X4 U3348 ( .A(n16684), .ZN(n16789) );
  INV_X4 U3350 ( .A(n3279), .ZN(n16942) );
  INV_X4 U3351 ( .A(n3118), .ZN(n16951) );
  INV_X4 U3353 ( .A(n3118), .ZN(n16953) );
  INV_X4 U3355 ( .A(n3275), .ZN(n16948) );
  INV_X4 U3356 ( .A(n3277), .ZN(n16945) );
  INV_X4 U3366 ( .A(n3277), .ZN(n16947) );
  INV_X4 U3383 ( .A(n3275), .ZN(n16950) );
  INV_X4 U3384 ( .A(n1622), .ZN(n1628) );
  INV_X4 U3386 ( .A(n2127), .ZN(n16993) );
  INV_X4 U3387 ( .A(n3279), .ZN(n16943) );
  INV_X4 U3389 ( .A(n3118), .ZN(n16952) );
  INV_X4 U3390 ( .A(n3275), .ZN(n16949) );
  INV_X4 U3392 ( .A(n3277), .ZN(n16946) );
  INV_X4 U3393 ( .A(n3279), .ZN(n16944) );
  NAND2_X2 U3396 ( .A1(n897), .A2(n16870), .ZN(n650) );
  INV_X4 U3397 ( .A(n499), .ZN(n195) );
  INV_X4 U3399 ( .A(n2243), .ZN(n17008) );
  INV_X4 U3400 ( .A(n2243), .ZN(n17007) );
  INV_X4 U3402 ( .A(n2243), .ZN(n17006) );
  INV_X4 U3403 ( .A(n2501), .ZN(n16994) );
  INV_X4 U3405 ( .A(n2501), .ZN(n16995) );
  AND2_X2 U3406 ( .A1(n3438), .A2(n3446), .ZN(n16739) );
  INV_X4 U3409 ( .A(n42), .ZN(n17113) );
  AND2_X2 U3410 ( .A1(n3445), .A2(n3435), .ZN(n16740) );
  AND2_X2 U3412 ( .A1(n3442), .A2(n3435), .ZN(n16741) );
  AND2_X2 U3413 ( .A1(n3435), .A2(n3446), .ZN(n16742) );
  AND2_X2 U3415 ( .A1(n3445), .A2(n3438), .ZN(n16743) );
  AND2_X2 U3416 ( .A1(n3442), .A2(n3438), .ZN(n16744) );
  AND2_X2 U3418 ( .A1(n3437), .A2(n3438), .ZN(n16745) );
  INV_X4 U3419 ( .A(n3213), .ZN(n3215) );
  INV_X4 U3423 ( .A(n16750), .ZN(n17017) );
  INV_X4 U3424 ( .A(n16748), .ZN(n17037) );
  INV_X4 U3427 ( .A(n16749), .ZN(n17062) );
  INV_X4 U3428 ( .A(n16751), .ZN(n17082) );
  INV_X4 U3431 ( .A(n16748), .ZN(n17036) );
  INV_X4 U3432 ( .A(n16749), .ZN(n17061) );
  INV_X4 U3436 ( .A(n16750), .ZN(n17016) );
  INV_X4 U3445 ( .A(n16751), .ZN(n17081) );
  INV_X4 U3447 ( .A(n16746), .ZN(n17046) );
  INV_X4 U3448 ( .A(n16747), .ZN(n17031) );
  INV_X4 U3450 ( .A(n17004), .ZN(n17001) );
  INV_X4 U3452 ( .A(n17004), .ZN(n17002) );
  INV_X4 U3453 ( .A(n17004), .ZN(n17003) );
  INV_X4 U3454 ( .A(n16752), .ZN(n17067) );
  INV_X4 U3459 ( .A(n16746), .ZN(n17047) );
  INV_X4 U3475 ( .A(n16747), .ZN(n17032) );
  INV_X4 U3476 ( .A(n16752), .ZN(n17066) );
  NAND2_X2 U3494 ( .A1(n16834), .A2(n16864), .ZN(n585) );
  INV_X4 U3562 ( .A(n2182), .ZN(n16964) );
  INV_X4 U3566 ( .A(n16754), .ZN(n16984) );
  INV_X4 U3568 ( .A(n2191), .ZN(n16963) );
  INV_X4 U3574 ( .A(n2182), .ZN(n16966) );
  INV_X4 U3577 ( .A(n16753), .ZN(n16969) );
  INV_X4 U3580 ( .A(n2190), .ZN(n16960) );
  INV_X4 U3581 ( .A(n16865), .ZN(n16864) );
  INV_X4 U3583 ( .A(n16839), .ZN(n16837) );
  INV_X4 U3637 ( .A(n16826), .ZN(n16825) );
  INV_X4 U3641 ( .A(n16861), .ZN(n16860) );
  INV_X4 U3642 ( .A(n16871), .ZN(n16870) );
  INV_X4 U3645 ( .A(n16850), .ZN(n16849) );
  INV_X4 U3646 ( .A(n797), .ZN(n17097) );
  NAND2_X2 U3649 ( .A1(n16851), .A2(n16856), .ZN(n715) );
  NAND2_X2 U3650 ( .A1(n16848), .A2(n16839), .ZN(n1086) );
  NAND2_X2 U3651 ( .A1(n16834), .A2(n17096), .ZN(n640) );
  NAND2_X2 U3652 ( .A1(n16845), .A2(n16860), .ZN(n617) );
  NAND2_X2 U3655 ( .A1(n16856), .A2(n16842), .ZN(n1104) );
  INV_X4 U3656 ( .A(n16755), .ZN(n16976) );
  INV_X4 U3658 ( .A(n16755), .ZN(n16978) );
  INV_X4 U3659 ( .A(n16759), .ZN(n16939) );
  INV_X4 U3660 ( .A(n16760), .ZN(n16916) );
  INV_X4 U3663 ( .A(n16756), .ZN(n16933) );
  INV_X4 U3665 ( .A(n16754), .ZN(n16982) );
  INV_X4 U3666 ( .A(n16763), .ZN(n16877) );
  INV_X4 U3669 ( .A(n16753), .ZN(n16967) );
  INV_X4 U3671 ( .A(n16753), .ZN(n16968) );
  INV_X4 U3673 ( .A(n2190), .ZN(n16958) );
  INV_X4 U3674 ( .A(n2190), .ZN(n16959) );
  INV_X4 U3675 ( .A(n16762), .ZN(n16913) );
  INV_X4 U3695 ( .A(n2191), .ZN(n16962) );
  INV_X4 U3696 ( .A(n2182), .ZN(n16965) );
  INV_X4 U3705 ( .A(n16757), .ZN(n16905) );
  INV_X4 U3721 ( .A(n16761), .ZN(n16908) );
  INV_X4 U3729 ( .A(n16758), .ZN(n16885) );
  INV_X4 U3732 ( .A(n16850), .ZN(n16848) );
  INV_X4 U3733 ( .A(n16844), .ZN(n16842) );
  INV_X4 U3737 ( .A(n16833), .ZN(n16828) );
  INV_X4 U3740 ( .A(n16832), .ZN(n16830) );
  INV_X4 U3741 ( .A(n16728), .ZN(n16836) );
  INV_X4 U3746 ( .A(n16832), .ZN(n16831) );
  INV_X4 U3749 ( .A(n16844), .ZN(n16843) );
  NAND2_X2 U3750 ( .A1(n16866), .A2(n16855), .ZN(n1519) );
  NAND2_X2 U3755 ( .A1(n16838), .A2(n16862), .ZN(n673) );
  NAND2_X2 U3758 ( .A1(n16855), .A2(n16839), .ZN(n918) );
  INV_X4 U3759 ( .A(n2543), .ZN(n2198) );
  INV_X4 U3765 ( .A(n4211), .ZN(n16911) );
  INV_X1 U3768 ( .A(n16755), .ZN(n16977) );
  INV_X4 U3769 ( .A(n2169), .ZN(n16991) );
  INV_X4 U3773 ( .A(n16759), .ZN(n16940) );
  INV_X4 U3776 ( .A(n16756), .ZN(n16934) );
  INV_X4 U3777 ( .A(n16767), .ZN(n16886) );
  INV_X4 U3782 ( .A(n16764), .ZN(n16897) );
  INV_X4 U3785 ( .A(n2191), .ZN(n16961) );
  INV_X4 U3786 ( .A(n16766), .ZN(n16891) );
  INV_X4 U3791 ( .A(n16765), .ZN(n16902) );
  INV_X4 U3794 ( .A(n16861), .ZN(n16859) );
  INV_X4 U3795 ( .A(n16861), .ZN(n16858) );
  INV_X4 U3825 ( .A(n16690), .ZN(n16824) );
  INV_X4 U3842 ( .A(n16694), .ZN(n16854) );
  INV_X4 U3865 ( .A(n16850), .ZN(n16847) );
  INV_X4 U3873 ( .A(n16694), .ZN(n16853) );
  INV_X4 U3874 ( .A(n16690), .ZN(n16823) );
  INV_X4 U3904 ( .A(n16844), .ZN(n16841) );
  INV_X4 U3937 ( .A(n16689), .ZN(n16868) );
  INV_X4 U3938 ( .A(n16694), .ZN(n16855) );
  INV_X4 U3940 ( .A(n16728), .ZN(n16838) );
  NOR2_X2 U3943 ( .A1(n2077), .A2(n2078), .ZN(n1808) );
  NAND2_X2 U3945 ( .A1(n16851), .A2(n16862), .ZN(n499) );
  INV_X4 U3946 ( .A(n16760), .ZN(n16915) );
  INV_X4 U3948 ( .A(n16754), .ZN(n16983) );
  INV_X4 U3950 ( .A(n16762), .ZN(n16912) );
  INV_X4 U3953 ( .A(n16760), .ZN(n16917) );
  INV_X4 U3963 ( .A(n16762), .ZN(n16914) );
  INV_X4 U3966 ( .A(n16757), .ZN(n16904) );
  INV_X4 U3967 ( .A(n16761), .ZN(n16907) );
  INV_X4 U3968 ( .A(n16759), .ZN(n16941) );
  INV_X4 U3975 ( .A(n16756), .ZN(n16935) );
  INV_X4 U3976 ( .A(n16651), .ZN(n16893) );
  INV_X4 U3981 ( .A(n16765), .ZN(n16901) );
  INV_X4 U3982 ( .A(n16766), .ZN(n16890) );
  INV_X4 U3984 ( .A(n16758), .ZN(n16884) );
  INV_X4 U3996 ( .A(n16767), .ZN(n16887) );
  INV_X4 U3997 ( .A(n16763), .ZN(n16878) );
  INV_X4 U3998 ( .A(n16764), .ZN(n16898) );
  INV_X4 U4000 ( .A(n16651), .ZN(n16892) );
  INV_X4 U4010 ( .A(n16686), .ZN(n17099) );
  INV_X4 U4013 ( .A(n16767), .ZN(n16888) );
  INV_X4 U4014 ( .A(n16763), .ZN(n16879) );
  INV_X4 U4018 ( .A(n16764), .ZN(n16899) );
  INV_X4 U4021 ( .A(n16790), .ZN(n16791) );
  INV_X4 U4022 ( .A(n2519), .ZN(n16790) );
  AOI211_X2 U4027 ( .C1(n2250), .C2(n17008), .A(n2520), .B(n2521), .ZN(n2519)
         );
  INV_X4 U4028 ( .A(n16757), .ZN(n16903) );
  INV_X4 U4031 ( .A(n16761), .ZN(n16906) );
  INV_X4 U4032 ( .A(n16765), .ZN(n16900) );
  INV_X4 U4037 ( .A(n16766), .ZN(n16889) );
  INV_X4 U4040 ( .A(n16758), .ZN(n16883) );
  NAND2_X2 U4041 ( .A1(n16806), .A2(n16820), .ZN(n851) );
  INV_X4 U4047 ( .A(n16681), .ZN(n16820) );
  INV_X4 U4050 ( .A(n16681), .ZN(n16819) );
  INV_X4 U4051 ( .A(n16689), .ZN(n16869) );
  NAND2_X2 U4055 ( .A1(n400), .A2(n1340), .ZN(n379) );
  INV_X4 U4058 ( .A(n16832), .ZN(n16829) );
  INV_X4 U4059 ( .A(n16813), .ZN(n16812) );
  INV_X4 U4064 ( .A(n2126), .ZN(n2131) );
  INV_X4 U4067 ( .A(n2926), .ZN(n2882) );
  INV_X4 U4068 ( .A(n2124), .ZN(n2055) );
  INV_X4 U4073 ( .A(n2981), .ZN(n2878) );
  INV_X4 U4076 ( .A(n4202), .ZN(n4203) );
  INV_X4 U4077 ( .A(n2998), .ZN(n2922) );
  AND2_X2 U4087 ( .A1(n3445), .A2(n3443), .ZN(n16746) );
  AND2_X2 U4090 ( .A1(n3442), .A2(n3443), .ZN(n16747) );
  OAI21_X2 U4091 ( .B1(n17096), .B2(n4070), .A(n3546), .ZN(n3213) );
  NOR2_X2 U4094 ( .A1(n17126), .A2(n1007), .ZN(n37) );
  NAND4_X2 U4114 ( .A1(n809), .A2(n760), .A3(n16819), .A4(n16856), .ZN(n200)
         );
  NAND2_X2 U4115 ( .A1(n791), .A2(n16725), .ZN(n819) );
  AND2_X2 U4118 ( .A1(n3437), .A2(n3439), .ZN(n16748) );
  AND2_X2 U4119 ( .A1(n3445), .A2(n3439), .ZN(n16749) );
  AND2_X2 U4123 ( .A1(n3442), .A2(n3439), .ZN(n16750) );
  AND2_X2 U4124 ( .A1(n3446), .A2(n3439), .ZN(n16751) );
  INV_X4 U4127 ( .A(n16768), .ZN(n17005) );
  INV_X4 U4128 ( .A(n16768), .ZN(n17004) );
  INV_X4 U4133 ( .A(n16999), .ZN(n16996) );
  INV_X4 U4134 ( .A(n16999), .ZN(n16997) );
  INV_X4 U4137 ( .A(n16687), .ZN(n16816) );
  INV_X4 U4138 ( .A(n16999), .ZN(n16998) );
  AND2_X2 U4143 ( .A1(n3443), .A2(n3446), .ZN(n16752) );
  NOR2_X2 U4144 ( .A1(n1125), .A2(n1124), .ZN(n1317) );
  INV_X4 U4147 ( .A(n16769), .ZN(n17109) );
  INV_X4 U4148 ( .A(n16769), .ZN(n17110) );
  INV_X4 U4154 ( .A(n17127), .ZN(n17124) );
  INV_X4 U4155 ( .A(n17095), .ZN(n17094) );
  INV_X4 U4158 ( .A(n16687), .ZN(n16815) );
  INV_X4 U4159 ( .A(n17126), .ZN(n17122) );
  INV_X4 U4163 ( .A(n17126), .ZN(n17123) );
  INV_X4 U4164 ( .A(n16647), .ZN(n17106) );
  INV_X4 U4167 ( .A(n16647), .ZN(n17105) );
  INV_X4 U4168 ( .A(n17126), .ZN(n17125) );
  NAND2_X2 U4174 ( .A1(n373), .A2(n1109), .ZN(n1131) );
  NAND3_X2 U4175 ( .A1(n3592), .A2(n3436), .A3(n3593), .ZN(n16753) );
  NAND2_X2 U4178 ( .A1(n3593), .A2(n3480), .ZN(n16754) );
  INV_X4 U4179 ( .A(n16770), .ZN(n16985) );
  INV_X4 U4194 ( .A(n16840), .ZN(n16839) );
  INV_X4 U4197 ( .A(n16827), .ZN(n16826) );
  OR2_X1 U4198 ( .A1(n16956), .A2(n3601), .ZN(n16755) );
  AND2_X2 U4204 ( .A1(n4162), .A2(n3492), .ZN(n16756) );
  AND2_X2 U4210 ( .A1(n4657), .A2(n4658), .ZN(n16757) );
  AND2_X2 U4224 ( .A1(n4662), .A2(n4657), .ZN(n16758) );
  NAND2_X2 U4226 ( .A1(n4163), .A2(n3480), .ZN(n16759) );
  NAND2_X2 U4230 ( .A1(n4663), .A2(n4659), .ZN(n16760) );
  AND2_X2 U4231 ( .A1(n4659), .A2(n4658), .ZN(n16761) );
  NAND2_X2 U4236 ( .A1(n4662), .A2(n4659), .ZN(n16762) );
  NAND2_X2 U4241 ( .A1(n4661), .A2(n4657), .ZN(n16763) );
  INV_X4 U4243 ( .A(n16852), .ZN(n16851) );
  INV_X4 U4249 ( .A(n16835), .ZN(n16833) );
  INV_X4 U4250 ( .A(n16835), .ZN(n16832) );
  INV_X4 U4260 ( .A(n16857), .ZN(n16856) );
  INV_X2 U4263 ( .A(n16770), .ZN(n16986) );
  INV_X1 U4264 ( .A(n16770), .ZN(n16987) );
  INV_X4 U4268 ( .A(n16846), .ZN(n16845) );
  INV_X4 U4271 ( .A(n16872), .ZN(n16871) );
  INV_X4 U4272 ( .A(n16822), .ZN(n16821) );
  INV_X4 U4277 ( .A(n16773), .ZN(n16973) );
  INV_X4 U4280 ( .A(n16772), .ZN(n16930) );
  INV_X4 U4281 ( .A(n16771), .ZN(n16918) );
  INV_X4 U4286 ( .A(n16775), .ZN(n16936) );
  INV_X4 U4289 ( .A(n16774), .ZN(n16927) );
  INV_X4 U4290 ( .A(n16773), .ZN(n16975) );
  NAND2_X2 U4291 ( .A1(n4665), .A2(n4658), .ZN(n16764) );
  NAND3_X2 U4297 ( .A1(n4662), .A2(n3436), .A3(n4660), .ZN(n16765) );
  NAND2_X2 U4300 ( .A1(n4665), .A2(n4662), .ZN(n16766) );
  NAND2_X2 U4301 ( .A1(n4660), .A2(n4663), .ZN(n16767) );
  INV_X4 U4302 ( .A(n16863), .ZN(n16862) );
  INV_X4 U4307 ( .A(n16777), .ZN(n16924) );
  INV_X2 U4310 ( .A(n16777), .ZN(n16925) );
  INV_X4 U4311 ( .A(n16776), .ZN(n16921) );
  INV_X2 U4312 ( .A(n16776), .ZN(n16922) );
  INV_X4 U4314 ( .A(n16867), .ZN(n16866) );
  INV_X4 U4315 ( .A(n16772), .ZN(n16931) );
  INV_X4 U4320 ( .A(n16771), .ZN(n16919) );
  INV_X4 U4323 ( .A(n16775), .ZN(n16937) );
  INV_X4 U4324 ( .A(n16774), .ZN(n16928) );
  INV_X4 U4325 ( .A(n16773), .ZN(n16974) );
  INV_X4 U4326 ( .A(n16772), .ZN(n16932) );
  INV_X4 U4335 ( .A(n16771), .ZN(n16920) );
  INV_X4 U4336 ( .A(n16775), .ZN(n16938) );
  INV_X4 U4338 ( .A(n16774), .ZN(n16929) );
  INV_X1 U4339 ( .A(n16777), .ZN(n16926) );
  INV_X1 U4340 ( .A(n16776), .ZN(n16923) );
  NOR2_X2 U4343 ( .A1(n179), .A2(n2001), .ZN(n1750) );
  INV_X4 U4344 ( .A(n16818), .ZN(n16817) );
  NOR2_X2 U4345 ( .A1(n503), .A2(n16659), .ZN(n475) );
  NAND2_X2 U4347 ( .A1(n16680), .A2(n16820), .ZN(n616) );
  INV_X4 U4348 ( .A(n16802), .ZN(n16804) );
  INV_X4 U4350 ( .A(n16814), .ZN(n16813) );
  NAND2_X2 U4351 ( .A1(n2231), .A2(n2172), .ZN(n1900) );
  INV_X4 U4352 ( .A(n17012), .ZN(n17009) );
  INV_X4 U4353 ( .A(n17012), .ZN(n17010) );
  INV_X4 U4354 ( .A(n17012), .ZN(n17011) );
  NAND2_X2 U4355 ( .A1(n252), .A2(n2882), .ZN(n2948) );
  NAND2_X2 U4362 ( .A1(n3873), .A2(n2882), .ZN(n3011) );
  INV_X4 U4365 ( .A(n2918), .ZN(n2879) );
  NAND2_X2 U4366 ( .A1(n336), .A2(n1002), .ZN(n334) );
  NAND2_X2 U4367 ( .A1(n1759), .A2(n4077), .ZN(n2998) );
  NAND2_X2 U4369 ( .A1(n1063), .A2(n1612), .ZN(n4202) );
  NAND2_X2 U4370 ( .A1(n2250), .A2(n1063), .ZN(n226) );
  NAND2_X2 U4374 ( .A1(n2196), .A2(n1063), .ZN(n229) );
  INV_X4 U4379 ( .A(n16779), .ZN(n17120) );
  INV_X4 U4381 ( .A(n16779), .ZN(n17121) );
  INV_X4 U4395 ( .A(n1385), .ZN(n1124) );
  NAND2_X2 U4402 ( .A1(n822), .A2(n16807), .ZN(n478) );
  AND3_X2 U4404 ( .A1(n3435), .A2(n3436), .A3(n3437), .ZN(n16768) );
  INV_X4 U4406 ( .A(n16780), .ZN(n17000) );
  INV_X4 U4417 ( .A(n16780), .ZN(n16999) );
  NAND2_X2 U4418 ( .A1(n1893), .A2(n253), .ZN(n1892) );
  NAND2_X2 U4419 ( .A1(n1897), .A2(n253), .ZN(n1895) );
  AND3_X2 U4424 ( .A1(n17107), .A2(n315), .A3(n314), .ZN(n16769) );
  INV_X4 U4425 ( .A(n16781), .ZN(n17095) );
  INV_X4 U4435 ( .A(hready_i), .ZN(n17126) );
  INV_X4 U4436 ( .A(n16798), .ZN(n16799) );
  NAND2_X2 U4440 ( .A1(n252), .A2(n253), .ZN(n213) );
  NAND2_X2 U4441 ( .A1(n1890), .A2(n253), .ZN(n1889) );
  NAND2_X2 U4444 ( .A1(n1887), .A2(n253), .ZN(n1886) );
  INV_X4 U4445 ( .A(n17108), .ZN(n17107) );
  INV_X4 U4448 ( .A(hready_i), .ZN(n17127) );
  BUF_X4 U4449 ( .A(n17188), .Z(n17130) );
  BUF_X4 U4452 ( .A(n17187), .Z(n17132) );
  BUF_X4 U4453 ( .A(n17195), .Z(n17129) );
  BUF_X4 U4454 ( .A(n17194), .Z(n17137) );
  BUF_X4 U4455 ( .A(n17194), .Z(n17136) );
  BUF_X4 U4459 ( .A(n17194), .Z(n17138) );
  BUF_X4 U4460 ( .A(n17186), .Z(n17134) );
  BUF_X4 U4463 ( .A(n17193), .Z(n17133) );
  BUF_X4 U4464 ( .A(n17192), .Z(n17135) );
  BUF_X4 U4467 ( .A(n17194), .Z(n17131) );
  BUF_X4 U4468 ( .A(n17195), .Z(n17128) );
  BUF_X4 U4471 ( .A(n17190), .Z(n17159) );
  BUF_X4 U4472 ( .A(n17194), .Z(n17140) );
  BUF_X4 U4473 ( .A(n17191), .Z(n17154) );
  BUF_X4 U4474 ( .A(n17192), .Z(n17151) );
  BUF_X4 U4478 ( .A(n17193), .Z(n17142) );
  BUF_X4 U4480 ( .A(n17194), .Z(n17141) );
  BUF_X4 U4481 ( .A(n17190), .Z(n17158) );
  BUF_X4 U4486 ( .A(n17188), .Z(n17172) );
  BUF_X4 U4487 ( .A(n17188), .Z(n17171) );
  BUF_X4 U4490 ( .A(n17188), .Z(n17170) );
  BUF_X4 U4491 ( .A(n17188), .Z(n17169) );
  BUF_X4 U4494 ( .A(n17189), .Z(n17168) );
  BUF_X4 U4495 ( .A(n17189), .Z(n17166) );
  BUF_X4 U4498 ( .A(n17189), .Z(n17165) );
  BUF_X4 U4499 ( .A(n17189), .Z(n17164) );
  BUF_X4 U4500 ( .A(n17189), .Z(n17163) );
  BUF_X4 U4504 ( .A(n17190), .Z(n17162) );
  BUF_X4 U4505 ( .A(n17190), .Z(n17161) );
  BUF_X4 U4508 ( .A(n17189), .Z(n17167) );
  BUF_X4 U4509 ( .A(n17186), .Z(n17185) );
  BUF_X4 U4512 ( .A(n17186), .Z(n17184) );
  BUF_X4 U4513 ( .A(n17186), .Z(n17183) );
  BUF_X4 U4516 ( .A(n17186), .Z(n17182) );
  BUF_X4 U4517 ( .A(n17186), .Z(n17181) );
  BUF_X4 U4519 ( .A(n17187), .Z(n17179) );
  BUF_X4 U4523 ( .A(n17187), .Z(n17178) );
  BUF_X4 U4527 ( .A(n17187), .Z(n17177) );
  BUF_X4 U4528 ( .A(n17187), .Z(n17176) );
  BUF_X4 U4531 ( .A(n17187), .Z(n17175) );
  BUF_X4 U4532 ( .A(n17188), .Z(n17174) );
  BUF_X4 U4535 ( .A(n17188), .Z(n17173) );
  BUF_X4 U4536 ( .A(n17187), .Z(n17180) );
  BUF_X4 U4539 ( .A(n17192), .Z(n17150) );
  BUF_X4 U4540 ( .A(n17192), .Z(n17149) );
  BUF_X4 U4543 ( .A(n17192), .Z(n17148) );
  BUF_X4 U4544 ( .A(n17193), .Z(n17147) );
  BUF_X4 U4546 ( .A(n17193), .Z(n17146) );
  BUF_X4 U4548 ( .A(n17193), .Z(n17145) );
  BUF_X4 U4552 ( .A(n17193), .Z(n17143) );
  BUF_X4 U4553 ( .A(n17193), .Z(n17144) );
  BUF_X4 U4556 ( .A(n17190), .Z(n17160) );
  BUF_X4 U4557 ( .A(n17191), .Z(n17157) );
  BUF_X4 U4560 ( .A(n17191), .Z(n17156) );
  BUF_X4 U4561 ( .A(n17191), .Z(n17155) );
  BUF_X4 U4564 ( .A(n17192), .Z(n17153) );
  BUF_X4 U4565 ( .A(n17192), .Z(n17152) );
  BUF_X4 U4566 ( .A(n17194), .Z(n17139) );
  OR4_X1 U4570 ( .A1(n2184), .A2(n5036), .A3(n4978), .A4(n4959), .ZN(n16770)
         );
  NAND3_X2 U4571 ( .A1(n4959), .A2(n3592), .A3(n5252), .ZN(n16771) );
  AND2_X2 U4574 ( .A1(n4162), .A2(n5252), .ZN(n16772) );
  NAND3_X2 U4575 ( .A1(n3592), .A2(n4968), .A3(n3593), .ZN(n16773) );
  NAND3_X2 U4578 ( .A1(n3592), .A2(n3492), .A3(n4959), .ZN(n16774) );
  NAND2_X2 U4579 ( .A1(n4163), .A2(n5036), .ZN(n16775) );
  OR4_X1 U4582 ( .A1(n3488), .A2(n3495), .A3(n5252), .A4(n5036), .ZN(n16776)
         );
  INV_X4 U4583 ( .A(n3180), .ZN(n16989) );
  OR4_X1 U4584 ( .A1(n3488), .A2(n3495), .A3(n3480), .A4(n5252), .ZN(n16777)
         );
  OAI21_X2 U4588 ( .B1(n1341), .B2(n1066), .A(n183), .ZN(n422) );
  INV_X4 U4589 ( .A(n2015), .ZN(n17012) );
  NAND2_X2 U4592 ( .A1(n5027), .A2(n2172), .ZN(n1821) );
  NAND2_X2 U4593 ( .A1(n5027), .A2(n5120), .ZN(n3566) );
  BUF_X4 U4596 ( .A(n4239), .Z(n16786) );
  NAND2_X2 U4597 ( .A1(n5120), .A2(n2231), .ZN(n1820) );
  NAND3_X2 U4600 ( .A1(n2882), .A2(n5149), .A3(n1111), .ZN(n2918) );
  INV_X4 U4601 ( .A(n16685), .ZN(n16787) );
  OR2_X1 U4607 ( .A1(n16778), .A2(n16647), .ZN(n266) );
  XOR2_X2 U4608 ( .A(sub_2068_A_23_), .B(sub_2068_carry_23_), .Z(n16778) );
  NAND2_X2 U4609 ( .A1(n37), .A2(n180), .ZN(n16779) );
  AND3_X2 U4610 ( .A1(n3435), .A2(n4968), .A3(n3437), .ZN(n16780) );
  INV_X4 U4622 ( .A(n265), .ZN(n17108) );
  OR3_X1 U4638 ( .A1(n5007), .A2(n4905), .A3(n261), .ZN(n16781) );
  BUF_X4 U4659 ( .A(hreset_n), .Z(n17189) );
  BUF_X4 U4660 ( .A(hreset_n), .Z(n17188) );
  BUF_X4 U4661 ( .A(hreset_n), .Z(n17187) );
  BUF_X4 U4666 ( .A(hreset_n), .Z(n17186) );
  BUF_X4 U4667 ( .A(hreset_n), .Z(n17193) );
  BUF_X4 U4668 ( .A(hreset_n), .Z(n17190) );
  BUF_X4 U4677 ( .A(hreset_n), .Z(n17192) );
  BUF_X4 U4678 ( .A(hreset_n), .Z(n17191) );
  BUF_X4 U4684 ( .A(hreset_n), .Z(n17194) );
  BUF_X4 U4689 ( .A(hreset_n), .Z(n17195) );
  XNOR2_X2 U4696 ( .A(add_2073_A_7_), .B(n16677), .ZN(n16782) );
  INV_X4 U4697 ( .A(n16782), .ZN(add_2073_SUM_7_) );
  XNOR2_X2 U4698 ( .A(add_2073_A_31_), .B(n16654), .ZN(n16783) );
  INV_X4 U4701 ( .A(n16783), .ZN(add_2073_SUM_31_) );
  NAND2_X2 U4702 ( .A1(add_2073_A_32_), .A2(n16660), .ZN(n16784) );
  XNOR2_X2 U4703 ( .A(add_2082_carry[33]), .B(n16784), .ZN(U4_DATA1_0) );
  XNOR2_X2 U4706 ( .A(add_2073_B_1_), .B(n16675), .ZN(n16785) );
  INV_X4 U4708 ( .A(n16785), .ZN(add_2073_SUM_1_) );
  INV_X4 U4711 ( .A(n1963), .ZN(n731) );
  INV_X4 U4713 ( .A(n1228), .ZN(n708) );
  INV_X4 U4715 ( .A(n945), .ZN(n483) );
  INV_X4 U4720 ( .A(n1882), .ZN(n897) );
  INV_X4 U4721 ( .A(n1198), .ZN(n473) );
  INV_X4 U4725 ( .A(n579), .ZN(n466) );
  NAND3_X2 U4726 ( .A1(n4706), .A2(n4707), .A3(n4708), .ZN(n610) );
  INV_X4 U4727 ( .A(n2719), .ZN(n2732) );
  NAND2_X2 U4728 ( .A1(n4663), .A2(n4657), .ZN(n4427) );
  INV_X4 U4732 ( .A(n4335), .ZN(n4192) );
  INV_X4 U4733 ( .A(n1234), .ZN(n563) );
  INV_X4 U4736 ( .A(n1125), .ZN(n1314) );
  INV_X4 U4774 ( .A(n2723), .ZN(n2074) );
  NAND2_X2 U4778 ( .A1(n3549), .A2(n3550), .ZN(n2126) );
  NAND4_X2 U4779 ( .A1(n3532), .A2(n16866), .A3(n16826), .A4(n1697), .ZN(n2501) );
  INV_X4 U4780 ( .A(n713), .ZN(n543) );
  AND2_X4 U4782 ( .A1(n44), .A2(n2103), .ZN(n3434) );
  AND3_X4 U4783 ( .A1(n48), .A2(n3403), .A3(n3404), .ZN(n3402) );
  AND3_X4 U4796 ( .A1(n144), .A2(n3352), .A3(n3353), .ZN(n3351) );
  INV_X4 U4797 ( .A(n2875), .ZN(n2912) );
  AND2_X4 U4804 ( .A1(n127), .A2(n2113), .ZN(n3286) );
  AND2_X4 U4805 ( .A1(n171), .A2(n2115), .ZN(n3171) );
  AND2_X4 U4813 ( .A1(n140), .A2(n2114), .ZN(n3144) );
  NOR4_X4 U4821 ( .A1(n2309), .A2(n2055), .A3(n2310), .A4(n3098), .ZN(n3097)
         );
  AND3_X4 U4822 ( .A1(n136), .A2(n3031), .A3(n3032), .ZN(n3030) );
  AND4_X4 U4830 ( .A1(n2124), .A2(n2306), .A3(n2974), .A4(n2975), .ZN(n2973)
         );
  AND4_X4 U4831 ( .A1(n2124), .A2(n2305), .A3(n2285), .A4(n2867), .ZN(n2866)
         );
  AND4_X4 U4835 ( .A1(n2696), .A2(n2844), .A3(n2845), .A4(n2846), .ZN(n2843)
         );
  AND3_X4 U4836 ( .A1(n2821), .A2(n2696), .A3(n2822), .ZN(n2820) );
  AND4_X4 U4839 ( .A1(n2696), .A2(n2798), .A3(n64), .A4(n2799), .ZN(n2797) );
  AND3_X4 U4840 ( .A1(n2776), .A2(n2696), .A3(n2777), .ZN(n2775) );
  AND4_X4 U4843 ( .A1(n2696), .A2(n2751), .A3(n2752), .A4(n2753), .ZN(n2750)
         );
  AND3_X4 U4844 ( .A1(n58), .A2(n2696), .A3(n2726), .ZN(n2725) );
  AND4_X4 U4847 ( .A1(n61), .A2(n2695), .A3(n2696), .A4(n2697), .ZN(n2694) );
  AND3_X4 U4848 ( .A1(n166), .A2(n2111), .A3(n2598), .ZN(n2597) );
  AND4_X4 U4851 ( .A1(n160), .A2(n2112), .A3(n2262), .A4(n2283), .ZN(n2573) );
  AND4_X4 U4852 ( .A1(n152), .A2(n2107), .A3(n2263), .A4(n2281), .ZN(n2549) );
  AND2_X4 U4853 ( .A1(n109), .A2(n2109), .ZN(n2494) );
  AND4_X4 U4855 ( .A1(n2124), .A2(n2291), .A3(n2234), .A4(n2471), .ZN(n2470)
         );
  AND3_X4 U4856 ( .A1(n100), .A2(n2443), .A3(n2444), .ZN(n2442) );
  NOR3_X4 U4858 ( .A1(n2110), .A2(n2055), .A3(n99), .ZN(n2416) );
  NOR3_X4 U4859 ( .A1(n117), .A2(n2080), .A3(n2081), .ZN(n2079) );
  AND4_X4 U4860 ( .A1(n76), .A2(n2063), .A3(n2064), .A4(n2065), .ZN(n1807) );
  NOR3_X4 U4865 ( .A1(n2054), .A2(n2055), .A3(n2056), .ZN(n1809) );
  AND3_X4 U4866 ( .A1(n192), .A2(n2013), .A3(n2014), .ZN(n1810) );
  INV_X4 U4869 ( .A(n1108), .ZN(n1109) );
  INV_X4 U4870 ( .A(n376), .ZN(n336) );
  INV_X4 U4871 ( .A(n378), .ZN(n338) );
  AND4_X4 U4878 ( .A1(n373), .A2(n336), .A3(n374), .A4(n375), .ZN(n341) );
  OR2_X4 U4882 ( .A1(n213), .A2(n251), .ZN(n211) );
  NOR2_X2 U4883 ( .A1(n42), .A2(n188), .ZN(n54) );
  INV_X4 U7 ( .A(1'b1), .ZN(htrans_o[0]) );
  INV_X4 U23 ( .A(1'b1), .ZN(hsize_o[2]) );
  INV_X4 U30 ( .A(1'b0), .ZN(hprot_o[1]) );
  INV_X4 U68 ( .A(1'b1), .ZN(hmastlock_o) );
  INV_X4 U77 ( .A(1'b1), .ZN(hburst_o[0]) );
  INV_X4 U90 ( .A(1'b1), .ZN(hburst_o[1]) );
  INV_X4 U99 ( .A(1'b1), .ZN(hburst_o[2]) );
  AOI211_X2 U198 ( .C1(n4964), .C2(n1426), .A(n1427), .B(n1428), .ZN(n13870)
         );
  AOI211_X2 U211 ( .C1(n5126), .C2(n1442), .A(n1443), .B(n1444), .ZN(n13795)
         );
  AOI211_X2 U222 ( .C1(n5582), .C2(n1438), .A(n1439), .B(n1440), .ZN(n13813)
         );
  AOI211_X2 U225 ( .C1(n5118), .C2(n1381), .A(n1382), .B(n1383), .ZN(n13989)
         );
  AOI211_X2 U234 ( .C1(n5061), .C2(n1433), .A(n1434), .B(n1435), .ZN(n13835)
         );
  AOI211_X2 U237 ( .C1(n5531), .C2(n1405), .A(n1406), .B(n1407), .ZN(n13919)
         );
  AOI211_X2 U240 ( .C1(n5529), .C2(n1399), .A(n1400), .B(n1401), .ZN(n13932)
         );
  AOI211_X2 U572 ( .C1(n5524), .C2(n1420), .A(n1421), .B(n1422), .ZN(n13894)
         );
  AOI211_X2 U578 ( .C1(n5525), .C2(n1387), .A(n1388), .B(n1389), .ZN(n13963)
         );
  AOI211_X2 U814 ( .C1(n5527), .C2(n1393), .A(n1394), .B(n1395), .ZN(n13951)
         );
  OAI222_X2 U815 ( .A1(n1148), .A2(n17103), .B1(n4821), .B2(n16792), .C1(n4761), .C2(n17101), .ZN(n4924) );
  OAI222_X2 U817 ( .A1(n1150), .A2(n17103), .B1(n4819), .B2(n16792), .C1(n4763), .C2(n17101), .ZN(n4926) );
  OAI222_X2 U829 ( .A1(n973), .A2(n17103), .B1(n4824), .B2(n16793), .C1(n4772), 
        .C2(n17100), .ZN(n4942) );
  OAI222_X2 U830 ( .A1(n956), .A2(n318), .B1(n4813), .B2(n16793), .C1(n4850), 
        .C2(n17100), .ZN(n4935) );
  OAI222_X2 U832 ( .A1(n957), .A2(n318), .B1(n4816), .B2(n16793), .C1(n4832), 
        .C2(n17100), .ZN(n4936) );
  OAI222_X2 U842 ( .A1(n963), .A2(n17103), .B1(n4815), .B2(n16793), .C1(n4831), 
        .C2(n17100), .ZN(n4938) );
  CLKBUF_X2 U843 ( .A(n4939), .Z(n17212) );
  OAI222_X2 U846 ( .A1(n1147), .A2(n17103), .B1(n4825), .B2(n16792), .C1(n4828), .C2(n17100), .ZN(n4923) );
  OAI221_X2 U987 ( .B1(n968), .B2(n17103), .C1(n4852), .C2(n17102), .A(n1164), 
        .ZN(n4943) );
  OAI221_X2 U1058 ( .B1(n967), .B2(n17103), .C1(n4853), .C2(n17102), .A(n1165), 
        .ZN(n4944) );
  OAI221_X2 U1062 ( .B1(n871), .B2(n17103), .C1(n5501), .C2(n17101), .A(n872), 
        .ZN(n5784) );
  OAI221_X2 U1066 ( .B1(n876), .B2(n17103), .C1(n5500), .C2(n17101), .A(n877), 
        .ZN(n5786) );
  AOI211_X2 U1070 ( .C1(n1310), .C2(n1311), .A(n1312), .B(n1313), .ZN(n14956)
         );
  AOI211_X2 U1074 ( .C1(n1447), .C2(n1448), .A(n1449), .B(n1450), .ZN(n13758)
         );
  AOI211_X2 U1078 ( .C1(n1411), .C2(n1412), .A(n1413), .B(n1414), .ZN(n13907)
         );
  OAI221_X2 U1082 ( .B1(n5515), .B2(n17109), .C1(n268), .C2(n265), .A(n269), 
        .ZN(n5714) );
  OAI221_X2 U1086 ( .B1(n5074), .B2(n17109), .C1(n280), .C2(n265), .A(n281), 
        .ZN(n5720) );
  OAI221_X2 U1091 ( .B1(n5571), .B2(n17110), .C1(n290), .C2(n17107), .A(n291), 
        .ZN(n5725) );
  OAI221_X2 U1095 ( .B1(n5508), .B2(n17110), .C1(n292), .C2(n17107), .A(n293), 
        .ZN(n5726) );
  OAI221_X2 U1100 ( .B1(n5509), .B2(n17110), .C1(n304), .C2(n17107), .A(n305), 
        .ZN(n5732) );
  OAI221_X2 U1103 ( .B1(n5514), .B2(n17110), .C1(n302), .C2(n17107), .A(n303), 
        .ZN(n5731) );
  OAI221_X2 U4884 ( .B1(n5517), .B2(n17110), .C1(n300), .C2(n17107), .A(n301), 
        .ZN(n5730) );
endmodule


module CORTEXM0DS ( HCLK, HRESETn, HADDR, HBURST, HMASTLOCK, HPROT, HSIZE, 
        HTRANS, HWDATA, HWRITE, HRDATA, HREADY, HRESP, NMI, IRQ, TXEV, RXEV, 
        LOCKUP, SYSRESETREQ, SLEEPING );
  output [31:0] HADDR;
  output [2:0] HBURST;
  output [3:0] HPROT;
  output [2:0] HSIZE;
  output [1:0] HTRANS;
  output [31:0] HWDATA;
  input [31:0] HRDATA;
  input [15:0] IRQ;
  input HCLK, HRESETn, HREADY, HRESP, NMI, RXEV;
  output HMASTLOCK, HWRITE, TXEV, LOCKUP, SYSRESETREQ, SLEEPING;
  wire   SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414,
         SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416,
         SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418,
         SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420,
         SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422,
         SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424,
         SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426,
         SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428,
         SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430,
         SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432,
         SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434,
         SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436,
         SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438,
         SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440,
         SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442,
         SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444,
         SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446,
         SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448,
         SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450,
         SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452,
         SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454,
         SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456,
         SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458,
         SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460,
         SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462,
         SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464,
         SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466,
         SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468,
         SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470,
         SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472,
         SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474,
         SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476,
         SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478,
         SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480,
         SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482,
         SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484,
         SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486,
         SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488,
         SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490,
         SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492,
         SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494,
         SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496,
         SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498,
         SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500,
         SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502,
         SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504,
         SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506,
         SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508,
         SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510,
         SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512,
         SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514,
         SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516,
         SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518,
         SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520,
         SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522,
         SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524,
         SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526,
         SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528,
         SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530,
         SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532,
         SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534,
         SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536,
         SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538,
         SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540,
         SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542,
         SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544,
         SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546,
         SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548,
         SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550,
         SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552,
         SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554,
         SYNOPSYS_UNCONNECTED_555;

  cortexm0ds_logic u_logic ( .hclk(HCLK), .hreset_n(HRESETn), .haddr_o(HADDR), 
        .hburst_o({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3}), .hprot_o({HPROT[3:2], SYNOPSYS_UNCONNECTED_4, 
        HPROT[0]}), .hsize_o({SYNOPSYS_UNCONNECTED_5, HSIZE[1:0]}), .htrans_o(
        {HTRANS[1], SYNOPSYS_UNCONNECTED_6}), .hwdata_o(HWDATA), .hwrite_o(
        HWRITE), .hrdata_i(HRDATA), .hready_i(HREADY), .hresp_i(HRESP), 
        .nmi_i(NMI), .irq_i(IRQ), .txev_o(TXEV), .rxev_i(RXEV), .lockup_o(
        LOCKUP), .sys_reset_req_o(SYSRESETREQ), .sleeping_o(SLEEPING), 
        .vis_r0_o({SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38}), .vis_r1_o({
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70}), .vis_r2_o({
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102}), .vis_r3_o({
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, 
        SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, 
        SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112, 
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114, 
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, 
        SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, 
        SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120, 
        SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130, 
        SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, 
        SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134}), .vis_r4_o({
        SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136, 
        SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, 
        SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166}), .vis_r5_o({
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184, 
        SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186, 
        SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188, 
        SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190, 
        SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192, 
        SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194, 
        SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196, 
        SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198}), .vis_r6_o({
        SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200, 
        SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202, 
        SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204, 
        SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206, 
        SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208, 
        SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210, 
        SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212, 
        SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214, 
        SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216, 
        SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218, 
        SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220, 
        SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222, 
        SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224, 
        SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226, 
        SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228, 
        SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230}), .vis_r7_o({
        SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232, 
        SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234, 
        SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236, 
        SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238, 
        SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240, 
        SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242, 
        SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244, 
        SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246, 
        SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248, 
        SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250, 
        SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252, 
        SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254, 
        SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256, 
        SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258, 
        SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260, 
        SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262}), .vis_r8_o({
        SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264, 
        SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266, 
        SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268, 
        SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270, 
        SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272, 
        SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274, 
        SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276, 
        SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278, 
        SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280, 
        SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282, 
        SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284, 
        SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286, 
        SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294}), .vis_r9_o({
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, 
        SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314, 
        SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316, 
        SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318, 
        SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320, 
        SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322, 
        SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324, 
        SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326}), .vis_r10_o({
        SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328, 
        SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330, 
        SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332, 
        SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334, 
        SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336, 
        SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, 
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358}), .vis_r11_o({
        SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, 
        SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380, 
        SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382, 
        SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384, 
        SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386, 
        SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388, 
        SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390}), .vis_r12_o({
        SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392, 
        SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394, 
        SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396, 
        SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398, 
        SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400, 
        SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402, 
        SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404, 
        SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406, 
        SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408, 
        SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410, 
        SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412, 
        SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414, 
        SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416, 
        SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418, 
        SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420, 
        SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422}), .vis_r14_o({
        SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424, 
        SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426, 
        SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428, 
        SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430, 
        SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432, 
        SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434, 
        SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436, 
        SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438, 
        SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440, 
        SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442, 
        SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444, 
        SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446, 
        SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448, 
        SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450, 
        SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452, 
        SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454}), .vis_msp_o({
        SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456, 
        SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458, 
        SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460, 
        SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462, 
        SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464, 
        SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466, 
        SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468, 
        SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470, 
        SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472, 
        SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474, 
        SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476, 
        SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478, 
        SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480, 
        SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482, 
        SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484}), .vis_psp_o({
        SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486, 
        SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488, 
        SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490, 
        SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492, 
        SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494, 
        SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496, 
        SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498, 
        SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500, 
        SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502, 
        SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504, 
        SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506, 
        SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508, 
        SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510, 
        SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512, 
        SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514}), .vis_pc_o({
        SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516, 
        SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518, 
        SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520, 
        SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522, 
        SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524, 
        SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526, 
        SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528, 
        SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530, 
        SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532, 
        SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534, 
        SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536, 
        SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538, 
        SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540, 
        SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542, 
        SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544, 
        SYNOPSYS_UNCONNECTED_545}), .vis_apsr_o({SYNOPSYS_UNCONNECTED_546, 
        SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548, 
        SYNOPSYS_UNCONNECTED_549}), .vis_ipsr_o({SYNOPSYS_UNCONNECTED_550, 
        SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552, 
        SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554, 
        SYNOPSYS_UNCONNECTED_555}) );
  INV_X4 U1 ( .A(1'b1), .ZN(HTRANS[0]) );
  INV_X4 U3 ( .A(1'b1), .ZN(HSIZE[2]) );
  INV_X4 U5 ( .A(1'b0), .ZN(HPROT[1]) );
  INV_X4 U7 ( .A(1'b1), .ZN(HMASTLOCK) );
  INV_X4 U9 ( .A(1'b1), .ZN(HBURST[0]) );
  INV_X4 U11 ( .A(1'b1), .ZN(HBURST[1]) );
  INV_X4 U13 ( .A(1'b1), .ZN(HBURST[2]) );
endmodule

